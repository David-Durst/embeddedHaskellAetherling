module FIFO(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7,
  output [31:0] O_8,
  output [31:0] O_9,
  output [31:0] O_10,
  output [31:0] O_11,
  output [31:0] O_12,
  output [31:0] O_13,
  output [31:0] O_14,
  output [31:0] O_15
);
  reg [31:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [31:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [31:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [31:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [31:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [31:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [31:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [31:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [31:0] _T__8; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [31:0] _T__9; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [31:0] _T__10; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [31:0] _T__11; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [31:0] _T__12; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [31:0] _T__13; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [31:0] _T__14; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [31:0] _T__15; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_16;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
  assign O_8 = _T__8; // @[FIFO.scala 14:7]
  assign O_9 = _T__9; // @[FIFO.scala 14:7]
  assign O_10 = _T__10; // @[FIFO.scala 14:7]
  assign O_11 = _T__11; // @[FIFO.scala 14:7]
  assign O_12 = _T__12; // @[FIFO.scala 14:7]
  assign O_13 = _T__13; // @[FIFO.scala 14:7]
  assign O_14 = _T__14; // @[FIFO.scala 14:7]
  assign O_15 = _T__15; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    _T__8 <= I_8;
    _T__9 <= I_9;
    _T__10 <= I_10;
    _T__11 <= I_11;
    _T__12 <= I_12;
    _T__13 <= I_13;
    _T__14 <= I_14;
    _T__15 <= I_15;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input         clock,
  input         RE,
  input  [6:0]  RADDR,
  output [31:0] RDATA_0,
  output [31:0] RDATA_1,
  output [31:0] RDATA_2,
  output [31:0] RDATA_3,
  output [31:0] RDATA_4,
  output [31:0] RDATA_5,
  output [31:0] RDATA_6,
  output [31:0] RDATA_7,
  output [31:0] RDATA_8,
  output [31:0] RDATA_9,
  output [31:0] RDATA_10,
  output [31:0] RDATA_11,
  output [31:0] RDATA_12,
  output [31:0] RDATA_13,
  output [31:0] RDATA_14,
  output [31:0] RDATA_15,
  input         WE,
  input  [6:0]  WADDR,
  input  [31:0] WDATA_0,
  input  [31:0] WDATA_1,
  input  [31:0] WDATA_2,
  input  [31:0] WDATA_3,
  input  [31:0] WDATA_4,
  input  [31:0] WDATA_5,
  input  [31:0] WDATA_6,
  input  [31:0] WDATA_7,
  input  [31:0] WDATA_8,
  input  [31:0] WDATA_9,
  input  [31:0] WDATA_10,
  input  [31:0] WDATA_11,
  input  [31:0] WDATA_12,
  input  [31:0] WDATA_13,
  input  [31:0] WDATA_14,
  input  [31:0] WDATA_15
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [511:0] ram [0:119]; // @[RAM_ST.scala 29:24]
  reg [511:0] _RAND_0;
  wire [511:0] ram__T_23_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram__T_23_addr; // @[RAM_ST.scala 29:24]
  reg [511:0] _RAND_1;
  wire [511:0] ram__T_17_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram__T_17_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_17_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_17_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_23_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [6:0] ram__T_23_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [6:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _T; // @[RAM_ST.scala 31:71]
  wire [255:0] _T_8; // @[RAM_ST.scala 31:115]
  wire [255:0] _T_15; // @[RAM_ST.scala 31:115]
  wire [6:0] _GEN_126; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_127; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_128; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_129; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_130; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_131; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_132; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_133; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_134; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_135; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_136; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_137; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_138; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_139; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_140; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_141; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_142; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_143; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_144; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_145; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_146; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_147; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_148; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_149; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_150; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_151; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_152; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_153; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_154; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_155; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_156; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_157; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_158; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_159; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_160; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_161; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_162; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_163; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_164; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_165; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_166; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_167; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_168; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_169; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_170; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_171; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_172; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_173; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_174; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_175; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_176; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_177; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_178; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_179; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_180; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_181; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_182; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_183; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_184; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_185; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_186; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_187; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_188; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_189; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_190; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_191; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_192; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_193; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_194; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_195; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_196; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_197; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_198; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_199; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_200; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_201; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_202; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_203; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_204; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_205; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_206; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_207; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_208; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_209; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_210; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_211; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_212; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_213; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_214; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_215; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_216; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_217; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_218; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_219; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_220; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_221; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_222; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_223; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_224; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_225; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_226; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_227; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_228; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_229; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_230; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_231; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_232; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_233; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_234; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_235; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_236; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_237; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_238; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_239; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_240; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_241; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_242; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_243; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_244; // @[RAM_ST.scala 32:46]
  wire [7:0] _T_18; // @[RAM_ST.scala 32:46]
  wire [511:0] _T_25;
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_23_addr = ram__T_23_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_23_data = ram[ram__T_23_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_23_data = ram__T_23_addr >= 7'h78 ? _RAND_1[511:0] : ram[ram__T_23_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_17_data = {_T_15,_T_8};
  assign ram__T_17_addr = _T[6:0];
  assign ram__T_17_mask = 1'h1;
  assign ram__T_17_en = write_elem_counter_valid;
  assign _GEN_1 = 7'h1 == WADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 7'h2 == WADDR ? 7'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 7'h3 == WADDR ? 7'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 7'h4 == WADDR ? 7'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 7'h5 == WADDR ? 7'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 7'h6 == WADDR ? 7'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 7'h7 == WADDR ? 7'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 7'h8 == WADDR ? 7'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 7'h9 == WADDR ? 7'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 7'ha == WADDR ? 7'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 7'hb == WADDR ? 7'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 7'hc == WADDR ? 7'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 7'hd == WADDR ? 7'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 7'he == WADDR ? 7'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 7'hf == WADDR ? 7'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 7'h10 == WADDR ? 7'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 7'h11 == WADDR ? 7'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 7'h12 == WADDR ? 7'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 7'h13 == WADDR ? 7'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 7'h14 == WADDR ? 7'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 7'h15 == WADDR ? 7'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 7'h16 == WADDR ? 7'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 7'h17 == WADDR ? 7'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 7'h18 == WADDR ? 7'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 7'h19 == WADDR ? 7'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 7'h1a == WADDR ? 7'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 7'h1b == WADDR ? 7'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 7'h1c == WADDR ? 7'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 7'h1d == WADDR ? 7'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 7'h1e == WADDR ? 7'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 7'h1f == WADDR ? 7'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 7'h20 == WADDR ? 7'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 7'h21 == WADDR ? 7'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 7'h22 == WADDR ? 7'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 7'h23 == WADDR ? 7'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 7'h24 == WADDR ? 7'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 7'h25 == WADDR ? 7'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 7'h26 == WADDR ? 7'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 7'h27 == WADDR ? 7'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 7'h28 == WADDR ? 7'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 7'h29 == WADDR ? 7'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 7'h2a == WADDR ? 7'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 7'h2b == WADDR ? 7'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 7'h2c == WADDR ? 7'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 7'h2d == WADDR ? 7'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 7'h2e == WADDR ? 7'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 7'h2f == WADDR ? 7'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 7'h30 == WADDR ? 7'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 7'h31 == WADDR ? 7'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 7'h32 == WADDR ? 7'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 7'h33 == WADDR ? 7'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 7'h34 == WADDR ? 7'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 7'h35 == WADDR ? 7'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 7'h36 == WADDR ? 7'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 7'h37 == WADDR ? 7'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 7'h38 == WADDR ? 7'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 7'h39 == WADDR ? 7'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 7'h3a == WADDR ? 7'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 7'h3b == WADDR ? 7'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 7'h3c == WADDR ? 7'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 7'h3d == WADDR ? 7'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 7'h3e == WADDR ? 7'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 7'h3f == WADDR ? 7'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 7'h40 == WADDR ? 7'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 7'h41 == WADDR ? 7'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 7'h42 == WADDR ? 7'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 7'h43 == WADDR ? 7'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 7'h44 == WADDR ? 7'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 7'h45 == WADDR ? 7'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 7'h46 == WADDR ? 7'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 7'h47 == WADDR ? 7'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 7'h48 == WADDR ? 7'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 7'h49 == WADDR ? 7'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 7'h4a == WADDR ? 7'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 7'h4b == WADDR ? 7'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 7'h4c == WADDR ? 7'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 7'h4d == WADDR ? 7'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 7'h4e == WADDR ? 7'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 7'h4f == WADDR ? 7'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 7'h50 == WADDR ? 7'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 7'h51 == WADDR ? 7'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 7'h52 == WADDR ? 7'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 7'h53 == WADDR ? 7'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 7'h54 == WADDR ? 7'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 7'h55 == WADDR ? 7'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 7'h56 == WADDR ? 7'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 7'h57 == WADDR ? 7'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 7'h58 == WADDR ? 7'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 7'h59 == WADDR ? 7'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 7'h5a == WADDR ? 7'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 7'h5b == WADDR ? 7'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 7'h5c == WADDR ? 7'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 7'h5d == WADDR ? 7'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 7'h5e == WADDR ? 7'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 7'h5f == WADDR ? 7'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 7'h60 == WADDR ? 7'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 7'h61 == WADDR ? 7'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 7'h62 == WADDR ? 7'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 7'h63 == WADDR ? 7'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 7'h64 == WADDR ? 7'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 7'h65 == WADDR ? 7'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 7'h66 == WADDR ? 7'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 7'h67 == WADDR ? 7'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 7'h68 == WADDR ? 7'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 7'h69 == WADDR ? 7'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 7'h6a == WADDR ? 7'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 7'h6b == WADDR ? 7'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 7'h6c == WADDR ? 7'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 7'h6d == WADDR ? 7'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 7'h6e == WADDR ? 7'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 7'h6f == WADDR ? 7'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 7'h70 == WADDR ? 7'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 7'h71 == WADDR ? 7'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 7'h72 == WADDR ? 7'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 7'h73 == WADDR ? 7'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 7'h74 == WADDR ? 7'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 7'h75 == WADDR ? 7'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 7'h76 == WADDR ? 7'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 7'h77 == WADDR ? 7'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_119}; // @[RAM_ST.scala 31:71]
  assign _T_8 = {WDATA_7,WDATA_6,WDATA_5,WDATA_4,WDATA_3,WDATA_2,WDATA_1,WDATA_0}; // @[RAM_ST.scala 31:115]
  assign _T_15 = {WDATA_15,WDATA_14,WDATA_13,WDATA_12,WDATA_11,WDATA_10,WDATA_9,WDATA_8}; // @[RAM_ST.scala 31:115]
  assign _GEN_126 = 7'h1 == RADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_127 = 7'h2 == RADDR ? 7'h2 : _GEN_126; // @[RAM_ST.scala 32:46]
  assign _GEN_128 = 7'h3 == RADDR ? 7'h3 : _GEN_127; // @[RAM_ST.scala 32:46]
  assign _GEN_129 = 7'h4 == RADDR ? 7'h4 : _GEN_128; // @[RAM_ST.scala 32:46]
  assign _GEN_130 = 7'h5 == RADDR ? 7'h5 : _GEN_129; // @[RAM_ST.scala 32:46]
  assign _GEN_131 = 7'h6 == RADDR ? 7'h6 : _GEN_130; // @[RAM_ST.scala 32:46]
  assign _GEN_132 = 7'h7 == RADDR ? 7'h7 : _GEN_131; // @[RAM_ST.scala 32:46]
  assign _GEN_133 = 7'h8 == RADDR ? 7'h8 : _GEN_132; // @[RAM_ST.scala 32:46]
  assign _GEN_134 = 7'h9 == RADDR ? 7'h9 : _GEN_133; // @[RAM_ST.scala 32:46]
  assign _GEN_135 = 7'ha == RADDR ? 7'ha : _GEN_134; // @[RAM_ST.scala 32:46]
  assign _GEN_136 = 7'hb == RADDR ? 7'hb : _GEN_135; // @[RAM_ST.scala 32:46]
  assign _GEN_137 = 7'hc == RADDR ? 7'hc : _GEN_136; // @[RAM_ST.scala 32:46]
  assign _GEN_138 = 7'hd == RADDR ? 7'hd : _GEN_137; // @[RAM_ST.scala 32:46]
  assign _GEN_139 = 7'he == RADDR ? 7'he : _GEN_138; // @[RAM_ST.scala 32:46]
  assign _GEN_140 = 7'hf == RADDR ? 7'hf : _GEN_139; // @[RAM_ST.scala 32:46]
  assign _GEN_141 = 7'h10 == RADDR ? 7'h10 : _GEN_140; // @[RAM_ST.scala 32:46]
  assign _GEN_142 = 7'h11 == RADDR ? 7'h11 : _GEN_141; // @[RAM_ST.scala 32:46]
  assign _GEN_143 = 7'h12 == RADDR ? 7'h12 : _GEN_142; // @[RAM_ST.scala 32:46]
  assign _GEN_144 = 7'h13 == RADDR ? 7'h13 : _GEN_143; // @[RAM_ST.scala 32:46]
  assign _GEN_145 = 7'h14 == RADDR ? 7'h14 : _GEN_144; // @[RAM_ST.scala 32:46]
  assign _GEN_146 = 7'h15 == RADDR ? 7'h15 : _GEN_145; // @[RAM_ST.scala 32:46]
  assign _GEN_147 = 7'h16 == RADDR ? 7'h16 : _GEN_146; // @[RAM_ST.scala 32:46]
  assign _GEN_148 = 7'h17 == RADDR ? 7'h17 : _GEN_147; // @[RAM_ST.scala 32:46]
  assign _GEN_149 = 7'h18 == RADDR ? 7'h18 : _GEN_148; // @[RAM_ST.scala 32:46]
  assign _GEN_150 = 7'h19 == RADDR ? 7'h19 : _GEN_149; // @[RAM_ST.scala 32:46]
  assign _GEN_151 = 7'h1a == RADDR ? 7'h1a : _GEN_150; // @[RAM_ST.scala 32:46]
  assign _GEN_152 = 7'h1b == RADDR ? 7'h1b : _GEN_151; // @[RAM_ST.scala 32:46]
  assign _GEN_153 = 7'h1c == RADDR ? 7'h1c : _GEN_152; // @[RAM_ST.scala 32:46]
  assign _GEN_154 = 7'h1d == RADDR ? 7'h1d : _GEN_153; // @[RAM_ST.scala 32:46]
  assign _GEN_155 = 7'h1e == RADDR ? 7'h1e : _GEN_154; // @[RAM_ST.scala 32:46]
  assign _GEN_156 = 7'h1f == RADDR ? 7'h1f : _GEN_155; // @[RAM_ST.scala 32:46]
  assign _GEN_157 = 7'h20 == RADDR ? 7'h20 : _GEN_156; // @[RAM_ST.scala 32:46]
  assign _GEN_158 = 7'h21 == RADDR ? 7'h21 : _GEN_157; // @[RAM_ST.scala 32:46]
  assign _GEN_159 = 7'h22 == RADDR ? 7'h22 : _GEN_158; // @[RAM_ST.scala 32:46]
  assign _GEN_160 = 7'h23 == RADDR ? 7'h23 : _GEN_159; // @[RAM_ST.scala 32:46]
  assign _GEN_161 = 7'h24 == RADDR ? 7'h24 : _GEN_160; // @[RAM_ST.scala 32:46]
  assign _GEN_162 = 7'h25 == RADDR ? 7'h25 : _GEN_161; // @[RAM_ST.scala 32:46]
  assign _GEN_163 = 7'h26 == RADDR ? 7'h26 : _GEN_162; // @[RAM_ST.scala 32:46]
  assign _GEN_164 = 7'h27 == RADDR ? 7'h27 : _GEN_163; // @[RAM_ST.scala 32:46]
  assign _GEN_165 = 7'h28 == RADDR ? 7'h28 : _GEN_164; // @[RAM_ST.scala 32:46]
  assign _GEN_166 = 7'h29 == RADDR ? 7'h29 : _GEN_165; // @[RAM_ST.scala 32:46]
  assign _GEN_167 = 7'h2a == RADDR ? 7'h2a : _GEN_166; // @[RAM_ST.scala 32:46]
  assign _GEN_168 = 7'h2b == RADDR ? 7'h2b : _GEN_167; // @[RAM_ST.scala 32:46]
  assign _GEN_169 = 7'h2c == RADDR ? 7'h2c : _GEN_168; // @[RAM_ST.scala 32:46]
  assign _GEN_170 = 7'h2d == RADDR ? 7'h2d : _GEN_169; // @[RAM_ST.scala 32:46]
  assign _GEN_171 = 7'h2e == RADDR ? 7'h2e : _GEN_170; // @[RAM_ST.scala 32:46]
  assign _GEN_172 = 7'h2f == RADDR ? 7'h2f : _GEN_171; // @[RAM_ST.scala 32:46]
  assign _GEN_173 = 7'h30 == RADDR ? 7'h30 : _GEN_172; // @[RAM_ST.scala 32:46]
  assign _GEN_174 = 7'h31 == RADDR ? 7'h31 : _GEN_173; // @[RAM_ST.scala 32:46]
  assign _GEN_175 = 7'h32 == RADDR ? 7'h32 : _GEN_174; // @[RAM_ST.scala 32:46]
  assign _GEN_176 = 7'h33 == RADDR ? 7'h33 : _GEN_175; // @[RAM_ST.scala 32:46]
  assign _GEN_177 = 7'h34 == RADDR ? 7'h34 : _GEN_176; // @[RAM_ST.scala 32:46]
  assign _GEN_178 = 7'h35 == RADDR ? 7'h35 : _GEN_177; // @[RAM_ST.scala 32:46]
  assign _GEN_179 = 7'h36 == RADDR ? 7'h36 : _GEN_178; // @[RAM_ST.scala 32:46]
  assign _GEN_180 = 7'h37 == RADDR ? 7'h37 : _GEN_179; // @[RAM_ST.scala 32:46]
  assign _GEN_181 = 7'h38 == RADDR ? 7'h38 : _GEN_180; // @[RAM_ST.scala 32:46]
  assign _GEN_182 = 7'h39 == RADDR ? 7'h39 : _GEN_181; // @[RAM_ST.scala 32:46]
  assign _GEN_183 = 7'h3a == RADDR ? 7'h3a : _GEN_182; // @[RAM_ST.scala 32:46]
  assign _GEN_184 = 7'h3b == RADDR ? 7'h3b : _GEN_183; // @[RAM_ST.scala 32:46]
  assign _GEN_185 = 7'h3c == RADDR ? 7'h3c : _GEN_184; // @[RAM_ST.scala 32:46]
  assign _GEN_186 = 7'h3d == RADDR ? 7'h3d : _GEN_185; // @[RAM_ST.scala 32:46]
  assign _GEN_187 = 7'h3e == RADDR ? 7'h3e : _GEN_186; // @[RAM_ST.scala 32:46]
  assign _GEN_188 = 7'h3f == RADDR ? 7'h3f : _GEN_187; // @[RAM_ST.scala 32:46]
  assign _GEN_189 = 7'h40 == RADDR ? 7'h40 : _GEN_188; // @[RAM_ST.scala 32:46]
  assign _GEN_190 = 7'h41 == RADDR ? 7'h41 : _GEN_189; // @[RAM_ST.scala 32:46]
  assign _GEN_191 = 7'h42 == RADDR ? 7'h42 : _GEN_190; // @[RAM_ST.scala 32:46]
  assign _GEN_192 = 7'h43 == RADDR ? 7'h43 : _GEN_191; // @[RAM_ST.scala 32:46]
  assign _GEN_193 = 7'h44 == RADDR ? 7'h44 : _GEN_192; // @[RAM_ST.scala 32:46]
  assign _GEN_194 = 7'h45 == RADDR ? 7'h45 : _GEN_193; // @[RAM_ST.scala 32:46]
  assign _GEN_195 = 7'h46 == RADDR ? 7'h46 : _GEN_194; // @[RAM_ST.scala 32:46]
  assign _GEN_196 = 7'h47 == RADDR ? 7'h47 : _GEN_195; // @[RAM_ST.scala 32:46]
  assign _GEN_197 = 7'h48 == RADDR ? 7'h48 : _GEN_196; // @[RAM_ST.scala 32:46]
  assign _GEN_198 = 7'h49 == RADDR ? 7'h49 : _GEN_197; // @[RAM_ST.scala 32:46]
  assign _GEN_199 = 7'h4a == RADDR ? 7'h4a : _GEN_198; // @[RAM_ST.scala 32:46]
  assign _GEN_200 = 7'h4b == RADDR ? 7'h4b : _GEN_199; // @[RAM_ST.scala 32:46]
  assign _GEN_201 = 7'h4c == RADDR ? 7'h4c : _GEN_200; // @[RAM_ST.scala 32:46]
  assign _GEN_202 = 7'h4d == RADDR ? 7'h4d : _GEN_201; // @[RAM_ST.scala 32:46]
  assign _GEN_203 = 7'h4e == RADDR ? 7'h4e : _GEN_202; // @[RAM_ST.scala 32:46]
  assign _GEN_204 = 7'h4f == RADDR ? 7'h4f : _GEN_203; // @[RAM_ST.scala 32:46]
  assign _GEN_205 = 7'h50 == RADDR ? 7'h50 : _GEN_204; // @[RAM_ST.scala 32:46]
  assign _GEN_206 = 7'h51 == RADDR ? 7'h51 : _GEN_205; // @[RAM_ST.scala 32:46]
  assign _GEN_207 = 7'h52 == RADDR ? 7'h52 : _GEN_206; // @[RAM_ST.scala 32:46]
  assign _GEN_208 = 7'h53 == RADDR ? 7'h53 : _GEN_207; // @[RAM_ST.scala 32:46]
  assign _GEN_209 = 7'h54 == RADDR ? 7'h54 : _GEN_208; // @[RAM_ST.scala 32:46]
  assign _GEN_210 = 7'h55 == RADDR ? 7'h55 : _GEN_209; // @[RAM_ST.scala 32:46]
  assign _GEN_211 = 7'h56 == RADDR ? 7'h56 : _GEN_210; // @[RAM_ST.scala 32:46]
  assign _GEN_212 = 7'h57 == RADDR ? 7'h57 : _GEN_211; // @[RAM_ST.scala 32:46]
  assign _GEN_213 = 7'h58 == RADDR ? 7'h58 : _GEN_212; // @[RAM_ST.scala 32:46]
  assign _GEN_214 = 7'h59 == RADDR ? 7'h59 : _GEN_213; // @[RAM_ST.scala 32:46]
  assign _GEN_215 = 7'h5a == RADDR ? 7'h5a : _GEN_214; // @[RAM_ST.scala 32:46]
  assign _GEN_216 = 7'h5b == RADDR ? 7'h5b : _GEN_215; // @[RAM_ST.scala 32:46]
  assign _GEN_217 = 7'h5c == RADDR ? 7'h5c : _GEN_216; // @[RAM_ST.scala 32:46]
  assign _GEN_218 = 7'h5d == RADDR ? 7'h5d : _GEN_217; // @[RAM_ST.scala 32:46]
  assign _GEN_219 = 7'h5e == RADDR ? 7'h5e : _GEN_218; // @[RAM_ST.scala 32:46]
  assign _GEN_220 = 7'h5f == RADDR ? 7'h5f : _GEN_219; // @[RAM_ST.scala 32:46]
  assign _GEN_221 = 7'h60 == RADDR ? 7'h60 : _GEN_220; // @[RAM_ST.scala 32:46]
  assign _GEN_222 = 7'h61 == RADDR ? 7'h61 : _GEN_221; // @[RAM_ST.scala 32:46]
  assign _GEN_223 = 7'h62 == RADDR ? 7'h62 : _GEN_222; // @[RAM_ST.scala 32:46]
  assign _GEN_224 = 7'h63 == RADDR ? 7'h63 : _GEN_223; // @[RAM_ST.scala 32:46]
  assign _GEN_225 = 7'h64 == RADDR ? 7'h64 : _GEN_224; // @[RAM_ST.scala 32:46]
  assign _GEN_226 = 7'h65 == RADDR ? 7'h65 : _GEN_225; // @[RAM_ST.scala 32:46]
  assign _GEN_227 = 7'h66 == RADDR ? 7'h66 : _GEN_226; // @[RAM_ST.scala 32:46]
  assign _GEN_228 = 7'h67 == RADDR ? 7'h67 : _GEN_227; // @[RAM_ST.scala 32:46]
  assign _GEN_229 = 7'h68 == RADDR ? 7'h68 : _GEN_228; // @[RAM_ST.scala 32:46]
  assign _GEN_230 = 7'h69 == RADDR ? 7'h69 : _GEN_229; // @[RAM_ST.scala 32:46]
  assign _GEN_231 = 7'h6a == RADDR ? 7'h6a : _GEN_230; // @[RAM_ST.scala 32:46]
  assign _GEN_232 = 7'h6b == RADDR ? 7'h6b : _GEN_231; // @[RAM_ST.scala 32:46]
  assign _GEN_233 = 7'h6c == RADDR ? 7'h6c : _GEN_232; // @[RAM_ST.scala 32:46]
  assign _GEN_234 = 7'h6d == RADDR ? 7'h6d : _GEN_233; // @[RAM_ST.scala 32:46]
  assign _GEN_235 = 7'h6e == RADDR ? 7'h6e : _GEN_234; // @[RAM_ST.scala 32:46]
  assign _GEN_236 = 7'h6f == RADDR ? 7'h6f : _GEN_235; // @[RAM_ST.scala 32:46]
  assign _GEN_237 = 7'h70 == RADDR ? 7'h70 : _GEN_236; // @[RAM_ST.scala 32:46]
  assign _GEN_238 = 7'h71 == RADDR ? 7'h71 : _GEN_237; // @[RAM_ST.scala 32:46]
  assign _GEN_239 = 7'h72 == RADDR ? 7'h72 : _GEN_238; // @[RAM_ST.scala 32:46]
  assign _GEN_240 = 7'h73 == RADDR ? 7'h73 : _GEN_239; // @[RAM_ST.scala 32:46]
  assign _GEN_241 = 7'h74 == RADDR ? 7'h74 : _GEN_240; // @[RAM_ST.scala 32:46]
  assign _GEN_242 = 7'h75 == RADDR ? 7'h75 : _GEN_241; // @[RAM_ST.scala 32:46]
  assign _GEN_243 = 7'h76 == RADDR ? 7'h76 : _GEN_242; // @[RAM_ST.scala 32:46]
  assign _GEN_244 = 7'h77 == RADDR ? 7'h77 : _GEN_243; // @[RAM_ST.scala 32:46]
  assign _T_18 = {{1'd0}, _GEN_244}; // @[RAM_ST.scala 32:46]
  assign _T_25 = ram__T_23_data;
  assign RDATA_0 = _T_25[31:0]; // @[RAM_ST.scala 32:9]
  assign RDATA_1 = _T_25[63:32]; // @[RAM_ST.scala 32:9]
  assign RDATA_2 = _T_25[95:64]; // @[RAM_ST.scala 32:9]
  assign RDATA_3 = _T_25[127:96]; // @[RAM_ST.scala 32:9]
  assign RDATA_4 = _T_25[159:128]; // @[RAM_ST.scala 32:9]
  assign RDATA_5 = _T_25[191:160]; // @[RAM_ST.scala 32:9]
  assign RDATA_6 = _T_25[223:192]; // @[RAM_ST.scala 32:9]
  assign RDATA_7 = _T_25[255:224]; // @[RAM_ST.scala 32:9]
  assign RDATA_8 = _T_25[287:256]; // @[RAM_ST.scala 32:9]
  assign RDATA_9 = _T_25[319:288]; // @[RAM_ST.scala 32:9]
  assign RDATA_10 = _T_25[351:320]; // @[RAM_ST.scala 32:9]
  assign RDATA_11 = _T_25[383:352]; // @[RAM_ST.scala 32:9]
  assign RDATA_12 = _T_25[415:384]; // @[RAM_ST.scala 32:9]
  assign RDATA_13 = _T_25[447:416]; // @[RAM_ST.scala 32:9]
  assign RDATA_14 = _T_25[479:448]; // @[RAM_ST.scala 32:9]
  assign RDATA_15 = _T_25[511:480]; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {16{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 120; initvar = initvar+1)
    ram[initvar] = _RAND_0[511:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {16{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_23_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_23_addr_pipe_0 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_17_en & ram__T_17_mask) begin
      ram[ram__T_17_addr] <= ram__T_17_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_23_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_23_addr_pipe_0 <= _T_18[6:0];
    end
  end
endmodule
module ShiftT(
  input         clock,
  input         reset,
  input         valid_up,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7,
  output [31:0] O_8,
  output [31:0] O_9,
  output [31:0] O_10,
  output [31:0] O_11,
  output [31:0] O_12,
  output [31:0] O_13,
  output [31:0] O_14,
  output [31:0] O_15
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_0; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_1; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_2; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_3; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_4; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_5; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_6; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_7; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_8; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_9; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_10; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_11; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_12; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_13; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_14; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_RDATA_15; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_0; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_1; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_2; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_3; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_4; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_5; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_6; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_7; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_8; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_9; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_10; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_11; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_12; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_13; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_14; // @[ShiftT.scala 39:29]
  wire [31:0] RAM_ST_WDATA_15; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [6:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [6:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0(RAM_ST_RDATA_0),
    .RDATA_1(RAM_ST_RDATA_1),
    .RDATA_2(RAM_ST_RDATA_2),
    .RDATA_3(RAM_ST_RDATA_3),
    .RDATA_4(RAM_ST_RDATA_4),
    .RDATA_5(RAM_ST_RDATA_5),
    .RDATA_6(RAM_ST_RDATA_6),
    .RDATA_7(RAM_ST_RDATA_7),
    .RDATA_8(RAM_ST_RDATA_8),
    .RDATA_9(RAM_ST_RDATA_9),
    .RDATA_10(RAM_ST_RDATA_10),
    .RDATA_11(RAM_ST_RDATA_11),
    .RDATA_12(RAM_ST_RDATA_12),
    .RDATA_13(RAM_ST_RDATA_13),
    .RDATA_14(RAM_ST_RDATA_14),
    .RDATA_15(RAM_ST_RDATA_15),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0(RAM_ST_WDATA_0),
    .WDATA_1(RAM_ST_WDATA_1),
    .WDATA_2(RAM_ST_WDATA_2),
    .WDATA_3(RAM_ST_WDATA_3),
    .WDATA_4(RAM_ST_WDATA_4),
    .WDATA_5(RAM_ST_WDATA_5),
    .WDATA_6(RAM_ST_WDATA_6),
    .WDATA_7(RAM_ST_WDATA_7),
    .WDATA_8(RAM_ST_WDATA_8),
    .WDATA_9(RAM_ST_WDATA_9),
    .WDATA_10(RAM_ST_WDATA_10),
    .WDATA_11(RAM_ST_WDATA_11),
    .WDATA_12(RAM_ST_WDATA_12),
    .WDATA_13(RAM_ST_WDATA_13),
    .WDATA_14(RAM_ST_WDATA_14),
    .WDATA_15(RAM_ST_WDATA_15)
  );
  NestedCounters_1 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 7'h77; // @[Counter.scala 37:24]
  assign _T_3 = value + 7'h1; // @[Counter.scala 38:22]
  assign O_0 = RAM_ST_RDATA_0; // @[ShiftT.scala 51:7]
  assign O_1 = RAM_ST_RDATA_1; // @[ShiftT.scala 51:7]
  assign O_2 = RAM_ST_RDATA_2; // @[ShiftT.scala 51:7]
  assign O_3 = RAM_ST_RDATA_3; // @[ShiftT.scala 51:7]
  assign O_4 = RAM_ST_RDATA_4; // @[ShiftT.scala 51:7]
  assign O_5 = RAM_ST_RDATA_5; // @[ShiftT.scala 51:7]
  assign O_6 = RAM_ST_RDATA_6; // @[ShiftT.scala 51:7]
  assign O_7 = RAM_ST_RDATA_7; // @[ShiftT.scala 51:7]
  assign O_8 = RAM_ST_RDATA_8; // @[ShiftT.scala 51:7]
  assign O_9 = RAM_ST_RDATA_9; // @[ShiftT.scala 51:7]
  assign O_10 = RAM_ST_RDATA_10; // @[ShiftT.scala 51:7]
  assign O_11 = RAM_ST_RDATA_11; // @[ShiftT.scala 51:7]
  assign O_12 = RAM_ST_RDATA_12; // @[ShiftT.scala 51:7]
  assign O_13 = RAM_ST_RDATA_13; // @[ShiftT.scala 51:7]
  assign O_14 = RAM_ST_RDATA_14; // @[ShiftT.scala 51:7]
  assign O_15 = RAM_ST_RDATA_15; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 7'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0 = I_0; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_1 = I_1; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_2 = I_2; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_3 = I_3; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_4 = I_4; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_5 = I_5; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_6 = I_6; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_7 = I_7; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_8 = I_8; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_9 = I_9; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_10 = I_10; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_11 = I_11; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_12 = I_12; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_13 = I_13; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_14 = I_14; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_15 = I_15; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 7'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 7'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7,
  output [31:0] O_8,
  output [31:0] O_9,
  output [31:0] O_10,
  output [31:0] O_11,
  output [31:0] O_12,
  output [31:0] O_13,
  output [31:0] O_14,
  output [31:0] O_15
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:26]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_1; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_2; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_3; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_4; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_5; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_6; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_7; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_8; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_9; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_10; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_11; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_12; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_13; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_14; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_15; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_1; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_2; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_3; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_4; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_5; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_6; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_7; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_8; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_9; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_10; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_11; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_12; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_13; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_14; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_15; // @[ShiftTS.scala 32:26]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0(ShiftT_I_0),
    .I_1(ShiftT_I_1),
    .I_2(ShiftT_I_2),
    .I_3(ShiftT_I_3),
    .I_4(ShiftT_I_4),
    .I_5(ShiftT_I_5),
    .I_6(ShiftT_I_6),
    .I_7(ShiftT_I_7),
    .I_8(ShiftT_I_8),
    .I_9(ShiftT_I_9),
    .I_10(ShiftT_I_10),
    .I_11(ShiftT_I_11),
    .I_12(ShiftT_I_12),
    .I_13(ShiftT_I_13),
    .I_14(ShiftT_I_14),
    .I_15(ShiftT_I_15),
    .O_0(ShiftT_O_0),
    .O_1(ShiftT_O_1),
    .O_2(ShiftT_O_2),
    .O_3(ShiftT_O_3),
    .O_4(ShiftT_O_4),
    .O_5(ShiftT_O_5),
    .O_6(ShiftT_O_6),
    .O_7(ShiftT_O_7),
    .O_8(ShiftT_O_8),
    .O_9(ShiftT_O_9),
    .O_10(ShiftT_O_10),
    .O_11(ShiftT_O_11),
    .O_12(ShiftT_O_12),
    .O_13(ShiftT_O_13),
    .O_14(ShiftT_O_14),
    .O_15(ShiftT_O_15)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = ShiftT_O_1; // @[ShiftTS.scala 51:36]
  assign O_2 = ShiftT_O_2; // @[ShiftTS.scala 51:36]
  assign O_3 = ShiftT_O_3; // @[ShiftTS.scala 51:36]
  assign O_4 = ShiftT_O_4; // @[ShiftTS.scala 51:36]
  assign O_5 = ShiftT_O_5; // @[ShiftTS.scala 51:36]
  assign O_6 = ShiftT_O_6; // @[ShiftTS.scala 51:36]
  assign O_7 = ShiftT_O_7; // @[ShiftTS.scala 51:36]
  assign O_8 = ShiftT_O_8; // @[ShiftTS.scala 51:36]
  assign O_9 = ShiftT_O_9; // @[ShiftTS.scala 51:36]
  assign O_10 = ShiftT_O_10; // @[ShiftTS.scala 51:36]
  assign O_11 = ShiftT_O_11; // @[ShiftTS.scala 51:36]
  assign O_12 = ShiftT_O_12; // @[ShiftTS.scala 51:36]
  assign O_13 = ShiftT_O_13; // @[ShiftTS.scala 51:36]
  assign O_14 = ShiftT_O_14; // @[ShiftTS.scala 51:36]
  assign O_15 = ShiftT_O_15; // @[ShiftTS.scala 51:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 53:29]
  assign ShiftT_I_0 = I_0; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_1 = I_1; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_2 = I_2; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_3 = I_3; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_4 = I_4; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_5 = I_5; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_6 = I_6; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_7 = I_7; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_8 = I_8; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_9 = I_9; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_10 = I_10; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_11 = I_11; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_12 = I_12; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_13 = I_13; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_14 = I_14; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_15 = I_15; // @[ShiftTS.scala 50:25]
endmodule
module ShiftT_2(
  input         clock,
  input  [31:0] I_0,
  output [31:0] O_0
);
  reg [31:0] _T_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0 = _T_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= I_0;
  end
endmodule
module ShiftTS_2(
  input         clock,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7,
  output [31:0] O_8,
  output [31:0] O_9,
  output [31:0] O_10,
  output [31:0] O_11,
  output [31:0] O_12,
  output [31:0] O_13,
  output [31:0] O_14,
  output [31:0] O_15
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [31:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  ShiftT_2 ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .I_0(ShiftT_I_0),
    .O_0(ShiftT_O_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = I_0; // @[ShiftTS.scala 40:36]
  assign O_2 = I_1; // @[ShiftTS.scala 40:36]
  assign O_3 = I_2; // @[ShiftTS.scala 40:36]
  assign O_4 = I_3; // @[ShiftTS.scala 40:36]
  assign O_5 = I_4; // @[ShiftTS.scala 40:36]
  assign O_6 = I_5; // @[ShiftTS.scala 40:36]
  assign O_7 = I_6; // @[ShiftTS.scala 40:36]
  assign O_8 = I_7; // @[ShiftTS.scala 40:36]
  assign O_9 = I_8; // @[ShiftTS.scala 40:36]
  assign O_10 = I_9; // @[ShiftTS.scala 40:36]
  assign O_11 = I_10; // @[ShiftTS.scala 40:36]
  assign O_12 = I_11; // @[ShiftTS.scala 40:36]
  assign O_13 = I_12; // @[ShiftTS.scala 40:36]
  assign O_14 = I_13; // @[ShiftTS.scala 40:36]
  assign O_15 = I_14; // @[ShiftTS.scala 40:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0 = I_15; // @[ShiftTS.scala 50:25]
endmodule
module SSeqTupleCreator(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1,
  output [31:0] O_0,
  output [31:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I0_8,
  input  [31:0] I0_9,
  input  [31:0] I0_10,
  input  [31:0] I0_11,
  input  [31:0] I0_12,
  input  [31:0] I0_13,
  input  [31:0] I0_14,
  input  [31:0] I0_15,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  input  [31:0] I1_8,
  input  [31:0] I1_9,
  input  [31:0] I1_10,
  input  [31:0] I1_11,
  input  [31:0] I1_12,
  input  [31:0] I1_13,
  input  [31:0] I1_14,
  input  [31:0] I1_15,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_8_0,
  output [31:0] O_8_1,
  output [31:0] O_9_0,
  output [31:0] O_9_1,
  output [31:0] O_10_0,
  output [31:0] O_10_1,
  output [31:0] O_11_0,
  output [31:0] O_11_1,
  output [31:0] O_12_0,
  output [31:0] O_12_1,
  output [31:0] O_13_0,
  output [31:0] O_13_1,
  output [31:0] O_14_0,
  output [31:0] O_14_1,
  output [31:0] O_15_0,
  output [31:0] O_15_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  SSeqTupleCreator other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  SSeqTupleCreator other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  SSeqTupleCreator other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  SSeqTupleCreator other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  SSeqTupleCreator other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0(other_ops_7_I0),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1)
  );
  SSeqTupleCreator other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0(other_ops_8_I0),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1)
  );
  SSeqTupleCreator other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0(other_ops_9_I0),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1)
  );
  SSeqTupleCreator other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0(other_ops_10_I0),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1)
  );
  SSeqTupleCreator other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0(other_ops_11_I0),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1)
  );
  SSeqTupleCreator other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0(other_ops_12_I0),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1)
  );
  SSeqTupleCreator other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0(other_ops_13_I0),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1)
  );
  SSeqTupleCreator other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0(other_ops_14_I0),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0 = I0_8; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0 = I0_9; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0 = I0_10; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0 = I0_11; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0 = I0_12; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0 = I0_13; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0 = I0_14; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0 = I0_15; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I0_3,
  input  [31:0] I0_4,
  input  [31:0] I0_5,
  input  [31:0] I0_6,
  input  [31:0] I0_7,
  input  [31:0] I0_8,
  input  [31:0] I0_9,
  input  [31:0] I0_10,
  input  [31:0] I0_11,
  input  [31:0] I0_12,
  input  [31:0] I0_13,
  input  [31:0] I0_14,
  input  [31:0] I0_15,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  input  [31:0] I1_8,
  input  [31:0] I1_9,
  input  [31:0] I1_10,
  input  [31:0] I1_11,
  input  [31:0] I1_12,
  input  [31:0] I1_13,
  input  [31:0] I1_14,
  input  [31:0] I1_15,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_8_0,
  output [31:0] O_8_1,
  output [31:0] O_9_0,
  output [31:0] O_9_1,
  output [31:0] O_10_0,
  output [31:0] O_10_1,
  output [31:0] O_11_0,
  output [31:0] O_11_1,
  output [31:0] O_12_0,
  output [31:0] O_12_1,
  output [31:0] O_13_0,
  output [31:0] O_13_1,
  output [31:0] O_14_0,
  output [31:0] O_14_1,
  output [31:0] O_15_0,
  output [31:0] O_15_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I0_8(op_I0_8),
    .I0_9(op_I0_9),
    .I0_10(op_I0_10),
    .I0_11(op_I0_11),
    .I0_12(op_I0_12),
    .I0_13(op_I0_13),
    .I0_14(op_I0_14),
    .I0_15(op_I0_15),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_8_0 = op_O_8_0; // @[Map2T.scala 17:7]
  assign O_8_1 = op_O_8_1; // @[Map2T.scala 17:7]
  assign O_9_0 = op_O_9_0; // @[Map2T.scala 17:7]
  assign O_9_1 = op_O_9_1; // @[Map2T.scala 17:7]
  assign O_10_0 = op_O_10_0; // @[Map2T.scala 17:7]
  assign O_10_1 = op_O_10_1; // @[Map2T.scala 17:7]
  assign O_11_0 = op_O_11_0; // @[Map2T.scala 17:7]
  assign O_11_1 = op_O_11_1; // @[Map2T.scala 17:7]
  assign O_12_0 = op_O_12_0; // @[Map2T.scala 17:7]
  assign O_12_1 = op_O_12_1; // @[Map2T.scala 17:7]
  assign O_13_0 = op_O_13_0; // @[Map2T.scala 17:7]
  assign O_13_1 = op_O_13_1; // @[Map2T.scala 17:7]
  assign O_14_0 = op_O_14_0; // @[Map2T.scala 17:7]
  assign O_14_1 = op_O_14_1; // @[Map2T.scala 17:7]
  assign O_15_0 = op_O_15_0; // @[Map2T.scala 17:7]
  assign O_15_1 = op_O_15_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I0_8 = I0_8; // @[Map2T.scala 15:11]
  assign op_I0_9 = I0_9; // @[Map2T.scala 15:11]
  assign op_I0_10 = I0_10; // @[Map2T.scala 15:11]
  assign op_I0_11 = I0_11; // @[Map2T.scala 15:11]
  assign op_I0_12 = I0_12; // @[Map2T.scala 15:11]
  assign op_I0_13 = I0_13; // @[Map2T.scala 15:11]
  assign op_I0_14 = I0_14; // @[Map2T.scala 15:11]
  assign op_I0_15 = I0_15; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I1,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I0_8_0,
  input  [31:0] I0_8_1,
  input  [31:0] I0_9_0,
  input  [31:0] I0_9_1,
  input  [31:0] I0_10_0,
  input  [31:0] I0_10_1,
  input  [31:0] I0_11_0,
  input  [31:0] I0_11_1,
  input  [31:0] I0_12_0,
  input  [31:0] I0_12_1,
  input  [31:0] I0_13_0,
  input  [31:0] I0_13_1,
  input  [31:0] I0_14_0,
  input  [31:0] I0_14_1,
  input  [31:0] I0_15_0,
  input  [31:0] I0_15_1,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  input  [31:0] I1_8,
  input  [31:0] I1_9,
  input  [31:0] I1_10,
  input  [31:0] I1_11,
  input  [31:0] I1_12,
  input  [31:0] I1_13,
  input  [31:0] I1_14,
  input  [31:0] I1_15,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2,
  output [31:0] O_8_0,
  output [31:0] O_8_1,
  output [31:0] O_8_2,
  output [31:0] O_9_0,
  output [31:0] O_9_1,
  output [31:0] O_9_2,
  output [31:0] O_10_0,
  output [31:0] O_10_1,
  output [31:0] O_10_2,
  output [31:0] O_11_0,
  output [31:0] O_11_1,
  output [31:0] O_11_2,
  output [31:0] O_12_0,
  output [31:0] O_12_1,
  output [31:0] O_12_2,
  output [31:0] O_13_0,
  output [31:0] O_13_1,
  output [31:0] O_13_2,
  output [31:0] O_14_0,
  output [31:0] O_14_1,
  output [31:0] O_14_2,
  output [31:0] O_15_0,
  output [31:0] O_15_1,
  output [31:0] O_15_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  SSeqTupleAppender other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  SSeqTupleAppender other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  SSeqTupleAppender other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  SSeqTupleAppender other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  SSeqTupleAppender other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  SSeqTupleAppender other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  SSeqTupleAppender other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  SSeqTupleAppender other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  SSeqTupleAppender other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  SSeqTupleAppender other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  SSeqTupleAppender other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  SSeqTupleAppender other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_4_2 = other_ops_3_O_2; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_5_2 = other_ops_4_O_2; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_6_2 = other_ops_5_O_2; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_7_2 = other_ops_6_O_2; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_8_2 = other_ops_7_O_2; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_9_2 = other_ops_8_O_2; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_10_2 = other_ops_9_O_2; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_11_2 = other_ops_10_O_2; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_12_2 = other_ops_11_O_2; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_13_2 = other_ops_12_O_2; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_14_2 = other_ops_13_O_2; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign O_15_2 = other_ops_14_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I0_8_0,
  input  [31:0] I0_8_1,
  input  [31:0] I0_9_0,
  input  [31:0] I0_9_1,
  input  [31:0] I0_10_0,
  input  [31:0] I0_10_1,
  input  [31:0] I0_11_0,
  input  [31:0] I0_11_1,
  input  [31:0] I0_12_0,
  input  [31:0] I0_12_1,
  input  [31:0] I0_13_0,
  input  [31:0] I0_13_1,
  input  [31:0] I0_14_0,
  input  [31:0] I0_14_1,
  input  [31:0] I0_15_0,
  input  [31:0] I0_15_1,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  input  [31:0] I1_3,
  input  [31:0] I1_4,
  input  [31:0] I1_5,
  input  [31:0] I1_6,
  input  [31:0] I1_7,
  input  [31:0] I1_8,
  input  [31:0] I1_9,
  input  [31:0] I1_10,
  input  [31:0] I1_11,
  input  [31:0] I1_12,
  input  [31:0] I1_13,
  input  [31:0] I1_14,
  input  [31:0] I1_15,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2,
  output [31:0] O_8_0,
  output [31:0] O_8_1,
  output [31:0] O_8_2,
  output [31:0] O_9_0,
  output [31:0] O_9_1,
  output [31:0] O_9_2,
  output [31:0] O_10_0,
  output [31:0] O_10_1,
  output [31:0] O_10_2,
  output [31:0] O_11_0,
  output [31:0] O_11_1,
  output [31:0] O_11_2,
  output [31:0] O_12_0,
  output [31:0] O_12_1,
  output [31:0] O_12_2,
  output [31:0] O_13_0,
  output [31:0] O_13_1,
  output [31:0] O_13_2,
  output [31:0] O_14_0,
  output [31:0] O_14_1,
  output [31:0] O_14_2,
  output [31:0] O_15_0,
  output [31:0] O_15_1,
  output [31:0] O_15_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_8_2(op_O_8_2),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_9_2(op_O_9_2),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_10_2(op_O_10_2),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_11_2(op_O_11_2),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_12_2(op_O_12_2),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_13_2(op_O_13_2),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_14_2(op_O_14_2),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1),
    .O_15_2(op_O_15_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_2_2 = op_O_2_2; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_3_2 = op_O_3_2; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_4_2 = op_O_4_2; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_5_2 = op_O_5_2; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_6_2 = op_O_6_2; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_7_2 = op_O_7_2; // @[Map2T.scala 17:7]
  assign O_8_0 = op_O_8_0; // @[Map2T.scala 17:7]
  assign O_8_1 = op_O_8_1; // @[Map2T.scala 17:7]
  assign O_8_2 = op_O_8_2; // @[Map2T.scala 17:7]
  assign O_9_0 = op_O_9_0; // @[Map2T.scala 17:7]
  assign O_9_1 = op_O_9_1; // @[Map2T.scala 17:7]
  assign O_9_2 = op_O_9_2; // @[Map2T.scala 17:7]
  assign O_10_0 = op_O_10_0; // @[Map2T.scala 17:7]
  assign O_10_1 = op_O_10_1; // @[Map2T.scala 17:7]
  assign O_10_2 = op_O_10_2; // @[Map2T.scala 17:7]
  assign O_11_0 = op_O_11_0; // @[Map2T.scala 17:7]
  assign O_11_1 = op_O_11_1; // @[Map2T.scala 17:7]
  assign O_11_2 = op_O_11_2; // @[Map2T.scala 17:7]
  assign O_12_0 = op_O_12_0; // @[Map2T.scala 17:7]
  assign O_12_1 = op_O_12_1; // @[Map2T.scala 17:7]
  assign O_12_2 = op_O_12_2; // @[Map2T.scala 17:7]
  assign O_13_0 = op_O_13_0; // @[Map2T.scala 17:7]
  assign O_13_1 = op_O_13_1; // @[Map2T.scala 17:7]
  assign O_13_2 = op_O_13_2; // @[Map2T.scala 17:7]
  assign O_14_0 = op_O_14_0; // @[Map2T.scala 17:7]
  assign O_14_1 = op_O_14_1; // @[Map2T.scala 17:7]
  assign O_14_2 = op_O_14_2; // @[Map2T.scala 17:7]
  assign O_15_0 = op_O_15_0; // @[Map2T.scala 17:7]
  assign O_15_1 = op_O_15_1; // @[Map2T.scala 17:7]
  assign O_15_2 = op_O_15_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  input  [31:0] I_3_0,
  input  [31:0] I_3_1,
  input  [31:0] I_3_2,
  input  [31:0] I_4_0,
  input  [31:0] I_4_1,
  input  [31:0] I_4_2,
  input  [31:0] I_5_0,
  input  [31:0] I_5_1,
  input  [31:0] I_5_2,
  input  [31:0] I_6_0,
  input  [31:0] I_6_1,
  input  [31:0] I_6_2,
  input  [31:0] I_7_0,
  input  [31:0] I_7_1,
  input  [31:0] I_7_2,
  input  [31:0] I_8_0,
  input  [31:0] I_8_1,
  input  [31:0] I_8_2,
  input  [31:0] I_9_0,
  input  [31:0] I_9_1,
  input  [31:0] I_9_2,
  input  [31:0] I_10_0,
  input  [31:0] I_10_1,
  input  [31:0] I_10_2,
  input  [31:0] I_11_0,
  input  [31:0] I_11_1,
  input  [31:0] I_11_2,
  input  [31:0] I_12_0,
  input  [31:0] I_12_1,
  input  [31:0] I_12_2,
  input  [31:0] I_13_0,
  input  [31:0] I_13_1,
  input  [31:0] I_13_2,
  input  [31:0] I_14_0,
  input  [31:0] I_14_1,
  input  [31:0] I_14_2,
  input  [31:0] I_15_0,
  input  [31:0] I_15_1,
  input  [31:0] I_15_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_4_0_2 = I_4_2; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_5_0_2 = I_5_2; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_6_0_2 = I_6_2; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_7_0_2 = I_7_2; // @[Partition.scala 15:39]
  assign O_8_0_0 = I_8_0; // @[Partition.scala 15:39]
  assign O_8_0_1 = I_8_1; // @[Partition.scala 15:39]
  assign O_8_0_2 = I_8_2; // @[Partition.scala 15:39]
  assign O_9_0_0 = I_9_0; // @[Partition.scala 15:39]
  assign O_9_0_1 = I_9_1; // @[Partition.scala 15:39]
  assign O_9_0_2 = I_9_2; // @[Partition.scala 15:39]
  assign O_10_0_0 = I_10_0; // @[Partition.scala 15:39]
  assign O_10_0_1 = I_10_1; // @[Partition.scala 15:39]
  assign O_10_0_2 = I_10_2; // @[Partition.scala 15:39]
  assign O_11_0_0 = I_11_0; // @[Partition.scala 15:39]
  assign O_11_0_1 = I_11_1; // @[Partition.scala 15:39]
  assign O_11_0_2 = I_11_2; // @[Partition.scala 15:39]
  assign O_12_0_0 = I_12_0; // @[Partition.scala 15:39]
  assign O_12_0_1 = I_12_1; // @[Partition.scala 15:39]
  assign O_12_0_2 = I_12_2; // @[Partition.scala 15:39]
  assign O_13_0_0 = I_13_0; // @[Partition.scala 15:39]
  assign O_13_0_1 = I_13_1; // @[Partition.scala 15:39]
  assign O_13_0_2 = I_13_2; // @[Partition.scala 15:39]
  assign O_14_0_0 = I_14_0; // @[Partition.scala 15:39]
  assign O_14_0_1 = I_14_1; // @[Partition.scala 15:39]
  assign O_14_0_2 = I_14_2; // @[Partition.scala 15:39]
  assign O_15_0_0 = I_15_0; // @[Partition.scala 15:39]
  assign O_15_0_1 = I_15_1; // @[Partition.scala 15:39]
  assign O_15_0_2 = I_15_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  input  [31:0] I_3_0,
  input  [31:0] I_3_1,
  input  [31:0] I_3_2,
  input  [31:0] I_4_0,
  input  [31:0] I_4_1,
  input  [31:0] I_4_2,
  input  [31:0] I_5_0,
  input  [31:0] I_5_1,
  input  [31:0] I_5_2,
  input  [31:0] I_6_0,
  input  [31:0] I_6_1,
  input  [31:0] I_6_2,
  input  [31:0] I_7_0,
  input  [31:0] I_7_1,
  input  [31:0] I_7_2,
  input  [31:0] I_8_0,
  input  [31:0] I_8_1,
  input  [31:0] I_8_2,
  input  [31:0] I_9_0,
  input  [31:0] I_9_1,
  input  [31:0] I_9_2,
  input  [31:0] I_10_0,
  input  [31:0] I_10_1,
  input  [31:0] I_10_2,
  input  [31:0] I_11_0,
  input  [31:0] I_11_1,
  input  [31:0] I_11_2,
  input  [31:0] I_12_0,
  input  [31:0] I_12_1,
  input  [31:0] I_12_2,
  input  [31:0] I_13_0,
  input  [31:0] I_13_1,
  input  [31:0] I_13_2,
  input  [31:0] I_14_0,
  input  [31:0] I_14_1,
  input  [31:0] I_14_2,
  input  [31:0] I_15_0,
  input  [31:0] I_15_1,
  input  [31:0] I_15_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_2_2(op_I_2_2),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_3_2(op_I_3_2),
    .I_4_0(op_I_4_0),
    .I_4_1(op_I_4_1),
    .I_4_2(op_I_4_2),
    .I_5_0(op_I_5_0),
    .I_5_1(op_I_5_1),
    .I_5_2(op_I_5_2),
    .I_6_0(op_I_6_0),
    .I_6_1(op_I_6_1),
    .I_6_2(op_I_6_2),
    .I_7_0(op_I_7_0),
    .I_7_1(op_I_7_1),
    .I_7_2(op_I_7_2),
    .I_8_0(op_I_8_0),
    .I_8_1(op_I_8_1),
    .I_8_2(op_I_8_2),
    .I_9_0(op_I_9_0),
    .I_9_1(op_I_9_1),
    .I_9_2(op_I_9_2),
    .I_10_0(op_I_10_0),
    .I_10_1(op_I_10_1),
    .I_10_2(op_I_10_2),
    .I_11_0(op_I_11_0),
    .I_11_1(op_I_11_1),
    .I_11_2(op_I_11_2),
    .I_12_0(op_I_12_0),
    .I_12_1(op_I_12_1),
    .I_12_2(op_I_12_2),
    .I_13_0(op_I_13_0),
    .I_13_1(op_I_13_1),
    .I_13_2(op_I_13_2),
    .I_14_0(op_I_14_0),
    .I_14_1(op_I_14_1),
    .I_14_2(op_I_14_2),
    .I_15_0(op_I_15_0),
    .I_15_1(op_I_15_1),
    .I_15_2(op_I_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2 = I_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_3_2 = I_3_2; // @[MapT.scala 14:10]
  assign op_I_4_0 = I_4_0; // @[MapT.scala 14:10]
  assign op_I_4_1 = I_4_1; // @[MapT.scala 14:10]
  assign op_I_4_2 = I_4_2; // @[MapT.scala 14:10]
  assign op_I_5_0 = I_5_0; // @[MapT.scala 14:10]
  assign op_I_5_1 = I_5_1; // @[MapT.scala 14:10]
  assign op_I_5_2 = I_5_2; // @[MapT.scala 14:10]
  assign op_I_6_0 = I_6_0; // @[MapT.scala 14:10]
  assign op_I_6_1 = I_6_1; // @[MapT.scala 14:10]
  assign op_I_6_2 = I_6_2; // @[MapT.scala 14:10]
  assign op_I_7_0 = I_7_0; // @[MapT.scala 14:10]
  assign op_I_7_1 = I_7_1; // @[MapT.scala 14:10]
  assign op_I_7_2 = I_7_2; // @[MapT.scala 14:10]
  assign op_I_8_0 = I_8_0; // @[MapT.scala 14:10]
  assign op_I_8_1 = I_8_1; // @[MapT.scala 14:10]
  assign op_I_8_2 = I_8_2; // @[MapT.scala 14:10]
  assign op_I_9_0 = I_9_0; // @[MapT.scala 14:10]
  assign op_I_9_1 = I_9_1; // @[MapT.scala 14:10]
  assign op_I_9_2 = I_9_2; // @[MapT.scala 14:10]
  assign op_I_10_0 = I_10_0; // @[MapT.scala 14:10]
  assign op_I_10_1 = I_10_1; // @[MapT.scala 14:10]
  assign op_I_10_2 = I_10_2; // @[MapT.scala 14:10]
  assign op_I_11_0 = I_11_0; // @[MapT.scala 14:10]
  assign op_I_11_1 = I_11_1; // @[MapT.scala 14:10]
  assign op_I_11_2 = I_11_2; // @[MapT.scala 14:10]
  assign op_I_12_0 = I_12_0; // @[MapT.scala 14:10]
  assign op_I_12_1 = I_12_1; // @[MapT.scala 14:10]
  assign op_I_12_2 = I_12_2; // @[MapT.scala 14:10]
  assign op_I_13_0 = I_13_0; // @[MapT.scala 14:10]
  assign op_I_13_1 = I_13_1; // @[MapT.scala 14:10]
  assign op_I_13_2 = I_13_2; // @[MapT.scala 14:10]
  assign op_I_14_0 = I_14_0; // @[MapT.scala 14:10]
  assign op_I_14_1 = I_14_1; // @[MapT.scala 14:10]
  assign op_I_14_2 = I_14_2; // @[MapT.scala 14:10]
  assign op_I_15_0 = I_15_0; // @[MapT.scala 14:10]
  assign op_I_15_1 = I_15_1; // @[MapT.scala 14:10]
  assign op_I_15_2 = I_15_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2,
  output [31:0] O_8_0,
  output [31:0] O_8_1,
  output [31:0] O_8_2,
  output [31:0] O_9_0,
  output [31:0] O_9_1,
  output [31:0] O_9_2,
  output [31:0] O_10_0,
  output [31:0] O_10_1,
  output [31:0] O_10_2,
  output [31:0] O_11_0,
  output [31:0] O_11_1,
  output [31:0] O_11_2,
  output [31:0] O_12_0,
  output [31:0] O_12_1,
  output [31:0] O_12_2,
  output [31:0] O_13_0,
  output [31:0] O_13_1,
  output [31:0] O_13_2,
  output [31:0] O_14_0,
  output [31:0] O_14_1,
  output [31:0] O_14_2,
  output [31:0] O_15_0,
  output [31:0] O_15_1,
  output [31:0] O_15_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  Remove1S other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  Remove1S other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  Remove1S other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  Remove1S other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  Remove1S other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  Remove1S other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  Remove1S other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  Remove1S other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  Remove1S other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  Remove1S other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  Remove1S other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  Remove1S other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_4_2 = other_ops_3_O_2; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_5_2 = other_ops_4_O_2; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_6_2 = other_ops_5_O_2; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_7_2 = other_ops_6_O_2; // @[MapS.scala 21:12]
  assign O_8_0 = other_ops_7_O_0; // @[MapS.scala 21:12]
  assign O_8_1 = other_ops_7_O_1; // @[MapS.scala 21:12]
  assign O_8_2 = other_ops_7_O_2; // @[MapS.scala 21:12]
  assign O_9_0 = other_ops_8_O_0; // @[MapS.scala 21:12]
  assign O_9_1 = other_ops_8_O_1; // @[MapS.scala 21:12]
  assign O_9_2 = other_ops_8_O_2; // @[MapS.scala 21:12]
  assign O_10_0 = other_ops_9_O_0; // @[MapS.scala 21:12]
  assign O_10_1 = other_ops_9_O_1; // @[MapS.scala 21:12]
  assign O_10_2 = other_ops_9_O_2; // @[MapS.scala 21:12]
  assign O_11_0 = other_ops_10_O_0; // @[MapS.scala 21:12]
  assign O_11_1 = other_ops_10_O_1; // @[MapS.scala 21:12]
  assign O_11_2 = other_ops_10_O_2; // @[MapS.scala 21:12]
  assign O_12_0 = other_ops_11_O_0; // @[MapS.scala 21:12]
  assign O_12_1 = other_ops_11_O_1; // @[MapS.scala 21:12]
  assign O_12_2 = other_ops_11_O_2; // @[MapS.scala 21:12]
  assign O_13_0 = other_ops_12_O_0; // @[MapS.scala 21:12]
  assign O_13_1 = other_ops_12_O_1; // @[MapS.scala 21:12]
  assign O_13_2 = other_ops_12_O_2; // @[MapS.scala 21:12]
  assign O_14_0 = other_ops_13_O_0; // @[MapS.scala 21:12]
  assign O_14_1 = other_ops_13_O_1; // @[MapS.scala 21:12]
  assign O_14_2 = other_ops_13_O_2; // @[MapS.scala 21:12]
  assign O_15_0 = other_ops_14_O_0; // @[MapS.scala 21:12]
  assign O_15_1 = other_ops_14_O_1; // @[MapS.scala 21:12]
  assign O_15_2 = other_ops_14_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2,
  output [31:0] O_3_0,
  output [31:0] O_3_1,
  output [31:0] O_3_2,
  output [31:0] O_4_0,
  output [31:0] O_4_1,
  output [31:0] O_4_2,
  output [31:0] O_5_0,
  output [31:0] O_5_1,
  output [31:0] O_5_2,
  output [31:0] O_6_0,
  output [31:0] O_6_1,
  output [31:0] O_6_2,
  output [31:0] O_7_0,
  output [31:0] O_7_1,
  output [31:0] O_7_2,
  output [31:0] O_8_0,
  output [31:0] O_8_1,
  output [31:0] O_8_2,
  output [31:0] O_9_0,
  output [31:0] O_9_1,
  output [31:0] O_9_2,
  output [31:0] O_10_0,
  output [31:0] O_10_1,
  output [31:0] O_10_2,
  output [31:0] O_11_0,
  output [31:0] O_11_1,
  output [31:0] O_11_2,
  output [31:0] O_12_0,
  output [31:0] O_12_1,
  output [31:0] O_12_2,
  output [31:0] O_13_0,
  output [31:0] O_13_1,
  output [31:0] O_13_2,
  output [31:0] O_14_0,
  output [31:0] O_14_1,
  output [31:0] O_14_2,
  output [31:0] O_15_0,
  output [31:0] O_15_1,
  output [31:0] O_15_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_8_2(op_O_8_2),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_9_2(op_O_9_2),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_10_2(op_O_10_2),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_11_2(op_O_11_2),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_12_2(op_O_12_2),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_13_2(op_O_13_2),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_14_2(op_O_14_2),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1),
    .O_15_2(op_O_15_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_2_2 = op_O_2_2; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_3_2 = op_O_3_2; // @[MapT.scala 15:7]
  assign O_4_0 = op_O_4_0; // @[MapT.scala 15:7]
  assign O_4_1 = op_O_4_1; // @[MapT.scala 15:7]
  assign O_4_2 = op_O_4_2; // @[MapT.scala 15:7]
  assign O_5_0 = op_O_5_0; // @[MapT.scala 15:7]
  assign O_5_1 = op_O_5_1; // @[MapT.scala 15:7]
  assign O_5_2 = op_O_5_2; // @[MapT.scala 15:7]
  assign O_6_0 = op_O_6_0; // @[MapT.scala 15:7]
  assign O_6_1 = op_O_6_1; // @[MapT.scala 15:7]
  assign O_6_2 = op_O_6_2; // @[MapT.scala 15:7]
  assign O_7_0 = op_O_7_0; // @[MapT.scala 15:7]
  assign O_7_1 = op_O_7_1; // @[MapT.scala 15:7]
  assign O_7_2 = op_O_7_2; // @[MapT.scala 15:7]
  assign O_8_0 = op_O_8_0; // @[MapT.scala 15:7]
  assign O_8_1 = op_O_8_1; // @[MapT.scala 15:7]
  assign O_8_2 = op_O_8_2; // @[MapT.scala 15:7]
  assign O_9_0 = op_O_9_0; // @[MapT.scala 15:7]
  assign O_9_1 = op_O_9_1; // @[MapT.scala 15:7]
  assign O_9_2 = op_O_9_2; // @[MapT.scala 15:7]
  assign O_10_0 = op_O_10_0; // @[MapT.scala 15:7]
  assign O_10_1 = op_O_10_1; // @[MapT.scala 15:7]
  assign O_10_2 = op_O_10_2; // @[MapT.scala 15:7]
  assign O_11_0 = op_O_11_0; // @[MapT.scala 15:7]
  assign O_11_1 = op_O_11_1; // @[MapT.scala 15:7]
  assign O_11_2 = op_O_11_2; // @[MapT.scala 15:7]
  assign O_12_0 = op_O_12_0; // @[MapT.scala 15:7]
  assign O_12_1 = op_O_12_1; // @[MapT.scala 15:7]
  assign O_12_2 = op_O_12_2; // @[MapT.scala 15:7]
  assign O_13_0 = op_O_13_0; // @[MapT.scala 15:7]
  assign O_13_1 = op_O_13_1; // @[MapT.scala 15:7]
  assign O_13_2 = op_O_13_2; // @[MapT.scala 15:7]
  assign O_14_0 = op_O_14_0; // @[MapT.scala 15:7]
  assign O_14_1 = op_O_14_1; // @[MapT.scala 15:7]
  assign O_14_2 = op_O_14_2; // @[MapT.scala 15:7]
  assign O_15_0 = op_O_15_0; // @[MapT.scala 15:7]
  assign O_15_1 = op_O_15_1; // @[MapT.scala 15:7]
  assign O_15_2 = op_O_15_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_3_2,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_4_2,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_5_2,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_6_2,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I0_7_2,
  input  [31:0] I0_8_0,
  input  [31:0] I0_8_1,
  input  [31:0] I0_8_2,
  input  [31:0] I0_9_0,
  input  [31:0] I0_9_1,
  input  [31:0] I0_9_2,
  input  [31:0] I0_10_0,
  input  [31:0] I0_10_1,
  input  [31:0] I0_10_2,
  input  [31:0] I0_11_0,
  input  [31:0] I0_11_1,
  input  [31:0] I0_11_2,
  input  [31:0] I0_12_0,
  input  [31:0] I0_12_1,
  input  [31:0] I0_12_2,
  input  [31:0] I0_13_0,
  input  [31:0] I0_13_1,
  input  [31:0] I0_13_2,
  input  [31:0] I0_14_0,
  input  [31:0] I0_14_1,
  input  [31:0] I0_14_2,
  input  [31:0] I0_15_0,
  input  [31:0] I0_15_1,
  input  [31:0] I0_15_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  input  [31:0] I1_8_0,
  input  [31:0] I1_8_1,
  input  [31:0] I1_8_2,
  input  [31:0] I1_9_0,
  input  [31:0] I1_9_1,
  input  [31:0] I1_9_2,
  input  [31:0] I1_10_0,
  input  [31:0] I1_10_1,
  input  [31:0] I1_10_2,
  input  [31:0] I1_11_0,
  input  [31:0] I1_11_1,
  input  [31:0] I1_11_2,
  input  [31:0] I1_12_0,
  input  [31:0] I1_12_1,
  input  [31:0] I1_12_2,
  input  [31:0] I1_13_0,
  input  [31:0] I1_13_1,
  input  [31:0] I1_13_2,
  input  [31:0] I1_14_0,
  input  [31:0] I1_14_1,
  input  [31:0] I1_14_2,
  input  [31:0] I1_15_0,
  input  [31:0] I1_15_1,
  input  [31:0] I1_15_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I0_2(other_ops_3_I0_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I0_2(other_ops_4_I0_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I0_2(other_ops_5_I0_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I0_2(other_ops_6_I0_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I0_2(other_ops_7_I0_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I0_2(other_ops_8_I0_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I0_2(other_ops_9_I0_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I0_2(other_ops_10_I0_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I0_2(other_ops_11_I0_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I0_2(other_ops_12_I0_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I0_2(other_ops_13_I0_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I0_2(other_ops_14_I0_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2 = I0_4_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2 = I0_5_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2 = I0_6_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2 = I0_7_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2 = I0_8_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2 = I0_9_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2 = I0_10_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2 = I0_11_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2 = I0_12_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2 = I0_13_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2 = I0_14_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2 = I0_15_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  input  [31:0] I0_3_0,
  input  [31:0] I0_3_1,
  input  [31:0] I0_3_2,
  input  [31:0] I0_4_0,
  input  [31:0] I0_4_1,
  input  [31:0] I0_4_2,
  input  [31:0] I0_5_0,
  input  [31:0] I0_5_1,
  input  [31:0] I0_5_2,
  input  [31:0] I0_6_0,
  input  [31:0] I0_6_1,
  input  [31:0] I0_6_2,
  input  [31:0] I0_7_0,
  input  [31:0] I0_7_1,
  input  [31:0] I0_7_2,
  input  [31:0] I0_8_0,
  input  [31:0] I0_8_1,
  input  [31:0] I0_8_2,
  input  [31:0] I0_9_0,
  input  [31:0] I0_9_1,
  input  [31:0] I0_9_2,
  input  [31:0] I0_10_0,
  input  [31:0] I0_10_1,
  input  [31:0] I0_10_2,
  input  [31:0] I0_11_0,
  input  [31:0] I0_11_1,
  input  [31:0] I0_11_2,
  input  [31:0] I0_12_0,
  input  [31:0] I0_12_1,
  input  [31:0] I0_12_2,
  input  [31:0] I0_13_0,
  input  [31:0] I0_13_1,
  input  [31:0] I0_13_2,
  input  [31:0] I0_14_0,
  input  [31:0] I0_14_1,
  input  [31:0] I0_14_2,
  input  [31:0] I0_15_0,
  input  [31:0] I0_15_1,
  input  [31:0] I0_15_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  input  [31:0] I1_8_0,
  input  [31:0] I1_8_1,
  input  [31:0] I1_8_2,
  input  [31:0] I1_9_0,
  input  [31:0] I1_9_1,
  input  [31:0] I1_9_2,
  input  [31:0] I1_10_0,
  input  [31:0] I1_10_1,
  input  [31:0] I1_10_2,
  input  [31:0] I1_11_0,
  input  [31:0] I1_11_1,
  input  [31:0] I1_11_2,
  input  [31:0] I1_12_0,
  input  [31:0] I1_12_1,
  input  [31:0] I1_12_2,
  input  [31:0] I1_13_0,
  input  [31:0] I1_13_1,
  input  [31:0] I1_13_2,
  input  [31:0] I1_14_0,
  input  [31:0] I1_14_1,
  input  [31:0] I1_14_2,
  input  [31:0] I1_15_0,
  input  [31:0] I1_15_1,
  input  [31:0] I1_15_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_2_2(op_I0_2_2),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_3_2(op_I0_3_2),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_4_2(op_I0_4_2),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_5_2(op_I0_5_2),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_6_2(op_I0_6_2),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_7_2(op_I0_7_2),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_8_2(op_I0_8_2),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_9_2(op_I0_9_2),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_10_2(op_I0_10_2),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_11_2(op_I0_11_2),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_12_2(op_I0_12_2),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_13_2(op_I0_13_2),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_14_2(op_I0_14_2),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I0_15_2(op_I0_15_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_8_2(op_I1_8_2),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_9_2(op_I1_9_2),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_10_2(op_I1_10_2),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_11_2(op_I1_11_2),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_12_2(op_I1_12_2),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_13_2(op_I1_13_2),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_14_2(op_I1_14_2),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .I1_15_2(op_I1_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_2 = op_O_8_0_2; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_8_1_2 = op_O_8_1_2; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_2 = op_O_9_0_2; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_9_1_2 = op_O_9_1_2; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_2 = op_O_10_0_2; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_10_1_2 = op_O_10_1_2; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_2 = op_O_11_0_2; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_11_1_2 = op_O_11_1_2; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_2 = op_O_12_0_2; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_12_1_2 = op_O_12_1_2; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_2 = op_O_13_0_2; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_13_1_2 = op_O_13_1_2; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_2 = op_O_14_0_2; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_14_1_2 = op_O_14_1_2; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_2 = op_O_15_0_2; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign O_15_1_2 = op_O_15_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2 = I0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2 = I0_3_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2 = I0_4_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2 = I0_5_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2 = I0_6_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2 = I0_7_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_8_2 = I0_8_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_9_2 = I0_9_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_10_2 = I0_10_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_11_2 = I0_11_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_12_2 = I0_12_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_13_2 = I0_13_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_14_2 = I0_14_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I0_15_2 = I0_15_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_8_2 = I1_8_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_9_2 = I1_9_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_10_2 = I1_10_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_11_2 = I1_11_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_12_2 = I1_12_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_13_2 = I1_13_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_14_2 = I1_14_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
  assign op_I1_15_2 = I1_15_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I1_0,
  input  [31:0] I1_1,
  input  [31:0] I1_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I0_8_0_0,
  input  [31:0] I0_8_0_1,
  input  [31:0] I0_8_0_2,
  input  [31:0] I0_8_1_0,
  input  [31:0] I0_8_1_1,
  input  [31:0] I0_8_1_2,
  input  [31:0] I0_9_0_0,
  input  [31:0] I0_9_0_1,
  input  [31:0] I0_9_0_2,
  input  [31:0] I0_9_1_0,
  input  [31:0] I0_9_1_1,
  input  [31:0] I0_9_1_2,
  input  [31:0] I0_10_0_0,
  input  [31:0] I0_10_0_1,
  input  [31:0] I0_10_0_2,
  input  [31:0] I0_10_1_0,
  input  [31:0] I0_10_1_1,
  input  [31:0] I0_10_1_2,
  input  [31:0] I0_11_0_0,
  input  [31:0] I0_11_0_1,
  input  [31:0] I0_11_0_2,
  input  [31:0] I0_11_1_0,
  input  [31:0] I0_11_1_1,
  input  [31:0] I0_11_1_2,
  input  [31:0] I0_12_0_0,
  input  [31:0] I0_12_0_1,
  input  [31:0] I0_12_0_2,
  input  [31:0] I0_12_1_0,
  input  [31:0] I0_12_1_1,
  input  [31:0] I0_12_1_2,
  input  [31:0] I0_13_0_0,
  input  [31:0] I0_13_0_1,
  input  [31:0] I0_13_0_2,
  input  [31:0] I0_13_1_0,
  input  [31:0] I0_13_1_1,
  input  [31:0] I0_13_1_2,
  input  [31:0] I0_14_0_0,
  input  [31:0] I0_14_0_1,
  input  [31:0] I0_14_0_2,
  input  [31:0] I0_14_1_0,
  input  [31:0] I0_14_1_1,
  input  [31:0] I0_14_1_2,
  input  [31:0] I0_15_0_0,
  input  [31:0] I0_15_0_1,
  input  [31:0] I0_15_0_2,
  input  [31:0] I0_15_1_0,
  input  [31:0] I0_15_1_1,
  input  [31:0] I0_15_1_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  input  [31:0] I1_8_0,
  input  [31:0] I1_8_1,
  input  [31:0] I1_8_2,
  input  [31:0] I1_9_0,
  input  [31:0] I1_9_1,
  input  [31:0] I1_9_2,
  input  [31:0] I1_10_0,
  input  [31:0] I1_10_1,
  input  [31:0] I1_10_2,
  input  [31:0] I1_11_0,
  input  [31:0] I1_11_1,
  input  [31:0] I1_11_2,
  input  [31:0] I1_12_0,
  input  [31:0] I1_12_1,
  input  [31:0] I1_12_2,
  input  [31:0] I1_13_0,
  input  [31:0] I1_13_1,
  input  [31:0] I1_13_2,
  input  [31:0] I1_14_0,
  input  [31:0] I1_14_1,
  input  [31:0] I1_14_2,
  input  [31:0] I1_15_0,
  input  [31:0] I1_15_1,
  input  [31:0] I1_15_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_8_2_0,
  output [31:0] O_8_2_1,
  output [31:0] O_8_2_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_9_2_0,
  output [31:0] O_9_2_1,
  output [31:0] O_9_2_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_10_2_0,
  output [31:0] O_10_2_1,
  output [31:0] O_10_2_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_11_2_0,
  output [31:0] O_11_2_1,
  output [31:0] O_11_2_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_12_2_0,
  output [31:0] O_12_2_1,
  output [31:0] O_12_2_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_13_2_0,
  output [31:0] O_13_2_1,
  output [31:0] O_13_2_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_14_2_0,
  output [31:0] O_14_2_1,
  output [31:0] O_14_2_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2,
  output [31:0] O_15_2_0,
  output [31:0] O_15_2_1,
  output [31:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I0_0_1(other_ops_7_I0_0_1),
    .I0_0_2(other_ops_7_I0_0_2),
    .I0_1_0(other_ops_7_I0_1_0),
    .I0_1_1(other_ops_7_I0_1_1),
    .I0_1_2(other_ops_7_I0_1_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I0_0_1(other_ops_8_I0_0_1),
    .I0_0_2(other_ops_8_I0_0_2),
    .I0_1_0(other_ops_8_I0_1_0),
    .I0_1_1(other_ops_8_I0_1_1),
    .I0_1_2(other_ops_8_I0_1_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I0_0_1(other_ops_9_I0_0_1),
    .I0_0_2(other_ops_9_I0_0_2),
    .I0_1_0(other_ops_9_I0_1_0),
    .I0_1_1(other_ops_9_I0_1_1),
    .I0_1_2(other_ops_9_I0_1_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I0_0_1(other_ops_10_I0_0_1),
    .I0_0_2(other_ops_10_I0_0_2),
    .I0_1_0(other_ops_10_I0_1_0),
    .I0_1_1(other_ops_10_I0_1_1),
    .I0_1_2(other_ops_10_I0_1_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I0_0_1(other_ops_11_I0_0_1),
    .I0_0_2(other_ops_11_I0_0_2),
    .I0_1_0(other_ops_11_I0_1_0),
    .I0_1_1(other_ops_11_I0_1_1),
    .I0_1_2(other_ops_11_I0_1_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I0_0_1(other_ops_12_I0_0_1),
    .I0_0_2(other_ops_12_I0_0_2),
    .I0_1_0(other_ops_12_I0_1_0),
    .I0_1_1(other_ops_12_I0_1_1),
    .I0_1_2(other_ops_12_I0_1_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I0_0_1(other_ops_13_I0_0_1),
    .I0_0_2(other_ops_13_I0_0_2),
    .I0_1_0(other_ops_13_I0_1_0),
    .I0_1_1(other_ops_13_I0_1_1),
    .I0_1_2(other_ops_13_I0_1_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I0_0_1(other_ops_14_I0_0_1),
    .I0_0_2(other_ops_14_I0_0_2),
    .I0_1_0(other_ops_14_I0_1_0),
    .I0_1_1(other_ops_14_I0_1_1),
    .I0_1_2(other_ops_14_I0_1_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[Map2S.scala 24:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[Map2S.scala 24:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[Map2S.scala 24:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[Map2S.scala 24:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[Map2S.scala 24:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[Map2S.scala 24:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[Map2S.scala 24:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[Map2S.scala 24:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[Map2S.scala 24:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[Map2S.scala 24:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[Map2S.scala 24:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[Map2S.scala 24:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[Map2S.scala 24:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[Map2S.scala 24:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[Map2S.scala 24:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[Map2S.scala 24:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[Map2S.scala 24:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[Map2S.scala 24:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[Map2S.scala 24:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[Map2S.scala 24:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[Map2S.scala 24:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[Map2S.scala 24:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[Map2S.scala 24:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[Map2S.scala 24:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1 = I0_8_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_2 = I0_8_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_0 = I0_8_1_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_1 = I0_8_1_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_2 = I0_8_1_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1 = I0_9_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_2 = I0_9_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_0 = I0_9_1_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_1 = I0_9_1_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_2 = I0_9_1_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1 = I0_10_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_2 = I0_10_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_0 = I0_10_1_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_1 = I0_10_1_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_2 = I0_10_1_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1 = I0_11_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_2 = I0_11_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_0 = I0_11_1_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_1 = I0_11_1_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_2 = I0_11_1_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1 = I0_12_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_2 = I0_12_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_0 = I0_12_1_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_1 = I0_12_1_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_2 = I0_12_1_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1 = I0_13_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_2 = I0_13_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_0 = I0_13_1_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_1 = I0_13_1_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_2 = I0_13_1_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1 = I0_14_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_2 = I0_14_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_0 = I0_14_1_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_1 = I0_14_1_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_2 = I0_14_1_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1 = I0_15_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_2 = I0_15_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_0 = I0_15_1_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_1 = I0_15_1_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_2 = I0_15_1_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I0_8_0_0,
  input  [31:0] I0_8_0_1,
  input  [31:0] I0_8_0_2,
  input  [31:0] I0_8_1_0,
  input  [31:0] I0_8_1_1,
  input  [31:0] I0_8_1_2,
  input  [31:0] I0_9_0_0,
  input  [31:0] I0_9_0_1,
  input  [31:0] I0_9_0_2,
  input  [31:0] I0_9_1_0,
  input  [31:0] I0_9_1_1,
  input  [31:0] I0_9_1_2,
  input  [31:0] I0_10_0_0,
  input  [31:0] I0_10_0_1,
  input  [31:0] I0_10_0_2,
  input  [31:0] I0_10_1_0,
  input  [31:0] I0_10_1_1,
  input  [31:0] I0_10_1_2,
  input  [31:0] I0_11_0_0,
  input  [31:0] I0_11_0_1,
  input  [31:0] I0_11_0_2,
  input  [31:0] I0_11_1_0,
  input  [31:0] I0_11_1_1,
  input  [31:0] I0_11_1_2,
  input  [31:0] I0_12_0_0,
  input  [31:0] I0_12_0_1,
  input  [31:0] I0_12_0_2,
  input  [31:0] I0_12_1_0,
  input  [31:0] I0_12_1_1,
  input  [31:0] I0_12_1_2,
  input  [31:0] I0_13_0_0,
  input  [31:0] I0_13_0_1,
  input  [31:0] I0_13_0_2,
  input  [31:0] I0_13_1_0,
  input  [31:0] I0_13_1_1,
  input  [31:0] I0_13_1_2,
  input  [31:0] I0_14_0_0,
  input  [31:0] I0_14_0_1,
  input  [31:0] I0_14_0_2,
  input  [31:0] I0_14_1_0,
  input  [31:0] I0_14_1_1,
  input  [31:0] I0_14_1_2,
  input  [31:0] I0_15_0_0,
  input  [31:0] I0_15_0_1,
  input  [31:0] I0_15_0_2,
  input  [31:0] I0_15_1_0,
  input  [31:0] I0_15_1_1,
  input  [31:0] I0_15_1_2,
  input  [31:0] I1_0_0,
  input  [31:0] I1_0_1,
  input  [31:0] I1_0_2,
  input  [31:0] I1_1_0,
  input  [31:0] I1_1_1,
  input  [31:0] I1_1_2,
  input  [31:0] I1_2_0,
  input  [31:0] I1_2_1,
  input  [31:0] I1_2_2,
  input  [31:0] I1_3_0,
  input  [31:0] I1_3_1,
  input  [31:0] I1_3_2,
  input  [31:0] I1_4_0,
  input  [31:0] I1_4_1,
  input  [31:0] I1_4_2,
  input  [31:0] I1_5_0,
  input  [31:0] I1_5_1,
  input  [31:0] I1_5_2,
  input  [31:0] I1_6_0,
  input  [31:0] I1_6_1,
  input  [31:0] I1_6_2,
  input  [31:0] I1_7_0,
  input  [31:0] I1_7_1,
  input  [31:0] I1_7_2,
  input  [31:0] I1_8_0,
  input  [31:0] I1_8_1,
  input  [31:0] I1_8_2,
  input  [31:0] I1_9_0,
  input  [31:0] I1_9_1,
  input  [31:0] I1_9_2,
  input  [31:0] I1_10_0,
  input  [31:0] I1_10_1,
  input  [31:0] I1_10_2,
  input  [31:0] I1_11_0,
  input  [31:0] I1_11_1,
  input  [31:0] I1_11_2,
  input  [31:0] I1_12_0,
  input  [31:0] I1_12_1,
  input  [31:0] I1_12_2,
  input  [31:0] I1_13_0,
  input  [31:0] I1_13_1,
  input  [31:0] I1_13_2,
  input  [31:0] I1_14_0,
  input  [31:0] I1_14_1,
  input  [31:0] I1_14_2,
  input  [31:0] I1_15_0,
  input  [31:0] I1_15_1,
  input  [31:0] I1_15_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_8_2_0,
  output [31:0] O_8_2_1,
  output [31:0] O_8_2_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_9_2_0,
  output [31:0] O_9_2_1,
  output [31:0] O_9_2_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_10_2_0,
  output [31:0] O_10_2_1,
  output [31:0] O_10_2_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_11_2_0,
  output [31:0] O_11_2_1,
  output [31:0] O_11_2_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_12_2_0,
  output [31:0] O_12_2_1,
  output [31:0] O_12_2_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_13_2_0,
  output [31:0] O_13_2_1,
  output [31:0] O_13_2_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_14_2_0,
  output [31:0] O_14_2_1,
  output [31:0] O_14_2_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2,
  output [31:0] O_15_2_0,
  output [31:0] O_15_2_1,
  output [31:0] O_15_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_8_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_9_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_10_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_11_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_12_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_13_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_14_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I1_15_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_8_0_1(op_I0_8_0_1),
    .I0_8_0_2(op_I0_8_0_2),
    .I0_8_1_0(op_I0_8_1_0),
    .I0_8_1_1(op_I0_8_1_1),
    .I0_8_1_2(op_I0_8_1_2),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_9_0_1(op_I0_9_0_1),
    .I0_9_0_2(op_I0_9_0_2),
    .I0_9_1_0(op_I0_9_1_0),
    .I0_9_1_1(op_I0_9_1_1),
    .I0_9_1_2(op_I0_9_1_2),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_10_0_1(op_I0_10_0_1),
    .I0_10_0_2(op_I0_10_0_2),
    .I0_10_1_0(op_I0_10_1_0),
    .I0_10_1_1(op_I0_10_1_1),
    .I0_10_1_2(op_I0_10_1_2),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_11_0_1(op_I0_11_0_1),
    .I0_11_0_2(op_I0_11_0_2),
    .I0_11_1_0(op_I0_11_1_0),
    .I0_11_1_1(op_I0_11_1_1),
    .I0_11_1_2(op_I0_11_1_2),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_12_0_1(op_I0_12_0_1),
    .I0_12_0_2(op_I0_12_0_2),
    .I0_12_1_0(op_I0_12_1_0),
    .I0_12_1_1(op_I0_12_1_1),
    .I0_12_1_2(op_I0_12_1_2),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_13_0_1(op_I0_13_0_1),
    .I0_13_0_2(op_I0_13_0_2),
    .I0_13_1_0(op_I0_13_1_0),
    .I0_13_1_1(op_I0_13_1_1),
    .I0_13_1_2(op_I0_13_1_2),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_14_0_1(op_I0_14_0_1),
    .I0_14_0_2(op_I0_14_0_2),
    .I0_14_1_0(op_I0_14_1_0),
    .I0_14_1_1(op_I0_14_1_1),
    .I0_14_1_2(op_I0_14_1_2),
    .I0_15_0_0(op_I0_15_0_0),
    .I0_15_0_1(op_I0_15_0_1),
    .I0_15_0_2(op_I0_15_0_2),
    .I0_15_1_0(op_I0_15_1_0),
    .I0_15_1_1(op_I0_15_1_1),
    .I0_15_1_2(op_I0_15_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_8_2(op_I1_8_2),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_9_2(op_I1_9_2),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_10_2(op_I1_10_2),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_11_2(op_I1_11_2),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_12_2(op_I1_12_2),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_13_2(op_I1_13_2),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_14_2(op_I1_14_2),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .I1_15_2(op_I1_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_2_2_0 = op_O_2_2_0; // @[Map2T.scala 17:7]
  assign O_2_2_1 = op_O_2_2_1; // @[Map2T.scala 17:7]
  assign O_2_2_2 = op_O_2_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_3_2_0 = op_O_3_2_0; // @[Map2T.scala 17:7]
  assign O_3_2_1 = op_O_3_2_1; // @[Map2T.scala 17:7]
  assign O_3_2_2 = op_O_3_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_4_2_0 = op_O_4_2_0; // @[Map2T.scala 17:7]
  assign O_4_2_1 = op_O_4_2_1; // @[Map2T.scala 17:7]
  assign O_4_2_2 = op_O_4_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_5_2_0 = op_O_5_2_0; // @[Map2T.scala 17:7]
  assign O_5_2_1 = op_O_5_2_1; // @[Map2T.scala 17:7]
  assign O_5_2_2 = op_O_5_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_6_2_0 = op_O_6_2_0; // @[Map2T.scala 17:7]
  assign O_6_2_1 = op_O_6_2_1; // @[Map2T.scala 17:7]
  assign O_6_2_2 = op_O_6_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_7_2_0 = op_O_7_2_0; // @[Map2T.scala 17:7]
  assign O_7_2_1 = op_O_7_2_1; // @[Map2T.scala 17:7]
  assign O_7_2_2 = op_O_7_2_2; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_2 = op_O_8_0_2; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_8_1_2 = op_O_8_1_2; // @[Map2T.scala 17:7]
  assign O_8_2_0 = op_O_8_2_0; // @[Map2T.scala 17:7]
  assign O_8_2_1 = op_O_8_2_1; // @[Map2T.scala 17:7]
  assign O_8_2_2 = op_O_8_2_2; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_2 = op_O_9_0_2; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_9_1_2 = op_O_9_1_2; // @[Map2T.scala 17:7]
  assign O_9_2_0 = op_O_9_2_0; // @[Map2T.scala 17:7]
  assign O_9_2_1 = op_O_9_2_1; // @[Map2T.scala 17:7]
  assign O_9_2_2 = op_O_9_2_2; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_2 = op_O_10_0_2; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_10_1_2 = op_O_10_1_2; // @[Map2T.scala 17:7]
  assign O_10_2_0 = op_O_10_2_0; // @[Map2T.scala 17:7]
  assign O_10_2_1 = op_O_10_2_1; // @[Map2T.scala 17:7]
  assign O_10_2_2 = op_O_10_2_2; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_2 = op_O_11_0_2; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_11_1_2 = op_O_11_1_2; // @[Map2T.scala 17:7]
  assign O_11_2_0 = op_O_11_2_0; // @[Map2T.scala 17:7]
  assign O_11_2_1 = op_O_11_2_1; // @[Map2T.scala 17:7]
  assign O_11_2_2 = op_O_11_2_2; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_2 = op_O_12_0_2; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_12_1_2 = op_O_12_1_2; // @[Map2T.scala 17:7]
  assign O_12_2_0 = op_O_12_2_0; // @[Map2T.scala 17:7]
  assign O_12_2_1 = op_O_12_2_1; // @[Map2T.scala 17:7]
  assign O_12_2_2 = op_O_12_2_2; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_2 = op_O_13_0_2; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_13_1_2 = op_O_13_1_2; // @[Map2T.scala 17:7]
  assign O_13_2_0 = op_O_13_2_0; // @[Map2T.scala 17:7]
  assign O_13_2_1 = op_O_13_2_1; // @[Map2T.scala 17:7]
  assign O_13_2_2 = op_O_13_2_2; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_2 = op_O_14_0_2; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_14_1_2 = op_O_14_1_2; // @[Map2T.scala 17:7]
  assign O_14_2_0 = op_O_14_2_0; // @[Map2T.scala 17:7]
  assign O_14_2_1 = op_O_14_2_1; // @[Map2T.scala 17:7]
  assign O_14_2_2 = op_O_14_2_2; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_2 = op_O_15_0_2; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign O_15_1_2 = op_O_15_1_2; // @[Map2T.scala 17:7]
  assign O_15_2_0 = op_O_15_2_0; // @[Map2T.scala 17:7]
  assign O_15_2_1 = op_O_15_2_1; // @[Map2T.scala 17:7]
  assign O_15_2_2 = op_O_15_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1 = I0_8_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_2 = I0_8_0_2; // @[Map2T.scala 15:11]
  assign op_I0_8_1_0 = I0_8_1_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1_1 = I0_8_1_1; // @[Map2T.scala 15:11]
  assign op_I0_8_1_2 = I0_8_1_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1 = I0_9_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_2 = I0_9_0_2; // @[Map2T.scala 15:11]
  assign op_I0_9_1_0 = I0_9_1_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1_1 = I0_9_1_1; // @[Map2T.scala 15:11]
  assign op_I0_9_1_2 = I0_9_1_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1 = I0_10_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_2 = I0_10_0_2; // @[Map2T.scala 15:11]
  assign op_I0_10_1_0 = I0_10_1_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1_1 = I0_10_1_1; // @[Map2T.scala 15:11]
  assign op_I0_10_1_2 = I0_10_1_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1 = I0_11_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_2 = I0_11_0_2; // @[Map2T.scala 15:11]
  assign op_I0_11_1_0 = I0_11_1_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1_1 = I0_11_1_1; // @[Map2T.scala 15:11]
  assign op_I0_11_1_2 = I0_11_1_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1 = I0_12_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_2 = I0_12_0_2; // @[Map2T.scala 15:11]
  assign op_I0_12_1_0 = I0_12_1_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1_1 = I0_12_1_1; // @[Map2T.scala 15:11]
  assign op_I0_12_1_2 = I0_12_1_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1 = I0_13_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_2 = I0_13_0_2; // @[Map2T.scala 15:11]
  assign op_I0_13_1_0 = I0_13_1_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1_1 = I0_13_1_1; // @[Map2T.scala 15:11]
  assign op_I0_13_1_2 = I0_13_1_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1 = I0_14_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_2 = I0_14_0_2; // @[Map2T.scala 15:11]
  assign op_I0_14_1_0 = I0_14_1_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1_1 = I0_14_1_1; // @[Map2T.scala 15:11]
  assign op_I0_14_1_2 = I0_14_1_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1 = I0_15_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_2 = I0_15_0_2; // @[Map2T.scala 15:11]
  assign op_I0_15_1_0 = I0_15_1_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1_1 = I0_15_1_1; // @[Map2T.scala 15:11]
  assign op_I0_15_1_2 = I0_15_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_8_2 = I1_8_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_9_2 = I1_9_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_10_2 = I1_10_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_11_2 = I1_11_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_12_2 = I1_12_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_13_2 = I1_13_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_14_2 = I1_14_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
  assign op_I1_15_2 = I1_15_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_8_1_0,
  input  [31:0] I_8_1_1,
  input  [31:0] I_8_1_2,
  input  [31:0] I_8_2_0,
  input  [31:0] I_8_2_1,
  input  [31:0] I_8_2_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_9_1_0,
  input  [31:0] I_9_1_1,
  input  [31:0] I_9_1_2,
  input  [31:0] I_9_2_0,
  input  [31:0] I_9_2_1,
  input  [31:0] I_9_2_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_10_1_0,
  input  [31:0] I_10_1_1,
  input  [31:0] I_10_1_2,
  input  [31:0] I_10_2_0,
  input  [31:0] I_10_2_1,
  input  [31:0] I_10_2_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_11_1_0,
  input  [31:0] I_11_1_1,
  input  [31:0] I_11_1_2,
  input  [31:0] I_11_2_0,
  input  [31:0] I_11_2_1,
  input  [31:0] I_11_2_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_12_1_0,
  input  [31:0] I_12_1_1,
  input  [31:0] I_12_1_2,
  input  [31:0] I_12_2_0,
  input  [31:0] I_12_2_1,
  input  [31:0] I_12_2_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_13_1_0,
  input  [31:0] I_13_1_1,
  input  [31:0] I_13_1_2,
  input  [31:0] I_13_2_0,
  input  [31:0] I_13_2_1,
  input  [31:0] I_13_2_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_14_1_0,
  input  [31:0] I_14_1_1,
  input  [31:0] I_14_1_2,
  input  [31:0] I_14_2_0,
  input  [31:0] I_14_2_1,
  input  [31:0] I_14_2_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  input  [31:0] I_15_1_0,
  input  [31:0] I_15_1_1,
  input  [31:0] I_15_1_2,
  input  [31:0] I_15_2_0,
  input  [31:0] I_15_2_1,
  input  [31:0] I_15_2_2,
  output [31:0] O_0_0_0_0,
  output [31:0] O_0_0_0_1,
  output [31:0] O_0_0_0_2,
  output [31:0] O_0_0_1_0,
  output [31:0] O_0_0_1_1,
  output [31:0] O_0_0_1_2,
  output [31:0] O_0_0_2_0,
  output [31:0] O_0_0_2_1,
  output [31:0] O_0_0_2_2,
  output [31:0] O_1_0_0_0,
  output [31:0] O_1_0_0_1,
  output [31:0] O_1_0_0_2,
  output [31:0] O_1_0_1_0,
  output [31:0] O_1_0_1_1,
  output [31:0] O_1_0_1_2,
  output [31:0] O_1_0_2_0,
  output [31:0] O_1_0_2_1,
  output [31:0] O_1_0_2_2,
  output [31:0] O_2_0_0_0,
  output [31:0] O_2_0_0_1,
  output [31:0] O_2_0_0_2,
  output [31:0] O_2_0_1_0,
  output [31:0] O_2_0_1_1,
  output [31:0] O_2_0_1_2,
  output [31:0] O_2_0_2_0,
  output [31:0] O_2_0_2_1,
  output [31:0] O_2_0_2_2,
  output [31:0] O_3_0_0_0,
  output [31:0] O_3_0_0_1,
  output [31:0] O_3_0_0_2,
  output [31:0] O_3_0_1_0,
  output [31:0] O_3_0_1_1,
  output [31:0] O_3_0_1_2,
  output [31:0] O_3_0_2_0,
  output [31:0] O_3_0_2_1,
  output [31:0] O_3_0_2_2,
  output [31:0] O_4_0_0_0,
  output [31:0] O_4_0_0_1,
  output [31:0] O_4_0_0_2,
  output [31:0] O_4_0_1_0,
  output [31:0] O_4_0_1_1,
  output [31:0] O_4_0_1_2,
  output [31:0] O_4_0_2_0,
  output [31:0] O_4_0_2_1,
  output [31:0] O_4_0_2_2,
  output [31:0] O_5_0_0_0,
  output [31:0] O_5_0_0_1,
  output [31:0] O_5_0_0_2,
  output [31:0] O_5_0_1_0,
  output [31:0] O_5_0_1_1,
  output [31:0] O_5_0_1_2,
  output [31:0] O_5_0_2_0,
  output [31:0] O_5_0_2_1,
  output [31:0] O_5_0_2_2,
  output [31:0] O_6_0_0_0,
  output [31:0] O_6_0_0_1,
  output [31:0] O_6_0_0_2,
  output [31:0] O_6_0_1_0,
  output [31:0] O_6_0_1_1,
  output [31:0] O_6_0_1_2,
  output [31:0] O_6_0_2_0,
  output [31:0] O_6_0_2_1,
  output [31:0] O_6_0_2_2,
  output [31:0] O_7_0_0_0,
  output [31:0] O_7_0_0_1,
  output [31:0] O_7_0_0_2,
  output [31:0] O_7_0_1_0,
  output [31:0] O_7_0_1_1,
  output [31:0] O_7_0_1_2,
  output [31:0] O_7_0_2_0,
  output [31:0] O_7_0_2_1,
  output [31:0] O_7_0_2_2,
  output [31:0] O_8_0_0_0,
  output [31:0] O_8_0_0_1,
  output [31:0] O_8_0_0_2,
  output [31:0] O_8_0_1_0,
  output [31:0] O_8_0_1_1,
  output [31:0] O_8_0_1_2,
  output [31:0] O_8_0_2_0,
  output [31:0] O_8_0_2_1,
  output [31:0] O_8_0_2_2,
  output [31:0] O_9_0_0_0,
  output [31:0] O_9_0_0_1,
  output [31:0] O_9_0_0_2,
  output [31:0] O_9_0_1_0,
  output [31:0] O_9_0_1_1,
  output [31:0] O_9_0_1_2,
  output [31:0] O_9_0_2_0,
  output [31:0] O_9_0_2_1,
  output [31:0] O_9_0_2_2,
  output [31:0] O_10_0_0_0,
  output [31:0] O_10_0_0_1,
  output [31:0] O_10_0_0_2,
  output [31:0] O_10_0_1_0,
  output [31:0] O_10_0_1_1,
  output [31:0] O_10_0_1_2,
  output [31:0] O_10_0_2_0,
  output [31:0] O_10_0_2_1,
  output [31:0] O_10_0_2_2,
  output [31:0] O_11_0_0_0,
  output [31:0] O_11_0_0_1,
  output [31:0] O_11_0_0_2,
  output [31:0] O_11_0_1_0,
  output [31:0] O_11_0_1_1,
  output [31:0] O_11_0_1_2,
  output [31:0] O_11_0_2_0,
  output [31:0] O_11_0_2_1,
  output [31:0] O_11_0_2_2,
  output [31:0] O_12_0_0_0,
  output [31:0] O_12_0_0_1,
  output [31:0] O_12_0_0_2,
  output [31:0] O_12_0_1_0,
  output [31:0] O_12_0_1_1,
  output [31:0] O_12_0_1_2,
  output [31:0] O_12_0_2_0,
  output [31:0] O_12_0_2_1,
  output [31:0] O_12_0_2_2,
  output [31:0] O_13_0_0_0,
  output [31:0] O_13_0_0_1,
  output [31:0] O_13_0_0_2,
  output [31:0] O_13_0_1_0,
  output [31:0] O_13_0_1_1,
  output [31:0] O_13_0_1_2,
  output [31:0] O_13_0_2_0,
  output [31:0] O_13_0_2_1,
  output [31:0] O_13_0_2_2,
  output [31:0] O_14_0_0_0,
  output [31:0] O_14_0_0_1,
  output [31:0] O_14_0_0_2,
  output [31:0] O_14_0_1_0,
  output [31:0] O_14_0_1_1,
  output [31:0] O_14_0_1_2,
  output [31:0] O_14_0_2_0,
  output [31:0] O_14_0_2_1,
  output [31:0] O_14_0_2_2,
  output [31:0] O_15_0_0_0,
  output [31:0] O_15_0_0_1,
  output [31:0] O_15_0_0_2,
  output [31:0] O_15_0_1_0,
  output [31:0] O_15_0_1_1,
  output [31:0] O_15_0_1_2,
  output [31:0] O_15_0_2_0,
  output [31:0] O_15_0_2_1,
  output [31:0] O_15_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_0_2 = I_4_0_2; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_4_0_1_2 = I_4_1_2; // @[Partition.scala 15:39]
  assign O_4_0_2_0 = I_4_2_0; // @[Partition.scala 15:39]
  assign O_4_0_2_1 = I_4_2_1; // @[Partition.scala 15:39]
  assign O_4_0_2_2 = I_4_2_2; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_0_2 = I_5_0_2; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_5_0_1_2 = I_5_1_2; // @[Partition.scala 15:39]
  assign O_5_0_2_0 = I_5_2_0; // @[Partition.scala 15:39]
  assign O_5_0_2_1 = I_5_2_1; // @[Partition.scala 15:39]
  assign O_5_0_2_2 = I_5_2_2; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_0_2 = I_6_0_2; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_6_0_1_2 = I_6_1_2; // @[Partition.scala 15:39]
  assign O_6_0_2_0 = I_6_2_0; // @[Partition.scala 15:39]
  assign O_6_0_2_1 = I_6_2_1; // @[Partition.scala 15:39]
  assign O_6_0_2_2 = I_6_2_2; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_0_2 = I_7_0_2; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_7_0_1_2 = I_7_1_2; // @[Partition.scala 15:39]
  assign O_7_0_2_0 = I_7_2_0; // @[Partition.scala 15:39]
  assign O_7_0_2_1 = I_7_2_1; // @[Partition.scala 15:39]
  assign O_7_0_2_2 = I_7_2_2; // @[Partition.scala 15:39]
  assign O_8_0_0_0 = I_8_0_0; // @[Partition.scala 15:39]
  assign O_8_0_0_1 = I_8_0_1; // @[Partition.scala 15:39]
  assign O_8_0_0_2 = I_8_0_2; // @[Partition.scala 15:39]
  assign O_8_0_1_0 = I_8_1_0; // @[Partition.scala 15:39]
  assign O_8_0_1_1 = I_8_1_1; // @[Partition.scala 15:39]
  assign O_8_0_1_2 = I_8_1_2; // @[Partition.scala 15:39]
  assign O_8_0_2_0 = I_8_2_0; // @[Partition.scala 15:39]
  assign O_8_0_2_1 = I_8_2_1; // @[Partition.scala 15:39]
  assign O_8_0_2_2 = I_8_2_2; // @[Partition.scala 15:39]
  assign O_9_0_0_0 = I_9_0_0; // @[Partition.scala 15:39]
  assign O_9_0_0_1 = I_9_0_1; // @[Partition.scala 15:39]
  assign O_9_0_0_2 = I_9_0_2; // @[Partition.scala 15:39]
  assign O_9_0_1_0 = I_9_1_0; // @[Partition.scala 15:39]
  assign O_9_0_1_1 = I_9_1_1; // @[Partition.scala 15:39]
  assign O_9_0_1_2 = I_9_1_2; // @[Partition.scala 15:39]
  assign O_9_0_2_0 = I_9_2_0; // @[Partition.scala 15:39]
  assign O_9_0_2_1 = I_9_2_1; // @[Partition.scala 15:39]
  assign O_9_0_2_2 = I_9_2_2; // @[Partition.scala 15:39]
  assign O_10_0_0_0 = I_10_0_0; // @[Partition.scala 15:39]
  assign O_10_0_0_1 = I_10_0_1; // @[Partition.scala 15:39]
  assign O_10_0_0_2 = I_10_0_2; // @[Partition.scala 15:39]
  assign O_10_0_1_0 = I_10_1_0; // @[Partition.scala 15:39]
  assign O_10_0_1_1 = I_10_1_1; // @[Partition.scala 15:39]
  assign O_10_0_1_2 = I_10_1_2; // @[Partition.scala 15:39]
  assign O_10_0_2_0 = I_10_2_0; // @[Partition.scala 15:39]
  assign O_10_0_2_1 = I_10_2_1; // @[Partition.scala 15:39]
  assign O_10_0_2_2 = I_10_2_2; // @[Partition.scala 15:39]
  assign O_11_0_0_0 = I_11_0_0; // @[Partition.scala 15:39]
  assign O_11_0_0_1 = I_11_0_1; // @[Partition.scala 15:39]
  assign O_11_0_0_2 = I_11_0_2; // @[Partition.scala 15:39]
  assign O_11_0_1_0 = I_11_1_0; // @[Partition.scala 15:39]
  assign O_11_0_1_1 = I_11_1_1; // @[Partition.scala 15:39]
  assign O_11_0_1_2 = I_11_1_2; // @[Partition.scala 15:39]
  assign O_11_0_2_0 = I_11_2_0; // @[Partition.scala 15:39]
  assign O_11_0_2_1 = I_11_2_1; // @[Partition.scala 15:39]
  assign O_11_0_2_2 = I_11_2_2; // @[Partition.scala 15:39]
  assign O_12_0_0_0 = I_12_0_0; // @[Partition.scala 15:39]
  assign O_12_0_0_1 = I_12_0_1; // @[Partition.scala 15:39]
  assign O_12_0_0_2 = I_12_0_2; // @[Partition.scala 15:39]
  assign O_12_0_1_0 = I_12_1_0; // @[Partition.scala 15:39]
  assign O_12_0_1_1 = I_12_1_1; // @[Partition.scala 15:39]
  assign O_12_0_1_2 = I_12_1_2; // @[Partition.scala 15:39]
  assign O_12_0_2_0 = I_12_2_0; // @[Partition.scala 15:39]
  assign O_12_0_2_1 = I_12_2_1; // @[Partition.scala 15:39]
  assign O_12_0_2_2 = I_12_2_2; // @[Partition.scala 15:39]
  assign O_13_0_0_0 = I_13_0_0; // @[Partition.scala 15:39]
  assign O_13_0_0_1 = I_13_0_1; // @[Partition.scala 15:39]
  assign O_13_0_0_2 = I_13_0_2; // @[Partition.scala 15:39]
  assign O_13_0_1_0 = I_13_1_0; // @[Partition.scala 15:39]
  assign O_13_0_1_1 = I_13_1_1; // @[Partition.scala 15:39]
  assign O_13_0_1_2 = I_13_1_2; // @[Partition.scala 15:39]
  assign O_13_0_2_0 = I_13_2_0; // @[Partition.scala 15:39]
  assign O_13_0_2_1 = I_13_2_1; // @[Partition.scala 15:39]
  assign O_13_0_2_2 = I_13_2_2; // @[Partition.scala 15:39]
  assign O_14_0_0_0 = I_14_0_0; // @[Partition.scala 15:39]
  assign O_14_0_0_1 = I_14_0_1; // @[Partition.scala 15:39]
  assign O_14_0_0_2 = I_14_0_2; // @[Partition.scala 15:39]
  assign O_14_0_1_0 = I_14_1_0; // @[Partition.scala 15:39]
  assign O_14_0_1_1 = I_14_1_1; // @[Partition.scala 15:39]
  assign O_14_0_1_2 = I_14_1_2; // @[Partition.scala 15:39]
  assign O_14_0_2_0 = I_14_2_0; // @[Partition.scala 15:39]
  assign O_14_0_2_1 = I_14_2_1; // @[Partition.scala 15:39]
  assign O_14_0_2_2 = I_14_2_2; // @[Partition.scala 15:39]
  assign O_15_0_0_0 = I_15_0_0; // @[Partition.scala 15:39]
  assign O_15_0_0_1 = I_15_0_1; // @[Partition.scala 15:39]
  assign O_15_0_0_2 = I_15_0_2; // @[Partition.scala 15:39]
  assign O_15_0_1_0 = I_15_1_0; // @[Partition.scala 15:39]
  assign O_15_0_1_1 = I_15_1_1; // @[Partition.scala 15:39]
  assign O_15_0_1_2 = I_15_1_2; // @[Partition.scala 15:39]
  assign O_15_0_2_0 = I_15_2_0; // @[Partition.scala 15:39]
  assign O_15_0_2_1 = I_15_2_1; // @[Partition.scala 15:39]
  assign O_15_0_2_2 = I_15_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_8_1_0,
  input  [31:0] I_8_1_1,
  input  [31:0] I_8_1_2,
  input  [31:0] I_8_2_0,
  input  [31:0] I_8_2_1,
  input  [31:0] I_8_2_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_9_1_0,
  input  [31:0] I_9_1_1,
  input  [31:0] I_9_1_2,
  input  [31:0] I_9_2_0,
  input  [31:0] I_9_2_1,
  input  [31:0] I_9_2_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_10_1_0,
  input  [31:0] I_10_1_1,
  input  [31:0] I_10_1_2,
  input  [31:0] I_10_2_0,
  input  [31:0] I_10_2_1,
  input  [31:0] I_10_2_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_11_1_0,
  input  [31:0] I_11_1_1,
  input  [31:0] I_11_1_2,
  input  [31:0] I_11_2_0,
  input  [31:0] I_11_2_1,
  input  [31:0] I_11_2_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_12_1_0,
  input  [31:0] I_12_1_1,
  input  [31:0] I_12_1_2,
  input  [31:0] I_12_2_0,
  input  [31:0] I_12_2_1,
  input  [31:0] I_12_2_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_13_1_0,
  input  [31:0] I_13_1_1,
  input  [31:0] I_13_1_2,
  input  [31:0] I_13_2_0,
  input  [31:0] I_13_2_1,
  input  [31:0] I_13_2_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_14_1_0,
  input  [31:0] I_14_1_1,
  input  [31:0] I_14_1_2,
  input  [31:0] I_14_2_0,
  input  [31:0] I_14_2_1,
  input  [31:0] I_14_2_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  input  [31:0] I_15_1_0,
  input  [31:0] I_15_1_1,
  input  [31:0] I_15_1_2,
  input  [31:0] I_15_2_0,
  input  [31:0] I_15_2_1,
  input  [31:0] I_15_2_2,
  output [31:0] O_0_0_0_0,
  output [31:0] O_0_0_0_1,
  output [31:0] O_0_0_0_2,
  output [31:0] O_0_0_1_0,
  output [31:0] O_0_0_1_1,
  output [31:0] O_0_0_1_2,
  output [31:0] O_0_0_2_0,
  output [31:0] O_0_0_2_1,
  output [31:0] O_0_0_2_2,
  output [31:0] O_1_0_0_0,
  output [31:0] O_1_0_0_1,
  output [31:0] O_1_0_0_2,
  output [31:0] O_1_0_1_0,
  output [31:0] O_1_0_1_1,
  output [31:0] O_1_0_1_2,
  output [31:0] O_1_0_2_0,
  output [31:0] O_1_0_2_1,
  output [31:0] O_1_0_2_2,
  output [31:0] O_2_0_0_0,
  output [31:0] O_2_0_0_1,
  output [31:0] O_2_0_0_2,
  output [31:0] O_2_0_1_0,
  output [31:0] O_2_0_1_1,
  output [31:0] O_2_0_1_2,
  output [31:0] O_2_0_2_0,
  output [31:0] O_2_0_2_1,
  output [31:0] O_2_0_2_2,
  output [31:0] O_3_0_0_0,
  output [31:0] O_3_0_0_1,
  output [31:0] O_3_0_0_2,
  output [31:0] O_3_0_1_0,
  output [31:0] O_3_0_1_1,
  output [31:0] O_3_0_1_2,
  output [31:0] O_3_0_2_0,
  output [31:0] O_3_0_2_1,
  output [31:0] O_3_0_2_2,
  output [31:0] O_4_0_0_0,
  output [31:0] O_4_0_0_1,
  output [31:0] O_4_0_0_2,
  output [31:0] O_4_0_1_0,
  output [31:0] O_4_0_1_1,
  output [31:0] O_4_0_1_2,
  output [31:0] O_4_0_2_0,
  output [31:0] O_4_0_2_1,
  output [31:0] O_4_0_2_2,
  output [31:0] O_5_0_0_0,
  output [31:0] O_5_0_0_1,
  output [31:0] O_5_0_0_2,
  output [31:0] O_5_0_1_0,
  output [31:0] O_5_0_1_1,
  output [31:0] O_5_0_1_2,
  output [31:0] O_5_0_2_0,
  output [31:0] O_5_0_2_1,
  output [31:0] O_5_0_2_2,
  output [31:0] O_6_0_0_0,
  output [31:0] O_6_0_0_1,
  output [31:0] O_6_0_0_2,
  output [31:0] O_6_0_1_0,
  output [31:0] O_6_0_1_1,
  output [31:0] O_6_0_1_2,
  output [31:0] O_6_0_2_0,
  output [31:0] O_6_0_2_1,
  output [31:0] O_6_0_2_2,
  output [31:0] O_7_0_0_0,
  output [31:0] O_7_0_0_1,
  output [31:0] O_7_0_0_2,
  output [31:0] O_7_0_1_0,
  output [31:0] O_7_0_1_1,
  output [31:0] O_7_0_1_2,
  output [31:0] O_7_0_2_0,
  output [31:0] O_7_0_2_1,
  output [31:0] O_7_0_2_2,
  output [31:0] O_8_0_0_0,
  output [31:0] O_8_0_0_1,
  output [31:0] O_8_0_0_2,
  output [31:0] O_8_0_1_0,
  output [31:0] O_8_0_1_1,
  output [31:0] O_8_0_1_2,
  output [31:0] O_8_0_2_0,
  output [31:0] O_8_0_2_1,
  output [31:0] O_8_0_2_2,
  output [31:0] O_9_0_0_0,
  output [31:0] O_9_0_0_1,
  output [31:0] O_9_0_0_2,
  output [31:0] O_9_0_1_0,
  output [31:0] O_9_0_1_1,
  output [31:0] O_9_0_1_2,
  output [31:0] O_9_0_2_0,
  output [31:0] O_9_0_2_1,
  output [31:0] O_9_0_2_2,
  output [31:0] O_10_0_0_0,
  output [31:0] O_10_0_0_1,
  output [31:0] O_10_0_0_2,
  output [31:0] O_10_0_1_0,
  output [31:0] O_10_0_1_1,
  output [31:0] O_10_0_1_2,
  output [31:0] O_10_0_2_0,
  output [31:0] O_10_0_2_1,
  output [31:0] O_10_0_2_2,
  output [31:0] O_11_0_0_0,
  output [31:0] O_11_0_0_1,
  output [31:0] O_11_0_0_2,
  output [31:0] O_11_0_1_0,
  output [31:0] O_11_0_1_1,
  output [31:0] O_11_0_1_2,
  output [31:0] O_11_0_2_0,
  output [31:0] O_11_0_2_1,
  output [31:0] O_11_0_2_2,
  output [31:0] O_12_0_0_0,
  output [31:0] O_12_0_0_1,
  output [31:0] O_12_0_0_2,
  output [31:0] O_12_0_1_0,
  output [31:0] O_12_0_1_1,
  output [31:0] O_12_0_1_2,
  output [31:0] O_12_0_2_0,
  output [31:0] O_12_0_2_1,
  output [31:0] O_12_0_2_2,
  output [31:0] O_13_0_0_0,
  output [31:0] O_13_0_0_1,
  output [31:0] O_13_0_0_2,
  output [31:0] O_13_0_1_0,
  output [31:0] O_13_0_1_1,
  output [31:0] O_13_0_1_2,
  output [31:0] O_13_0_2_0,
  output [31:0] O_13_0_2_1,
  output [31:0] O_13_0_2_2,
  output [31:0] O_14_0_0_0,
  output [31:0] O_14_0_0_1,
  output [31:0] O_14_0_0_2,
  output [31:0] O_14_0_1_0,
  output [31:0] O_14_0_1_1,
  output [31:0] O_14_0_1_2,
  output [31:0] O_14_0_2_0,
  output [31:0] O_14_0_2_1,
  output [31:0] O_14_0_2_2,
  output [31:0] O_15_0_0_0,
  output [31:0] O_15_0_0_1,
  output [31:0] O_15_0_0_2,
  output [31:0] O_15_0_1_0,
  output [31:0] O_15_0_1_1,
  output [31:0] O_15_0_1_2,
  output [31:0] O_15_0_2_0,
  output [31:0] O_15_0_2_1,
  output [31:0] O_15_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_0_2(op_O_8_0_0_2),
    .O_8_0_1_0(op_O_8_0_1_0),
    .O_8_0_1_1(op_O_8_0_1_1),
    .O_8_0_1_2(op_O_8_0_1_2),
    .O_8_0_2_0(op_O_8_0_2_0),
    .O_8_0_2_1(op_O_8_0_2_1),
    .O_8_0_2_2(op_O_8_0_2_2),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_0_2(op_O_9_0_0_2),
    .O_9_0_1_0(op_O_9_0_1_0),
    .O_9_0_1_1(op_O_9_0_1_1),
    .O_9_0_1_2(op_O_9_0_1_2),
    .O_9_0_2_0(op_O_9_0_2_0),
    .O_9_0_2_1(op_O_9_0_2_1),
    .O_9_0_2_2(op_O_9_0_2_2),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_0_2(op_O_10_0_0_2),
    .O_10_0_1_0(op_O_10_0_1_0),
    .O_10_0_1_1(op_O_10_0_1_1),
    .O_10_0_1_2(op_O_10_0_1_2),
    .O_10_0_2_0(op_O_10_0_2_0),
    .O_10_0_2_1(op_O_10_0_2_1),
    .O_10_0_2_2(op_O_10_0_2_2),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_0_2(op_O_11_0_0_2),
    .O_11_0_1_0(op_O_11_0_1_0),
    .O_11_0_1_1(op_O_11_0_1_1),
    .O_11_0_1_2(op_O_11_0_1_2),
    .O_11_0_2_0(op_O_11_0_2_0),
    .O_11_0_2_1(op_O_11_0_2_1),
    .O_11_0_2_2(op_O_11_0_2_2),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_0_2(op_O_12_0_0_2),
    .O_12_0_1_0(op_O_12_0_1_0),
    .O_12_0_1_1(op_O_12_0_1_1),
    .O_12_0_1_2(op_O_12_0_1_2),
    .O_12_0_2_0(op_O_12_0_2_0),
    .O_12_0_2_1(op_O_12_0_2_1),
    .O_12_0_2_2(op_O_12_0_2_2),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_0_2(op_O_13_0_0_2),
    .O_13_0_1_0(op_O_13_0_1_0),
    .O_13_0_1_1(op_O_13_0_1_1),
    .O_13_0_1_2(op_O_13_0_1_2),
    .O_13_0_2_0(op_O_13_0_2_0),
    .O_13_0_2_1(op_O_13_0_2_1),
    .O_13_0_2_2(op_O_13_0_2_2),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_0_2(op_O_14_0_0_2),
    .O_14_0_1_0(op_O_14_0_1_0),
    .O_14_0_1_1(op_O_14_0_1_1),
    .O_14_0_1_2(op_O_14_0_1_2),
    .O_14_0_2_0(op_O_14_0_2_0),
    .O_14_0_2_1(op_O_14_0_2_1),
    .O_14_0_2_2(op_O_14_0_2_2),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_0_2(op_O_15_0_0_2),
    .O_15_0_1_0(op_O_15_0_1_0),
    .O_15_0_1_1(op_O_15_0_1_1),
    .O_15_0_1_2(op_O_15_0_1_2),
    .O_15_0_2_0(op_O_15_0_2_0),
    .O_15_0_2_1(op_O_15_0_2_1),
    .O_15_0_2_2(op_O_15_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[MapT.scala 15:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[MapT.scala 15:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[MapT.scala 15:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[MapT.scala 15:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[MapT.scala 15:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[MapT.scala 15:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[MapT.scala 15:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[MapT.scala 15:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[MapT.scala 15:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[MapT.scala 15:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[MapT.scala 15:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[MapT.scala 15:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[MapT.scala 15:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[MapT.scala 15:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[MapT.scala 15:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[MapT.scala 15:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[MapT.scala 15:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[MapT.scala 15:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[MapT.scala 15:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[MapT.scala 15:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[MapT.scala 15:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[MapT.scala 15:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[MapT.scala 15:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[MapT.scala 15:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[MapT.scala 15:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[MapT.scala 15:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[MapT.scala 15:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[MapT.scala 15:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[MapT.scala 15:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[MapT.scala 15:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[MapT.scala 15:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[MapT.scala 15:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[MapT.scala 15:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[MapT.scala 15:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[MapT.scala 15:7]
  assign O_8_0_0_2 = op_O_8_0_0_2; // @[MapT.scala 15:7]
  assign O_8_0_1_0 = op_O_8_0_1_0; // @[MapT.scala 15:7]
  assign O_8_0_1_1 = op_O_8_0_1_1; // @[MapT.scala 15:7]
  assign O_8_0_1_2 = op_O_8_0_1_2; // @[MapT.scala 15:7]
  assign O_8_0_2_0 = op_O_8_0_2_0; // @[MapT.scala 15:7]
  assign O_8_0_2_1 = op_O_8_0_2_1; // @[MapT.scala 15:7]
  assign O_8_0_2_2 = op_O_8_0_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[MapT.scala 15:7]
  assign O_9_0_0_2 = op_O_9_0_0_2; // @[MapT.scala 15:7]
  assign O_9_0_1_0 = op_O_9_0_1_0; // @[MapT.scala 15:7]
  assign O_9_0_1_1 = op_O_9_0_1_1; // @[MapT.scala 15:7]
  assign O_9_0_1_2 = op_O_9_0_1_2; // @[MapT.scala 15:7]
  assign O_9_0_2_0 = op_O_9_0_2_0; // @[MapT.scala 15:7]
  assign O_9_0_2_1 = op_O_9_0_2_1; // @[MapT.scala 15:7]
  assign O_9_0_2_2 = op_O_9_0_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[MapT.scala 15:7]
  assign O_10_0_0_2 = op_O_10_0_0_2; // @[MapT.scala 15:7]
  assign O_10_0_1_0 = op_O_10_0_1_0; // @[MapT.scala 15:7]
  assign O_10_0_1_1 = op_O_10_0_1_1; // @[MapT.scala 15:7]
  assign O_10_0_1_2 = op_O_10_0_1_2; // @[MapT.scala 15:7]
  assign O_10_0_2_0 = op_O_10_0_2_0; // @[MapT.scala 15:7]
  assign O_10_0_2_1 = op_O_10_0_2_1; // @[MapT.scala 15:7]
  assign O_10_0_2_2 = op_O_10_0_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[MapT.scala 15:7]
  assign O_11_0_0_2 = op_O_11_0_0_2; // @[MapT.scala 15:7]
  assign O_11_0_1_0 = op_O_11_0_1_0; // @[MapT.scala 15:7]
  assign O_11_0_1_1 = op_O_11_0_1_1; // @[MapT.scala 15:7]
  assign O_11_0_1_2 = op_O_11_0_1_2; // @[MapT.scala 15:7]
  assign O_11_0_2_0 = op_O_11_0_2_0; // @[MapT.scala 15:7]
  assign O_11_0_2_1 = op_O_11_0_2_1; // @[MapT.scala 15:7]
  assign O_11_0_2_2 = op_O_11_0_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[MapT.scala 15:7]
  assign O_12_0_0_2 = op_O_12_0_0_2; // @[MapT.scala 15:7]
  assign O_12_0_1_0 = op_O_12_0_1_0; // @[MapT.scala 15:7]
  assign O_12_0_1_1 = op_O_12_0_1_1; // @[MapT.scala 15:7]
  assign O_12_0_1_2 = op_O_12_0_1_2; // @[MapT.scala 15:7]
  assign O_12_0_2_0 = op_O_12_0_2_0; // @[MapT.scala 15:7]
  assign O_12_0_2_1 = op_O_12_0_2_1; // @[MapT.scala 15:7]
  assign O_12_0_2_2 = op_O_12_0_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[MapT.scala 15:7]
  assign O_13_0_0_2 = op_O_13_0_0_2; // @[MapT.scala 15:7]
  assign O_13_0_1_0 = op_O_13_0_1_0; // @[MapT.scala 15:7]
  assign O_13_0_1_1 = op_O_13_0_1_1; // @[MapT.scala 15:7]
  assign O_13_0_1_2 = op_O_13_0_1_2; // @[MapT.scala 15:7]
  assign O_13_0_2_0 = op_O_13_0_2_0; // @[MapT.scala 15:7]
  assign O_13_0_2_1 = op_O_13_0_2_1; // @[MapT.scala 15:7]
  assign O_13_0_2_2 = op_O_13_0_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[MapT.scala 15:7]
  assign O_14_0_0_2 = op_O_14_0_0_2; // @[MapT.scala 15:7]
  assign O_14_0_1_0 = op_O_14_0_1_0; // @[MapT.scala 15:7]
  assign O_14_0_1_1 = op_O_14_0_1_1; // @[MapT.scala 15:7]
  assign O_14_0_1_2 = op_O_14_0_1_2; // @[MapT.scala 15:7]
  assign O_14_0_2_0 = op_O_14_0_2_0; // @[MapT.scala 15:7]
  assign O_14_0_2_1 = op_O_14_0_2_1; // @[MapT.scala 15:7]
  assign O_14_0_2_2 = op_O_14_0_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[MapT.scala 15:7]
  assign O_15_0_0_2 = op_O_15_0_0_2; // @[MapT.scala 15:7]
  assign O_15_0_1_0 = op_O_15_0_1_0; // @[MapT.scala 15:7]
  assign O_15_0_1_1 = op_O_15_0_1_1; // @[MapT.scala 15:7]
  assign O_15_0_1_2 = op_O_15_0_1_2; // @[MapT.scala 15:7]
  assign O_15_0_2_0 = op_O_15_0_2_0; // @[MapT.scala 15:7]
  assign O_15_0_2_1 = op_O_15_0_2_1; // @[MapT.scala 15:7]
  assign O_15_0_2_2 = op_O_15_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_1_0,
  output [31:0] O_1_1,
  output [31:0] O_1_2,
  output [31:0] O_2_0,
  output [31:0] O_2_1,
  output [31:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_0,
  input  [31:0] I_0_0_0_1,
  input  [31:0] I_0_0_0_2,
  input  [31:0] I_0_0_1_0,
  input  [31:0] I_0_0_1_1,
  input  [31:0] I_0_0_1_2,
  input  [31:0] I_0_0_2_0,
  input  [31:0] I_0_0_2_1,
  input  [31:0] I_0_0_2_2,
  input  [31:0] I_1_0_0_0,
  input  [31:0] I_1_0_0_1,
  input  [31:0] I_1_0_0_2,
  input  [31:0] I_1_0_1_0,
  input  [31:0] I_1_0_1_1,
  input  [31:0] I_1_0_1_2,
  input  [31:0] I_1_0_2_0,
  input  [31:0] I_1_0_2_1,
  input  [31:0] I_1_0_2_2,
  input  [31:0] I_2_0_0_0,
  input  [31:0] I_2_0_0_1,
  input  [31:0] I_2_0_0_2,
  input  [31:0] I_2_0_1_0,
  input  [31:0] I_2_0_1_1,
  input  [31:0] I_2_0_1_2,
  input  [31:0] I_2_0_2_0,
  input  [31:0] I_2_0_2_1,
  input  [31:0] I_2_0_2_2,
  input  [31:0] I_3_0_0_0,
  input  [31:0] I_3_0_0_1,
  input  [31:0] I_3_0_0_2,
  input  [31:0] I_3_0_1_0,
  input  [31:0] I_3_0_1_1,
  input  [31:0] I_3_0_1_2,
  input  [31:0] I_3_0_2_0,
  input  [31:0] I_3_0_2_1,
  input  [31:0] I_3_0_2_2,
  input  [31:0] I_4_0_0_0,
  input  [31:0] I_4_0_0_1,
  input  [31:0] I_4_0_0_2,
  input  [31:0] I_4_0_1_0,
  input  [31:0] I_4_0_1_1,
  input  [31:0] I_4_0_1_2,
  input  [31:0] I_4_0_2_0,
  input  [31:0] I_4_0_2_1,
  input  [31:0] I_4_0_2_2,
  input  [31:0] I_5_0_0_0,
  input  [31:0] I_5_0_0_1,
  input  [31:0] I_5_0_0_2,
  input  [31:0] I_5_0_1_0,
  input  [31:0] I_5_0_1_1,
  input  [31:0] I_5_0_1_2,
  input  [31:0] I_5_0_2_0,
  input  [31:0] I_5_0_2_1,
  input  [31:0] I_5_0_2_2,
  input  [31:0] I_6_0_0_0,
  input  [31:0] I_6_0_0_1,
  input  [31:0] I_6_0_0_2,
  input  [31:0] I_6_0_1_0,
  input  [31:0] I_6_0_1_1,
  input  [31:0] I_6_0_1_2,
  input  [31:0] I_6_0_2_0,
  input  [31:0] I_6_0_2_1,
  input  [31:0] I_6_0_2_2,
  input  [31:0] I_7_0_0_0,
  input  [31:0] I_7_0_0_1,
  input  [31:0] I_7_0_0_2,
  input  [31:0] I_7_0_1_0,
  input  [31:0] I_7_0_1_1,
  input  [31:0] I_7_0_1_2,
  input  [31:0] I_7_0_2_0,
  input  [31:0] I_7_0_2_1,
  input  [31:0] I_7_0_2_2,
  input  [31:0] I_8_0_0_0,
  input  [31:0] I_8_0_0_1,
  input  [31:0] I_8_0_0_2,
  input  [31:0] I_8_0_1_0,
  input  [31:0] I_8_0_1_1,
  input  [31:0] I_8_0_1_2,
  input  [31:0] I_8_0_2_0,
  input  [31:0] I_8_0_2_1,
  input  [31:0] I_8_0_2_2,
  input  [31:0] I_9_0_0_0,
  input  [31:0] I_9_0_0_1,
  input  [31:0] I_9_0_0_2,
  input  [31:0] I_9_0_1_0,
  input  [31:0] I_9_0_1_1,
  input  [31:0] I_9_0_1_2,
  input  [31:0] I_9_0_2_0,
  input  [31:0] I_9_0_2_1,
  input  [31:0] I_9_0_2_2,
  input  [31:0] I_10_0_0_0,
  input  [31:0] I_10_0_0_1,
  input  [31:0] I_10_0_0_2,
  input  [31:0] I_10_0_1_0,
  input  [31:0] I_10_0_1_1,
  input  [31:0] I_10_0_1_2,
  input  [31:0] I_10_0_2_0,
  input  [31:0] I_10_0_2_1,
  input  [31:0] I_10_0_2_2,
  input  [31:0] I_11_0_0_0,
  input  [31:0] I_11_0_0_1,
  input  [31:0] I_11_0_0_2,
  input  [31:0] I_11_0_1_0,
  input  [31:0] I_11_0_1_1,
  input  [31:0] I_11_0_1_2,
  input  [31:0] I_11_0_2_0,
  input  [31:0] I_11_0_2_1,
  input  [31:0] I_11_0_2_2,
  input  [31:0] I_12_0_0_0,
  input  [31:0] I_12_0_0_1,
  input  [31:0] I_12_0_0_2,
  input  [31:0] I_12_0_1_0,
  input  [31:0] I_12_0_1_1,
  input  [31:0] I_12_0_1_2,
  input  [31:0] I_12_0_2_0,
  input  [31:0] I_12_0_2_1,
  input  [31:0] I_12_0_2_2,
  input  [31:0] I_13_0_0_0,
  input  [31:0] I_13_0_0_1,
  input  [31:0] I_13_0_0_2,
  input  [31:0] I_13_0_1_0,
  input  [31:0] I_13_0_1_1,
  input  [31:0] I_13_0_1_2,
  input  [31:0] I_13_0_2_0,
  input  [31:0] I_13_0_2_1,
  input  [31:0] I_13_0_2_2,
  input  [31:0] I_14_0_0_0,
  input  [31:0] I_14_0_0_1,
  input  [31:0] I_14_0_0_2,
  input  [31:0] I_14_0_1_0,
  input  [31:0] I_14_0_1_1,
  input  [31:0] I_14_0_1_2,
  input  [31:0] I_14_0_2_0,
  input  [31:0] I_14_0_2_1,
  input  [31:0] I_14_0_2_2,
  input  [31:0] I_15_0_0_0,
  input  [31:0] I_15_0_0_1,
  input  [31:0] I_15_0_0_2,
  input  [31:0] I_15_0_1_0,
  input  [31:0] I_15_0_1_1,
  input  [31:0] I_15_0_1_2,
  input  [31:0] I_15_0_2_0,
  input  [31:0] I_15_0_2_1,
  input  [31:0] I_15_0_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_8_2_0,
  output [31:0] O_8_2_1,
  output [31:0] O_8_2_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_9_2_0,
  output [31:0] O_9_2_1,
  output [31:0] O_9_2_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_10_2_0,
  output [31:0] O_10_2_1,
  output [31:0] O_10_2_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_11_2_0,
  output [31:0] O_11_2_1,
  output [31:0] O_11_2_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_12_2_0,
  output [31:0] O_12_2_1,
  output [31:0] O_12_2_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_13_2_0,
  output [31:0] O_13_2_1,
  output [31:0] O_13_2_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_14_2_0,
  output [31:0] O_14_2_1,
  output [31:0] O_14_2_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2,
  output [31:0] O_15_2_0,
  output [31:0] O_15_2_1,
  output [31:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I_0_2_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_0_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_1_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_1_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_1_2; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_2_0; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_2_1; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  Remove1S_3 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_0_2(other_ops_7_I_0_0_2),
    .I_0_1_0(other_ops_7_I_0_1_0),
    .I_0_1_1(other_ops_7_I_0_1_1),
    .I_0_1_2(other_ops_7_I_0_1_2),
    .I_0_2_0(other_ops_7_I_0_2_0),
    .I_0_2_1(other_ops_7_I_0_2_1),
    .I_0_2_2(other_ops_7_I_0_2_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  Remove1S_3 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_0_2(other_ops_8_I_0_0_2),
    .I_0_1_0(other_ops_8_I_0_1_0),
    .I_0_1_1(other_ops_8_I_0_1_1),
    .I_0_1_2(other_ops_8_I_0_1_2),
    .I_0_2_0(other_ops_8_I_0_2_0),
    .I_0_2_1(other_ops_8_I_0_2_1),
    .I_0_2_2(other_ops_8_I_0_2_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  Remove1S_3 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_0_2(other_ops_9_I_0_0_2),
    .I_0_1_0(other_ops_9_I_0_1_0),
    .I_0_1_1(other_ops_9_I_0_1_1),
    .I_0_1_2(other_ops_9_I_0_1_2),
    .I_0_2_0(other_ops_9_I_0_2_0),
    .I_0_2_1(other_ops_9_I_0_2_1),
    .I_0_2_2(other_ops_9_I_0_2_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  Remove1S_3 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_0_2(other_ops_10_I_0_0_2),
    .I_0_1_0(other_ops_10_I_0_1_0),
    .I_0_1_1(other_ops_10_I_0_1_1),
    .I_0_1_2(other_ops_10_I_0_1_2),
    .I_0_2_0(other_ops_10_I_0_2_0),
    .I_0_2_1(other_ops_10_I_0_2_1),
    .I_0_2_2(other_ops_10_I_0_2_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  Remove1S_3 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_0_2(other_ops_11_I_0_0_2),
    .I_0_1_0(other_ops_11_I_0_1_0),
    .I_0_1_1(other_ops_11_I_0_1_1),
    .I_0_1_2(other_ops_11_I_0_1_2),
    .I_0_2_0(other_ops_11_I_0_2_0),
    .I_0_2_1(other_ops_11_I_0_2_1),
    .I_0_2_2(other_ops_11_I_0_2_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  Remove1S_3 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_0_2(other_ops_12_I_0_0_2),
    .I_0_1_0(other_ops_12_I_0_1_0),
    .I_0_1_1(other_ops_12_I_0_1_1),
    .I_0_1_2(other_ops_12_I_0_1_2),
    .I_0_2_0(other_ops_12_I_0_2_0),
    .I_0_2_1(other_ops_12_I_0_2_1),
    .I_0_2_2(other_ops_12_I_0_2_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  Remove1S_3 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_0_2(other_ops_13_I_0_0_2),
    .I_0_1_0(other_ops_13_I_0_1_0),
    .I_0_1_1(other_ops_13_I_0_1_1),
    .I_0_1_2(other_ops_13_I_0_1_2),
    .I_0_2_0(other_ops_13_I_0_2_0),
    .I_0_2_1(other_ops_13_I_0_2_1),
    .I_0_2_2(other_ops_13_I_0_2_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  Remove1S_3 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_0_2(other_ops_14_I_0_0_2),
    .I_0_1_0(other_ops_14_I_0_1_0),
    .I_0_1_1(other_ops_14_I_0_1_1),
    .I_0_1_2(other_ops_14_I_0_1_2),
    .I_0_2_0(other_ops_14_I_0_2_0),
    .I_0_2_1(other_ops_14_I_0_2_1),
    .I_0_2_2(other_ops_14_I_0_2_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[MapS.scala 21:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[MapS.scala 21:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[MapS.scala 21:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[MapS.scala 21:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[MapS.scala 21:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[MapS.scala 21:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[MapS.scala 21:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[MapS.scala 21:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[MapS.scala 21:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[MapS.scala 21:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[MapS.scala 21:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[MapS.scala 21:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[MapS.scala 21:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[MapS.scala 21:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[MapS.scala 21:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[MapS.scala 21:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[MapS.scala 21:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[MapS.scala 21:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[MapS.scala 21:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[MapS.scala 21:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[MapS.scala 21:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[MapS.scala 21:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[MapS.scala 21:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[MapS.scala 21:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[MapS.scala 21:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[MapS.scala 21:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[MapS.scala 21:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[MapS.scala 21:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[MapS.scala 21:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[MapS.scala 21:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[MapS.scala 21:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[MapS.scala 21:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[MapS.scala 21:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[MapS.scala 21:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[MapS.scala 21:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[MapS.scala 21:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[MapS.scala 21:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[MapS.scala 21:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[MapS.scala 21:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[MapS.scala 21:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[MapS.scala 21:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[MapS.scala 21:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[MapS.scala 21:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[MapS.scala 21:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[MapS.scala 21:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[MapS.scala 21:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[MapS.scala 21:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[MapS.scala 21:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_2 = I_8_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_0 = I_8_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_1 = I_8_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_2 = I_8_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_0 = I_8_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_1 = I_8_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_2 = I_8_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_2 = I_9_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_0 = I_9_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_1 = I_9_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_2 = I_9_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_0 = I_9_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_1 = I_9_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_2 = I_9_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_2 = I_10_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_0 = I_10_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_1 = I_10_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_2 = I_10_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_0 = I_10_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_1 = I_10_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_2 = I_10_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_2 = I_11_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_0 = I_11_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_1 = I_11_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_2 = I_11_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_0 = I_11_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_1 = I_11_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_2 = I_11_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_2 = I_12_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_0 = I_12_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_1 = I_12_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_2 = I_12_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_0 = I_12_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_1 = I_12_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_2 = I_12_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_2 = I_13_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_0 = I_13_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_1 = I_13_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_2 = I_13_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_0 = I_13_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_1 = I_13_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_2 = I_13_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_2 = I_14_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_0 = I_14_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_1 = I_14_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_2 = I_14_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_0 = I_14_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_1 = I_14_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_2 = I_14_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_2 = I_15_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_0 = I_15_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_1 = I_15_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_2 = I_15_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_0 = I_15_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_1 = I_15_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_2 = I_15_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_0,
  input  [31:0] I_0_0_0_1,
  input  [31:0] I_0_0_0_2,
  input  [31:0] I_0_0_1_0,
  input  [31:0] I_0_0_1_1,
  input  [31:0] I_0_0_1_2,
  input  [31:0] I_0_0_2_0,
  input  [31:0] I_0_0_2_1,
  input  [31:0] I_0_0_2_2,
  input  [31:0] I_1_0_0_0,
  input  [31:0] I_1_0_0_1,
  input  [31:0] I_1_0_0_2,
  input  [31:0] I_1_0_1_0,
  input  [31:0] I_1_0_1_1,
  input  [31:0] I_1_0_1_2,
  input  [31:0] I_1_0_2_0,
  input  [31:0] I_1_0_2_1,
  input  [31:0] I_1_0_2_2,
  input  [31:0] I_2_0_0_0,
  input  [31:0] I_2_0_0_1,
  input  [31:0] I_2_0_0_2,
  input  [31:0] I_2_0_1_0,
  input  [31:0] I_2_0_1_1,
  input  [31:0] I_2_0_1_2,
  input  [31:0] I_2_0_2_0,
  input  [31:0] I_2_0_2_1,
  input  [31:0] I_2_0_2_2,
  input  [31:0] I_3_0_0_0,
  input  [31:0] I_3_0_0_1,
  input  [31:0] I_3_0_0_2,
  input  [31:0] I_3_0_1_0,
  input  [31:0] I_3_0_1_1,
  input  [31:0] I_3_0_1_2,
  input  [31:0] I_3_0_2_0,
  input  [31:0] I_3_0_2_1,
  input  [31:0] I_3_0_2_2,
  input  [31:0] I_4_0_0_0,
  input  [31:0] I_4_0_0_1,
  input  [31:0] I_4_0_0_2,
  input  [31:0] I_4_0_1_0,
  input  [31:0] I_4_0_1_1,
  input  [31:0] I_4_0_1_2,
  input  [31:0] I_4_0_2_0,
  input  [31:0] I_4_0_2_1,
  input  [31:0] I_4_0_2_2,
  input  [31:0] I_5_0_0_0,
  input  [31:0] I_5_0_0_1,
  input  [31:0] I_5_0_0_2,
  input  [31:0] I_5_0_1_0,
  input  [31:0] I_5_0_1_1,
  input  [31:0] I_5_0_1_2,
  input  [31:0] I_5_0_2_0,
  input  [31:0] I_5_0_2_1,
  input  [31:0] I_5_0_2_2,
  input  [31:0] I_6_0_0_0,
  input  [31:0] I_6_0_0_1,
  input  [31:0] I_6_0_0_2,
  input  [31:0] I_6_0_1_0,
  input  [31:0] I_6_0_1_1,
  input  [31:0] I_6_0_1_2,
  input  [31:0] I_6_0_2_0,
  input  [31:0] I_6_0_2_1,
  input  [31:0] I_6_0_2_2,
  input  [31:0] I_7_0_0_0,
  input  [31:0] I_7_0_0_1,
  input  [31:0] I_7_0_0_2,
  input  [31:0] I_7_0_1_0,
  input  [31:0] I_7_0_1_1,
  input  [31:0] I_7_0_1_2,
  input  [31:0] I_7_0_2_0,
  input  [31:0] I_7_0_2_1,
  input  [31:0] I_7_0_2_2,
  input  [31:0] I_8_0_0_0,
  input  [31:0] I_8_0_0_1,
  input  [31:0] I_8_0_0_2,
  input  [31:0] I_8_0_1_0,
  input  [31:0] I_8_0_1_1,
  input  [31:0] I_8_0_1_2,
  input  [31:0] I_8_0_2_0,
  input  [31:0] I_8_0_2_1,
  input  [31:0] I_8_0_2_2,
  input  [31:0] I_9_0_0_0,
  input  [31:0] I_9_0_0_1,
  input  [31:0] I_9_0_0_2,
  input  [31:0] I_9_0_1_0,
  input  [31:0] I_9_0_1_1,
  input  [31:0] I_9_0_1_2,
  input  [31:0] I_9_0_2_0,
  input  [31:0] I_9_0_2_1,
  input  [31:0] I_9_0_2_2,
  input  [31:0] I_10_0_0_0,
  input  [31:0] I_10_0_0_1,
  input  [31:0] I_10_0_0_2,
  input  [31:0] I_10_0_1_0,
  input  [31:0] I_10_0_1_1,
  input  [31:0] I_10_0_1_2,
  input  [31:0] I_10_0_2_0,
  input  [31:0] I_10_0_2_1,
  input  [31:0] I_10_0_2_2,
  input  [31:0] I_11_0_0_0,
  input  [31:0] I_11_0_0_1,
  input  [31:0] I_11_0_0_2,
  input  [31:0] I_11_0_1_0,
  input  [31:0] I_11_0_1_1,
  input  [31:0] I_11_0_1_2,
  input  [31:0] I_11_0_2_0,
  input  [31:0] I_11_0_2_1,
  input  [31:0] I_11_0_2_2,
  input  [31:0] I_12_0_0_0,
  input  [31:0] I_12_0_0_1,
  input  [31:0] I_12_0_0_2,
  input  [31:0] I_12_0_1_0,
  input  [31:0] I_12_0_1_1,
  input  [31:0] I_12_0_1_2,
  input  [31:0] I_12_0_2_0,
  input  [31:0] I_12_0_2_1,
  input  [31:0] I_12_0_2_2,
  input  [31:0] I_13_0_0_0,
  input  [31:0] I_13_0_0_1,
  input  [31:0] I_13_0_0_2,
  input  [31:0] I_13_0_1_0,
  input  [31:0] I_13_0_1_1,
  input  [31:0] I_13_0_1_2,
  input  [31:0] I_13_0_2_0,
  input  [31:0] I_13_0_2_1,
  input  [31:0] I_13_0_2_2,
  input  [31:0] I_14_0_0_0,
  input  [31:0] I_14_0_0_1,
  input  [31:0] I_14_0_0_2,
  input  [31:0] I_14_0_1_0,
  input  [31:0] I_14_0_1_1,
  input  [31:0] I_14_0_1_2,
  input  [31:0] I_14_0_2_0,
  input  [31:0] I_14_0_2_1,
  input  [31:0] I_14_0_2_2,
  input  [31:0] I_15_0_0_0,
  input  [31:0] I_15_0_0_1,
  input  [31:0] I_15_0_0_2,
  input  [31:0] I_15_0_1_0,
  input  [31:0] I_15_0_1_1,
  input  [31:0] I_15_0_1_2,
  input  [31:0] I_15_0_2_0,
  input  [31:0] I_15_0_2_1,
  input  [31:0] I_15_0_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_8_2_0,
  output [31:0] O_8_2_1,
  output [31:0] O_8_2_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_9_2_0,
  output [31:0] O_9_2_1,
  output [31:0] O_9_2_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_10_2_0,
  output [31:0] O_10_2_1,
  output [31:0] O_10_2_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_11_2_0,
  output [31:0] O_11_2_1,
  output [31:0] O_11_2_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_12_2_0,
  output [31:0] O_12_2_1,
  output [31:0] O_12_2_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_13_2_0,
  output [31:0] O_13_2_1,
  output [31:0] O_13_2_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_14_2_0,
  output [31:0] O_14_2_1,
  output [31:0] O_14_2_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2,
  output [31:0] O_15_2_0,
  output [31:0] O_15_2_1,
  output [31:0] O_15_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .I_8_0_0_0(op_I_8_0_0_0),
    .I_8_0_0_1(op_I_8_0_0_1),
    .I_8_0_0_2(op_I_8_0_0_2),
    .I_8_0_1_0(op_I_8_0_1_0),
    .I_8_0_1_1(op_I_8_0_1_1),
    .I_8_0_1_2(op_I_8_0_1_2),
    .I_8_0_2_0(op_I_8_0_2_0),
    .I_8_0_2_1(op_I_8_0_2_1),
    .I_8_0_2_2(op_I_8_0_2_2),
    .I_9_0_0_0(op_I_9_0_0_0),
    .I_9_0_0_1(op_I_9_0_0_1),
    .I_9_0_0_2(op_I_9_0_0_2),
    .I_9_0_1_0(op_I_9_0_1_0),
    .I_9_0_1_1(op_I_9_0_1_1),
    .I_9_0_1_2(op_I_9_0_1_2),
    .I_9_0_2_0(op_I_9_0_2_0),
    .I_9_0_2_1(op_I_9_0_2_1),
    .I_9_0_2_2(op_I_9_0_2_2),
    .I_10_0_0_0(op_I_10_0_0_0),
    .I_10_0_0_1(op_I_10_0_0_1),
    .I_10_0_0_2(op_I_10_0_0_2),
    .I_10_0_1_0(op_I_10_0_1_0),
    .I_10_0_1_1(op_I_10_0_1_1),
    .I_10_0_1_2(op_I_10_0_1_2),
    .I_10_0_2_0(op_I_10_0_2_0),
    .I_10_0_2_1(op_I_10_0_2_1),
    .I_10_0_2_2(op_I_10_0_2_2),
    .I_11_0_0_0(op_I_11_0_0_0),
    .I_11_0_0_1(op_I_11_0_0_1),
    .I_11_0_0_2(op_I_11_0_0_2),
    .I_11_0_1_0(op_I_11_0_1_0),
    .I_11_0_1_1(op_I_11_0_1_1),
    .I_11_0_1_2(op_I_11_0_1_2),
    .I_11_0_2_0(op_I_11_0_2_0),
    .I_11_0_2_1(op_I_11_0_2_1),
    .I_11_0_2_2(op_I_11_0_2_2),
    .I_12_0_0_0(op_I_12_0_0_0),
    .I_12_0_0_1(op_I_12_0_0_1),
    .I_12_0_0_2(op_I_12_0_0_2),
    .I_12_0_1_0(op_I_12_0_1_0),
    .I_12_0_1_1(op_I_12_0_1_1),
    .I_12_0_1_2(op_I_12_0_1_2),
    .I_12_0_2_0(op_I_12_0_2_0),
    .I_12_0_2_1(op_I_12_0_2_1),
    .I_12_0_2_2(op_I_12_0_2_2),
    .I_13_0_0_0(op_I_13_0_0_0),
    .I_13_0_0_1(op_I_13_0_0_1),
    .I_13_0_0_2(op_I_13_0_0_2),
    .I_13_0_1_0(op_I_13_0_1_0),
    .I_13_0_1_1(op_I_13_0_1_1),
    .I_13_0_1_2(op_I_13_0_1_2),
    .I_13_0_2_0(op_I_13_0_2_0),
    .I_13_0_2_1(op_I_13_0_2_1),
    .I_13_0_2_2(op_I_13_0_2_2),
    .I_14_0_0_0(op_I_14_0_0_0),
    .I_14_0_0_1(op_I_14_0_0_1),
    .I_14_0_0_2(op_I_14_0_0_2),
    .I_14_0_1_0(op_I_14_0_1_0),
    .I_14_0_1_1(op_I_14_0_1_1),
    .I_14_0_1_2(op_I_14_0_1_2),
    .I_14_0_2_0(op_I_14_0_2_0),
    .I_14_0_2_1(op_I_14_0_2_1),
    .I_14_0_2_2(op_I_14_0_2_2),
    .I_15_0_0_0(op_I_15_0_0_0),
    .I_15_0_0_1(op_I_15_0_0_1),
    .I_15_0_0_2(op_I_15_0_0_2),
    .I_15_0_1_0(op_I_15_0_1_0),
    .I_15_0_1_1(op_I_15_0_1_1),
    .I_15_0_1_2(op_I_15_0_1_2),
    .I_15_0_2_0(op_I_15_0_2_0),
    .I_15_0_2_1(op_I_15_0_2_1),
    .I_15_0_2_2(op_I_15_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_8_1_0 = op_O_8_1_0; // @[MapT.scala 15:7]
  assign O_8_1_1 = op_O_8_1_1; // @[MapT.scala 15:7]
  assign O_8_1_2 = op_O_8_1_2; // @[MapT.scala 15:7]
  assign O_8_2_0 = op_O_8_2_0; // @[MapT.scala 15:7]
  assign O_8_2_1 = op_O_8_2_1; // @[MapT.scala 15:7]
  assign O_8_2_2 = op_O_8_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_9_1_0 = op_O_9_1_0; // @[MapT.scala 15:7]
  assign O_9_1_1 = op_O_9_1_1; // @[MapT.scala 15:7]
  assign O_9_1_2 = op_O_9_1_2; // @[MapT.scala 15:7]
  assign O_9_2_0 = op_O_9_2_0; // @[MapT.scala 15:7]
  assign O_9_2_1 = op_O_9_2_1; // @[MapT.scala 15:7]
  assign O_9_2_2 = op_O_9_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_10_1_0 = op_O_10_1_0; // @[MapT.scala 15:7]
  assign O_10_1_1 = op_O_10_1_1; // @[MapT.scala 15:7]
  assign O_10_1_2 = op_O_10_1_2; // @[MapT.scala 15:7]
  assign O_10_2_0 = op_O_10_2_0; // @[MapT.scala 15:7]
  assign O_10_2_1 = op_O_10_2_1; // @[MapT.scala 15:7]
  assign O_10_2_2 = op_O_10_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_11_1_0 = op_O_11_1_0; // @[MapT.scala 15:7]
  assign O_11_1_1 = op_O_11_1_1; // @[MapT.scala 15:7]
  assign O_11_1_2 = op_O_11_1_2; // @[MapT.scala 15:7]
  assign O_11_2_0 = op_O_11_2_0; // @[MapT.scala 15:7]
  assign O_11_2_1 = op_O_11_2_1; // @[MapT.scala 15:7]
  assign O_11_2_2 = op_O_11_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_12_1_0 = op_O_12_1_0; // @[MapT.scala 15:7]
  assign O_12_1_1 = op_O_12_1_1; // @[MapT.scala 15:7]
  assign O_12_1_2 = op_O_12_1_2; // @[MapT.scala 15:7]
  assign O_12_2_0 = op_O_12_2_0; // @[MapT.scala 15:7]
  assign O_12_2_1 = op_O_12_2_1; // @[MapT.scala 15:7]
  assign O_12_2_2 = op_O_12_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_13_1_0 = op_O_13_1_0; // @[MapT.scala 15:7]
  assign O_13_1_1 = op_O_13_1_1; // @[MapT.scala 15:7]
  assign O_13_1_2 = op_O_13_1_2; // @[MapT.scala 15:7]
  assign O_13_2_0 = op_O_13_2_0; // @[MapT.scala 15:7]
  assign O_13_2_1 = op_O_13_2_1; // @[MapT.scala 15:7]
  assign O_13_2_2 = op_O_13_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_14_1_0 = op_O_14_1_0; // @[MapT.scala 15:7]
  assign O_14_1_1 = op_O_14_1_1; // @[MapT.scala 15:7]
  assign O_14_1_2 = op_O_14_1_2; // @[MapT.scala 15:7]
  assign O_14_2_0 = op_O_14_2_0; // @[MapT.scala 15:7]
  assign O_14_2_1 = op_O_14_2_1; // @[MapT.scala 15:7]
  assign O_14_2_2 = op_O_14_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign O_15_1_0 = op_O_15_1_0; // @[MapT.scala 15:7]
  assign O_15_1_1 = op_O_15_1_1; // @[MapT.scala 15:7]
  assign O_15_1_2 = op_O_15_1_2; // @[MapT.scala 15:7]
  assign O_15_2_0 = op_O_15_2_0; // @[MapT.scala 15:7]
  assign O_15_2_1 = op_O_15_2_1; // @[MapT.scala 15:7]
  assign O_15_2_2 = op_O_15_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0_0 = I_8_0_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_0_1 = I_8_0_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0_2 = I_8_0_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_1_0 = I_8_0_1_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1_1 = I_8_0_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_1_2 = I_8_0_1_2; // @[MapT.scala 14:10]
  assign op_I_8_0_2_0 = I_8_0_2_0; // @[MapT.scala 14:10]
  assign op_I_8_0_2_1 = I_8_0_2_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2_2 = I_8_0_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0_0 = I_9_0_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_0_1 = I_9_0_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0_2 = I_9_0_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_1_0 = I_9_0_1_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1_1 = I_9_0_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_1_2 = I_9_0_1_2; // @[MapT.scala 14:10]
  assign op_I_9_0_2_0 = I_9_0_2_0; // @[MapT.scala 14:10]
  assign op_I_9_0_2_1 = I_9_0_2_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2_2 = I_9_0_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0_0 = I_10_0_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_0_1 = I_10_0_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0_2 = I_10_0_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_1_0 = I_10_0_1_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1_1 = I_10_0_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_1_2 = I_10_0_1_2; // @[MapT.scala 14:10]
  assign op_I_10_0_2_0 = I_10_0_2_0; // @[MapT.scala 14:10]
  assign op_I_10_0_2_1 = I_10_0_2_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2_2 = I_10_0_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0_0 = I_11_0_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_0_1 = I_11_0_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0_2 = I_11_0_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_1_0 = I_11_0_1_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1_1 = I_11_0_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_1_2 = I_11_0_1_2; // @[MapT.scala 14:10]
  assign op_I_11_0_2_0 = I_11_0_2_0; // @[MapT.scala 14:10]
  assign op_I_11_0_2_1 = I_11_0_2_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2_2 = I_11_0_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0_0 = I_12_0_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_0_1 = I_12_0_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0_2 = I_12_0_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_1_0 = I_12_0_1_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1_1 = I_12_0_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_1_2 = I_12_0_1_2; // @[MapT.scala 14:10]
  assign op_I_12_0_2_0 = I_12_0_2_0; // @[MapT.scala 14:10]
  assign op_I_12_0_2_1 = I_12_0_2_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2_2 = I_12_0_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0_0 = I_13_0_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_0_1 = I_13_0_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0_2 = I_13_0_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_1_0 = I_13_0_1_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1_1 = I_13_0_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_1_2 = I_13_0_1_2; // @[MapT.scala 14:10]
  assign op_I_13_0_2_0 = I_13_0_2_0; // @[MapT.scala 14:10]
  assign op_I_13_0_2_1 = I_13_0_2_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2_2 = I_13_0_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0_0 = I_14_0_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_0_1 = I_14_0_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0_2 = I_14_0_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_1_0 = I_14_0_1_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1_1 = I_14_0_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_1_2 = I_14_0_1_2; // @[MapT.scala 14:10]
  assign op_I_14_0_2_0 = I_14_0_2_0; // @[MapT.scala 14:10]
  assign op_I_14_0_2_1 = I_14_0_2_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2_2 = I_14_0_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0_0 = I_15_0_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_0_1 = I_15_0_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0_2 = I_15_0_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_1_0 = I_15_0_1_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1_1 = I_15_0_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_1_2 = I_15_0_1_2; // @[MapT.scala 14:10]
  assign op_I_15_0_2_0 = I_15_0_2_0; // @[MapT.scala 14:10]
  assign op_I_15_0_2_1 = I_15_0_2_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2_2 = I_15_0_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_8_1_0,
  input  [31:0] I_8_1_1,
  input  [31:0] I_8_1_2,
  input  [31:0] I_8_2_0,
  input  [31:0] I_8_2_1,
  input  [31:0] I_8_2_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_9_1_0,
  input  [31:0] I_9_1_1,
  input  [31:0] I_9_1_2,
  input  [31:0] I_9_2_0,
  input  [31:0] I_9_2_1,
  input  [31:0] I_9_2_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_10_1_0,
  input  [31:0] I_10_1_1,
  input  [31:0] I_10_1_2,
  input  [31:0] I_10_2_0,
  input  [31:0] I_10_2_1,
  input  [31:0] I_10_2_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_11_1_0,
  input  [31:0] I_11_1_1,
  input  [31:0] I_11_1_2,
  input  [31:0] I_11_2_0,
  input  [31:0] I_11_2_1,
  input  [31:0] I_11_2_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_12_1_0,
  input  [31:0] I_12_1_1,
  input  [31:0] I_12_1_2,
  input  [31:0] I_12_2_0,
  input  [31:0] I_12_2_1,
  input  [31:0] I_12_2_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_13_1_0,
  input  [31:0] I_13_1_1,
  input  [31:0] I_13_1_2,
  input  [31:0] I_13_2_0,
  input  [31:0] I_13_2_1,
  input  [31:0] I_13_2_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_14_1_0,
  input  [31:0] I_14_1_1,
  input  [31:0] I_14_1_2,
  input  [31:0] I_14_2_0,
  input  [31:0] I_14_2_1,
  input  [31:0] I_14_2_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  input  [31:0] I_15_1_0,
  input  [31:0] I_15_1_1,
  input  [31:0] I_15_1_2,
  input  [31:0] I_15_2_0,
  input  [31:0] I_15_2_1,
  input  [31:0] I_15_2_2,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_1_0,
  output [31:0] O_0_1_1,
  output [31:0] O_0_1_2,
  output [31:0] O_0_2_0,
  output [31:0] O_0_2_1,
  output [31:0] O_0_2_2,
  output [31:0] O_1_0_0,
  output [31:0] O_1_0_1,
  output [31:0] O_1_0_2,
  output [31:0] O_1_1_0,
  output [31:0] O_1_1_1,
  output [31:0] O_1_1_2,
  output [31:0] O_1_2_0,
  output [31:0] O_1_2_1,
  output [31:0] O_1_2_2,
  output [31:0] O_2_0_0,
  output [31:0] O_2_0_1,
  output [31:0] O_2_0_2,
  output [31:0] O_2_1_0,
  output [31:0] O_2_1_1,
  output [31:0] O_2_1_2,
  output [31:0] O_2_2_0,
  output [31:0] O_2_2_1,
  output [31:0] O_2_2_2,
  output [31:0] O_3_0_0,
  output [31:0] O_3_0_1,
  output [31:0] O_3_0_2,
  output [31:0] O_3_1_0,
  output [31:0] O_3_1_1,
  output [31:0] O_3_1_2,
  output [31:0] O_3_2_0,
  output [31:0] O_3_2_1,
  output [31:0] O_3_2_2,
  output [31:0] O_4_0_0,
  output [31:0] O_4_0_1,
  output [31:0] O_4_0_2,
  output [31:0] O_4_1_0,
  output [31:0] O_4_1_1,
  output [31:0] O_4_1_2,
  output [31:0] O_4_2_0,
  output [31:0] O_4_2_1,
  output [31:0] O_4_2_2,
  output [31:0] O_5_0_0,
  output [31:0] O_5_0_1,
  output [31:0] O_5_0_2,
  output [31:0] O_5_1_0,
  output [31:0] O_5_1_1,
  output [31:0] O_5_1_2,
  output [31:0] O_5_2_0,
  output [31:0] O_5_2_1,
  output [31:0] O_5_2_2,
  output [31:0] O_6_0_0,
  output [31:0] O_6_0_1,
  output [31:0] O_6_0_2,
  output [31:0] O_6_1_0,
  output [31:0] O_6_1_1,
  output [31:0] O_6_1_2,
  output [31:0] O_6_2_0,
  output [31:0] O_6_2_1,
  output [31:0] O_6_2_2,
  output [31:0] O_7_0_0,
  output [31:0] O_7_0_1,
  output [31:0] O_7_0_2,
  output [31:0] O_7_1_0,
  output [31:0] O_7_1_1,
  output [31:0] O_7_1_2,
  output [31:0] O_7_2_0,
  output [31:0] O_7_2_1,
  output [31:0] O_7_2_2,
  output [31:0] O_8_0_0,
  output [31:0] O_8_0_1,
  output [31:0] O_8_0_2,
  output [31:0] O_8_1_0,
  output [31:0] O_8_1_1,
  output [31:0] O_8_1_2,
  output [31:0] O_8_2_0,
  output [31:0] O_8_2_1,
  output [31:0] O_8_2_2,
  output [31:0] O_9_0_0,
  output [31:0] O_9_0_1,
  output [31:0] O_9_0_2,
  output [31:0] O_9_1_0,
  output [31:0] O_9_1_1,
  output [31:0] O_9_1_2,
  output [31:0] O_9_2_0,
  output [31:0] O_9_2_1,
  output [31:0] O_9_2_2,
  output [31:0] O_10_0_0,
  output [31:0] O_10_0_1,
  output [31:0] O_10_0_2,
  output [31:0] O_10_1_0,
  output [31:0] O_10_1_1,
  output [31:0] O_10_1_2,
  output [31:0] O_10_2_0,
  output [31:0] O_10_2_1,
  output [31:0] O_10_2_2,
  output [31:0] O_11_0_0,
  output [31:0] O_11_0_1,
  output [31:0] O_11_0_2,
  output [31:0] O_11_1_0,
  output [31:0] O_11_1_1,
  output [31:0] O_11_1_2,
  output [31:0] O_11_2_0,
  output [31:0] O_11_2_1,
  output [31:0] O_11_2_2,
  output [31:0] O_12_0_0,
  output [31:0] O_12_0_1,
  output [31:0] O_12_0_2,
  output [31:0] O_12_1_0,
  output [31:0] O_12_1_1,
  output [31:0] O_12_1_2,
  output [31:0] O_12_2_0,
  output [31:0] O_12_2_1,
  output [31:0] O_12_2_2,
  output [31:0] O_13_0_0,
  output [31:0] O_13_0_1,
  output [31:0] O_13_0_2,
  output [31:0] O_13_1_0,
  output [31:0] O_13_1_1,
  output [31:0] O_13_1_2,
  output [31:0] O_13_2_0,
  output [31:0] O_13_2_1,
  output [31:0] O_13_2_2,
  output [31:0] O_14_0_0,
  output [31:0] O_14_0_1,
  output [31:0] O_14_0_2,
  output [31:0] O_14_1_0,
  output [31:0] O_14_1_1,
  output [31:0] O_14_1_2,
  output [31:0] O_14_2_0,
  output [31:0] O_14_2_1,
  output [31:0] O_14_2_2,
  output [31:0] O_15_0_0,
  output [31:0] O_15_0_1,
  output [31:0] O_15_0_2,
  output [31:0] O_15_1_0,
  output [31:0] O_15_1_1,
  output [31:0] O_15_1_2,
  output [31:0] O_15_2_0,
  output [31:0] O_15_2_1,
  output [31:0] O_15_2_2
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_0_0_1 = I_0_0_1; // @[Passthrough.scala 17:68]
  assign O_0_0_2 = I_0_0_2; // @[Passthrough.scala 17:68]
  assign O_0_1_0 = I_0_1_0; // @[Passthrough.scala 17:68]
  assign O_0_1_1 = I_0_1_1; // @[Passthrough.scala 17:68]
  assign O_0_1_2 = I_0_1_2; // @[Passthrough.scala 17:68]
  assign O_0_2_0 = I_0_2_0; // @[Passthrough.scala 17:68]
  assign O_0_2_1 = I_0_2_1; // @[Passthrough.scala 17:68]
  assign O_0_2_2 = I_0_2_2; // @[Passthrough.scala 17:68]
  assign O_1_0_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0_1 = I_1_0_1; // @[Passthrough.scala 17:68]
  assign O_1_0_2 = I_1_0_2; // @[Passthrough.scala 17:68]
  assign O_1_1_0 = I_1_1_0; // @[Passthrough.scala 17:68]
  assign O_1_1_1 = I_1_1_1; // @[Passthrough.scala 17:68]
  assign O_1_1_2 = I_1_1_2; // @[Passthrough.scala 17:68]
  assign O_1_2_0 = I_1_2_0; // @[Passthrough.scala 17:68]
  assign O_1_2_1 = I_1_2_1; // @[Passthrough.scala 17:68]
  assign O_1_2_2 = I_1_2_2; // @[Passthrough.scala 17:68]
  assign O_2_0_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0_1 = I_2_0_1; // @[Passthrough.scala 17:68]
  assign O_2_0_2 = I_2_0_2; // @[Passthrough.scala 17:68]
  assign O_2_1_0 = I_2_1_0; // @[Passthrough.scala 17:68]
  assign O_2_1_1 = I_2_1_1; // @[Passthrough.scala 17:68]
  assign O_2_1_2 = I_2_1_2; // @[Passthrough.scala 17:68]
  assign O_2_2_0 = I_2_2_0; // @[Passthrough.scala 17:68]
  assign O_2_2_1 = I_2_2_1; // @[Passthrough.scala 17:68]
  assign O_2_2_2 = I_2_2_2; // @[Passthrough.scala 17:68]
  assign O_3_0_0 = I_3_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0_1 = I_3_0_1; // @[Passthrough.scala 17:68]
  assign O_3_0_2 = I_3_0_2; // @[Passthrough.scala 17:68]
  assign O_3_1_0 = I_3_1_0; // @[Passthrough.scala 17:68]
  assign O_3_1_1 = I_3_1_1; // @[Passthrough.scala 17:68]
  assign O_3_1_2 = I_3_1_2; // @[Passthrough.scala 17:68]
  assign O_3_2_0 = I_3_2_0; // @[Passthrough.scala 17:68]
  assign O_3_2_1 = I_3_2_1; // @[Passthrough.scala 17:68]
  assign O_3_2_2 = I_3_2_2; // @[Passthrough.scala 17:68]
  assign O_4_0_0 = I_4_0_0; // @[Passthrough.scala 17:68]
  assign O_4_0_1 = I_4_0_1; // @[Passthrough.scala 17:68]
  assign O_4_0_2 = I_4_0_2; // @[Passthrough.scala 17:68]
  assign O_4_1_0 = I_4_1_0; // @[Passthrough.scala 17:68]
  assign O_4_1_1 = I_4_1_1; // @[Passthrough.scala 17:68]
  assign O_4_1_2 = I_4_1_2; // @[Passthrough.scala 17:68]
  assign O_4_2_0 = I_4_2_0; // @[Passthrough.scala 17:68]
  assign O_4_2_1 = I_4_2_1; // @[Passthrough.scala 17:68]
  assign O_4_2_2 = I_4_2_2; // @[Passthrough.scala 17:68]
  assign O_5_0_0 = I_5_0_0; // @[Passthrough.scala 17:68]
  assign O_5_0_1 = I_5_0_1; // @[Passthrough.scala 17:68]
  assign O_5_0_2 = I_5_0_2; // @[Passthrough.scala 17:68]
  assign O_5_1_0 = I_5_1_0; // @[Passthrough.scala 17:68]
  assign O_5_1_1 = I_5_1_1; // @[Passthrough.scala 17:68]
  assign O_5_1_2 = I_5_1_2; // @[Passthrough.scala 17:68]
  assign O_5_2_0 = I_5_2_0; // @[Passthrough.scala 17:68]
  assign O_5_2_1 = I_5_2_1; // @[Passthrough.scala 17:68]
  assign O_5_2_2 = I_5_2_2; // @[Passthrough.scala 17:68]
  assign O_6_0_0 = I_6_0_0; // @[Passthrough.scala 17:68]
  assign O_6_0_1 = I_6_0_1; // @[Passthrough.scala 17:68]
  assign O_6_0_2 = I_6_0_2; // @[Passthrough.scala 17:68]
  assign O_6_1_0 = I_6_1_0; // @[Passthrough.scala 17:68]
  assign O_6_1_1 = I_6_1_1; // @[Passthrough.scala 17:68]
  assign O_6_1_2 = I_6_1_2; // @[Passthrough.scala 17:68]
  assign O_6_2_0 = I_6_2_0; // @[Passthrough.scala 17:68]
  assign O_6_2_1 = I_6_2_1; // @[Passthrough.scala 17:68]
  assign O_6_2_2 = I_6_2_2; // @[Passthrough.scala 17:68]
  assign O_7_0_0 = I_7_0_0; // @[Passthrough.scala 17:68]
  assign O_7_0_1 = I_7_0_1; // @[Passthrough.scala 17:68]
  assign O_7_0_2 = I_7_0_2; // @[Passthrough.scala 17:68]
  assign O_7_1_0 = I_7_1_0; // @[Passthrough.scala 17:68]
  assign O_7_1_1 = I_7_1_1; // @[Passthrough.scala 17:68]
  assign O_7_1_2 = I_7_1_2; // @[Passthrough.scala 17:68]
  assign O_7_2_0 = I_7_2_0; // @[Passthrough.scala 17:68]
  assign O_7_2_1 = I_7_2_1; // @[Passthrough.scala 17:68]
  assign O_7_2_2 = I_7_2_2; // @[Passthrough.scala 17:68]
  assign O_8_0_0 = I_8_0_0; // @[Passthrough.scala 17:68]
  assign O_8_0_1 = I_8_0_1; // @[Passthrough.scala 17:68]
  assign O_8_0_2 = I_8_0_2; // @[Passthrough.scala 17:68]
  assign O_8_1_0 = I_8_1_0; // @[Passthrough.scala 17:68]
  assign O_8_1_1 = I_8_1_1; // @[Passthrough.scala 17:68]
  assign O_8_1_2 = I_8_1_2; // @[Passthrough.scala 17:68]
  assign O_8_2_0 = I_8_2_0; // @[Passthrough.scala 17:68]
  assign O_8_2_1 = I_8_2_1; // @[Passthrough.scala 17:68]
  assign O_8_2_2 = I_8_2_2; // @[Passthrough.scala 17:68]
  assign O_9_0_0 = I_9_0_0; // @[Passthrough.scala 17:68]
  assign O_9_0_1 = I_9_0_1; // @[Passthrough.scala 17:68]
  assign O_9_0_2 = I_9_0_2; // @[Passthrough.scala 17:68]
  assign O_9_1_0 = I_9_1_0; // @[Passthrough.scala 17:68]
  assign O_9_1_1 = I_9_1_1; // @[Passthrough.scala 17:68]
  assign O_9_1_2 = I_9_1_2; // @[Passthrough.scala 17:68]
  assign O_9_2_0 = I_9_2_0; // @[Passthrough.scala 17:68]
  assign O_9_2_1 = I_9_2_1; // @[Passthrough.scala 17:68]
  assign O_9_2_2 = I_9_2_2; // @[Passthrough.scala 17:68]
  assign O_10_0_0 = I_10_0_0; // @[Passthrough.scala 17:68]
  assign O_10_0_1 = I_10_0_1; // @[Passthrough.scala 17:68]
  assign O_10_0_2 = I_10_0_2; // @[Passthrough.scala 17:68]
  assign O_10_1_0 = I_10_1_0; // @[Passthrough.scala 17:68]
  assign O_10_1_1 = I_10_1_1; // @[Passthrough.scala 17:68]
  assign O_10_1_2 = I_10_1_2; // @[Passthrough.scala 17:68]
  assign O_10_2_0 = I_10_2_0; // @[Passthrough.scala 17:68]
  assign O_10_2_1 = I_10_2_1; // @[Passthrough.scala 17:68]
  assign O_10_2_2 = I_10_2_2; // @[Passthrough.scala 17:68]
  assign O_11_0_0 = I_11_0_0; // @[Passthrough.scala 17:68]
  assign O_11_0_1 = I_11_0_1; // @[Passthrough.scala 17:68]
  assign O_11_0_2 = I_11_0_2; // @[Passthrough.scala 17:68]
  assign O_11_1_0 = I_11_1_0; // @[Passthrough.scala 17:68]
  assign O_11_1_1 = I_11_1_1; // @[Passthrough.scala 17:68]
  assign O_11_1_2 = I_11_1_2; // @[Passthrough.scala 17:68]
  assign O_11_2_0 = I_11_2_0; // @[Passthrough.scala 17:68]
  assign O_11_2_1 = I_11_2_1; // @[Passthrough.scala 17:68]
  assign O_11_2_2 = I_11_2_2; // @[Passthrough.scala 17:68]
  assign O_12_0_0 = I_12_0_0; // @[Passthrough.scala 17:68]
  assign O_12_0_1 = I_12_0_1; // @[Passthrough.scala 17:68]
  assign O_12_0_2 = I_12_0_2; // @[Passthrough.scala 17:68]
  assign O_12_1_0 = I_12_1_0; // @[Passthrough.scala 17:68]
  assign O_12_1_1 = I_12_1_1; // @[Passthrough.scala 17:68]
  assign O_12_1_2 = I_12_1_2; // @[Passthrough.scala 17:68]
  assign O_12_2_0 = I_12_2_0; // @[Passthrough.scala 17:68]
  assign O_12_2_1 = I_12_2_1; // @[Passthrough.scala 17:68]
  assign O_12_2_2 = I_12_2_2; // @[Passthrough.scala 17:68]
  assign O_13_0_0 = I_13_0_0; // @[Passthrough.scala 17:68]
  assign O_13_0_1 = I_13_0_1; // @[Passthrough.scala 17:68]
  assign O_13_0_2 = I_13_0_2; // @[Passthrough.scala 17:68]
  assign O_13_1_0 = I_13_1_0; // @[Passthrough.scala 17:68]
  assign O_13_1_1 = I_13_1_1; // @[Passthrough.scala 17:68]
  assign O_13_1_2 = I_13_1_2; // @[Passthrough.scala 17:68]
  assign O_13_2_0 = I_13_2_0; // @[Passthrough.scala 17:68]
  assign O_13_2_1 = I_13_2_1; // @[Passthrough.scala 17:68]
  assign O_13_2_2 = I_13_2_2; // @[Passthrough.scala 17:68]
  assign O_14_0_0 = I_14_0_0; // @[Passthrough.scala 17:68]
  assign O_14_0_1 = I_14_0_1; // @[Passthrough.scala 17:68]
  assign O_14_0_2 = I_14_0_2; // @[Passthrough.scala 17:68]
  assign O_14_1_0 = I_14_1_0; // @[Passthrough.scala 17:68]
  assign O_14_1_1 = I_14_1_1; // @[Passthrough.scala 17:68]
  assign O_14_1_2 = I_14_1_2; // @[Passthrough.scala 17:68]
  assign O_14_2_0 = I_14_2_0; // @[Passthrough.scala 17:68]
  assign O_14_2_1 = I_14_2_1; // @[Passthrough.scala 17:68]
  assign O_14_2_2 = I_14_2_2; // @[Passthrough.scala 17:68]
  assign O_15_0_0 = I_15_0_0; // @[Passthrough.scala 17:68]
  assign O_15_0_1 = I_15_0_1; // @[Passthrough.scala 17:68]
  assign O_15_0_2 = I_15_0_2; // @[Passthrough.scala 17:68]
  assign O_15_1_0 = I_15_1_0; // @[Passthrough.scala 17:68]
  assign O_15_1_1 = I_15_1_1; // @[Passthrough.scala 17:68]
  assign O_15_1_2 = I_15_1_2; // @[Passthrough.scala 17:68]
  assign O_15_2_0 = I_15_2_0; // @[Passthrough.scala 17:68]
  assign O_15_2_1 = I_15_2_1; // @[Passthrough.scala 17:68]
  assign O_15_2_2 = I_15_2_2; // @[Passthrough.scala 17:68]
endmodule
module Counter_T(
  input         clock,
  input         reset,
  output [31:0] O
);
  reg [31:0] counter_value; // @[Counter.scala 53:30]
  reg [31:0] _RAND_0;
  wire  _T; // @[Counter.scala 61:49]
  wire [31:0] _T_3; // @[Counter.scala 63:70]
  assign _T = counter_value == 32'hef0; // @[Counter.scala 61:49]
  assign _T_3 = counter_value + 32'h10; // @[Counter.scala 63:70]
  assign O = counter_value; // @[Counter.scala 66:5]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counter_value = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      counter_value <= 32'h0;
    end else if (_T) begin
      counter_value <= 32'h0;
    end else begin
      counter_value <= _T_3;
    end
  end
endmodule
module Counter_TS(
  input         clock,
  input         reset,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3,
  output [31:0] O_4,
  output [31:0] O_5,
  output [31:0] O_6,
  output [31:0] O_7,
  output [31:0] O_8,
  output [31:0] O_9,
  output [31:0] O_10,
  output [31:0] O_11,
  output [31:0] O_12,
  output [31:0] O_13,
  output [31:0] O_14,
  output [31:0] O_15
);
  wire  counter_t_clock; // @[Counter.scala 84:25]
  wire  counter_t_reset; // @[Counter.scala 84:25]
  wire [31:0] counter_t_O; // @[Counter.scala 84:25]
  wire [32:0] _T; // @[Counter.scala 95:49]
  Counter_T counter_t ( // @[Counter.scala 84:25]
    .clock(counter_t_clock),
    .reset(counter_t_reset),
    .O(counter_t_O)
  );
  assign _T = {{1'd0}, counter_t_O}; // @[Counter.scala 95:49]
  assign O_0 = _T[31:0]; // @[Counter.scala 95:12]
  assign O_1 = 32'h1 + counter_t_O; // @[Counter.scala 95:12]
  assign O_2 = 32'h2 + counter_t_O; // @[Counter.scala 95:12]
  assign O_3 = 32'h3 + counter_t_O; // @[Counter.scala 95:12]
  assign O_4 = 32'h4 + counter_t_O; // @[Counter.scala 95:12]
  assign O_5 = 32'h5 + counter_t_O; // @[Counter.scala 95:12]
  assign O_6 = 32'h6 + counter_t_O; // @[Counter.scala 95:12]
  assign O_7 = 32'h7 + counter_t_O; // @[Counter.scala 95:12]
  assign O_8 = 32'h8 + counter_t_O; // @[Counter.scala 95:12]
  assign O_9 = 32'h9 + counter_t_O; // @[Counter.scala 95:12]
  assign O_10 = 32'ha + counter_t_O; // @[Counter.scala 95:12]
  assign O_11 = 32'hb + counter_t_O; // @[Counter.scala 95:12]
  assign O_12 = 32'hc + counter_t_O; // @[Counter.scala 95:12]
  assign O_13 = 32'hd + counter_t_O; // @[Counter.scala 95:12]
  assign O_14 = 32'he + counter_t_O; // @[Counter.scala 95:12]
  assign O_15 = 32'hf + counter_t_O; // @[Counter.scala 95:12]
  assign counter_t_clock = clock;
  assign counter_t_reset = reset;
endmodule
module AtomTuple(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1,
  output [31:0] O_t0b,
  output [31:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Lt(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  wire  _T; // @[Arithmetic.scala 462:25]
  assign _T = I_t0b < I_t1b; // @[Arithmetic.scala 462:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 464:14]
  assign O = {{31'd0}, _T}; // @[Arithmetic.scala 462:7]
endmodule
module Not(
  input   valid_up,
  output  valid_down,
  input   I,
  output  O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 45:14]
  assign O = ~I; // @[Arithmetic.scala 44:5]
endmodule
module Module_0(
  output        valid_down,
  input  [31:0] I,
  output        O
);
  wire  n112_valid_up; // @[Top.scala 18:22]
  wire  n112_valid_down; // @[Top.scala 18:22]
  wire [31:0] n112_I0; // @[Top.scala 18:22]
  wire [31:0] n112_I1; // @[Top.scala 18:22]
  wire [31:0] n112_O_t0b; // @[Top.scala 18:22]
  wire [31:0] n112_O_t1b; // @[Top.scala 18:22]
  wire  n113_valid_up; // @[Top.scala 22:22]
  wire  n113_valid_down; // @[Top.scala 22:22]
  wire [31:0] n113_I_t0b; // @[Top.scala 22:22]
  wire [31:0] n113_I_t1b; // @[Top.scala 22:22]
  wire [31:0] n113_O; // @[Top.scala 22:22]
  wire  n114_valid_up; // @[Top.scala 25:22]
  wire  n114_valid_down; // @[Top.scala 25:22]
  wire  n114_I; // @[Top.scala 25:22]
  wire  n114_O; // @[Top.scala 25:22]
  AtomTuple n112 ( // @[Top.scala 18:22]
    .valid_up(n112_valid_up),
    .valid_down(n112_valid_down),
    .I0(n112_I0),
    .I1(n112_I1),
    .O_t0b(n112_O_t0b),
    .O_t1b(n112_O_t1b)
  );
  Lt n113 ( // @[Top.scala 22:22]
    .valid_up(n113_valid_up),
    .valid_down(n113_valid_down),
    .I_t0b(n113_I_t0b),
    .I_t1b(n113_I_t1b),
    .O(n113_O)
  );
  Not n114 ( // @[Top.scala 25:22]
    .valid_up(n114_valid_up),
    .valid_down(n114_valid_down),
    .I(n114_I),
    .O(n114_O)
  );
  assign valid_down = n114_valid_down; // @[Top.scala 29:16]
  assign O = n114_O; // @[Top.scala 28:7]
  assign n112_valid_up = 1'h1; // @[Top.scala 21:19]
  assign n112_I0 = I; // @[Top.scala 19:13]
  assign n112_I1 = 32'h780; // @[Top.scala 20:13]
  assign n113_valid_up = n112_valid_down; // @[Top.scala 24:19]
  assign n113_I_t0b = n112_O_t0b; // @[Top.scala 23:12]
  assign n113_I_t1b = n112_O_t1b; // @[Top.scala 23:12]
  assign n114_valid_up = n113_valid_down; // @[Top.scala 27:19]
  assign n114_I = n113_O[0]; // @[Top.scala 26:12]
endmodule
module MapS_4(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7,
  output        O_8,
  output        O_9,
  output        O_10,
  output        O_11,
  output        O_12,
  output        O_13,
  output        O_14,
  output        O_15
);
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire  other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire  other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I; // @[MapS.scala 10:86]
  wire  other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I; // @[MapS.scala 10:86]
  wire  other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I; // @[MapS.scala 10:86]
  wire  other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I; // @[MapS.scala 10:86]
  wire  other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I; // @[MapS.scala 10:86]
  wire  other_ops_6_O; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I; // @[MapS.scala 10:86]
  wire  other_ops_7_O; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I; // @[MapS.scala 10:86]
  wire  other_ops_8_O; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I; // @[MapS.scala 10:86]
  wire  other_ops_9_O; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I; // @[MapS.scala 10:86]
  wire  other_ops_10_O; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I; // @[MapS.scala 10:86]
  wire  other_ops_11_O; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I; // @[MapS.scala 10:86]
  wire  other_ops_12_O; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I; // @[MapS.scala 10:86]
  wire  other_ops_13_O; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I; // @[MapS.scala 10:86]
  wire  other_ops_14_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_2_valid_down),
    .I(other_ops_2_I),
    .O(other_ops_2_O)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_3_valid_down),
    .I(other_ops_3_I),
    .O(other_ops_3_O)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_4_valid_down),
    .I(other_ops_4_I),
    .O(other_ops_4_O)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_5_valid_down),
    .I(other_ops_5_I),
    .O(other_ops_5_O)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_6_valid_down),
    .I(other_ops_6_I),
    .O(other_ops_6_O)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_7_valid_down),
    .I(other_ops_7_I),
    .O(other_ops_7_O)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_8_valid_down),
    .I(other_ops_8_I),
    .O(other_ops_8_O)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_9_valid_down),
    .I(other_ops_9_I),
    .O(other_ops_9_O)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_10_valid_down),
    .I(other_ops_10_I),
    .O(other_ops_10_O)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_11_valid_down),
    .I(other_ops_11_I),
    .O(other_ops_11_O)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_12_valid_down),
    .I(other_ops_12_I),
    .O(other_ops_12_O)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_13_valid_down),
    .I(other_ops_13_I),
    .O(other_ops_13_O)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_14_valid_down),
    .I(other_ops_14_I),
    .O(other_ops_14_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign O_8 = other_ops_7_O; // @[MapS.scala 21:12]
  assign O_9 = other_ops_8_O; // @[MapS.scala 21:12]
  assign O_10 = other_ops_9_O; // @[MapS.scala 21:12]
  assign O_11 = other_ops_10_O; // @[MapS.scala 21:12]
  assign O_12 = other_ops_11_O; // @[MapS.scala 21:12]
  assign O_13 = other_ops_12_O; // @[MapS.scala 21:12]
  assign O_14 = other_ops_13_O; // @[MapS.scala 21:12]
  assign O_15 = other_ops_14_O; // @[MapS.scala 21:12]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
  assign other_ops_2_I = I_3; // @[MapS.scala 20:41]
  assign other_ops_3_I = I_4; // @[MapS.scala 20:41]
  assign other_ops_4_I = I_5; // @[MapS.scala 20:41]
  assign other_ops_5_I = I_6; // @[MapS.scala 20:41]
  assign other_ops_6_I = I_7; // @[MapS.scala 20:41]
  assign other_ops_7_I = I_8; // @[MapS.scala 20:41]
  assign other_ops_8_I = I_9; // @[MapS.scala 20:41]
  assign other_ops_9_I = I_10; // @[MapS.scala 20:41]
  assign other_ops_10_I = I_11; // @[MapS.scala 20:41]
  assign other_ops_11_I = I_12; // @[MapS.scala 20:41]
  assign other_ops_12_I = I_13; // @[MapS.scala 20:41]
  assign other_ops_13_I = I_14; // @[MapS.scala 20:41]
  assign other_ops_14_I = I_15; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7,
  output        O_8,
  output        O_9,
  output        O_10,
  output        O_11,
  output        O_12,
  output        O_13,
  output        O_14,
  output        O_15
);
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3; // @[MapT.scala 8:20]
  wire [31:0] op_I_4; // @[MapT.scala 8:20]
  wire [31:0] op_I_5; // @[MapT.scala 8:20]
  wire [31:0] op_I_6; // @[MapT.scala 8:20]
  wire [31:0] op_I_7; // @[MapT.scala 8:20]
  wire [31:0] op_I_8; // @[MapT.scala 8:20]
  wire [31:0] op_I_9; // @[MapT.scala 8:20]
  wire [31:0] op_I_10; // @[MapT.scala 8:20]
  wire [31:0] op_I_11; // @[MapT.scala 8:20]
  wire [31:0] op_I_12; // @[MapT.scala 8:20]
  wire [31:0] op_I_13; // @[MapT.scala 8:20]
  wire [31:0] op_I_14; // @[MapT.scala 8:20]
  wire [31:0] op_I_15; // @[MapT.scala 8:20]
  wire  op_O_0; // @[MapT.scala 8:20]
  wire  op_O_1; // @[MapT.scala 8:20]
  wire  op_O_2; // @[MapT.scala 8:20]
  wire  op_O_3; // @[MapT.scala 8:20]
  wire  op_O_4; // @[MapT.scala 8:20]
  wire  op_O_5; // @[MapT.scala 8:20]
  wire  op_O_6; // @[MapT.scala 8:20]
  wire  op_O_7; // @[MapT.scala 8:20]
  wire  op_O_8; // @[MapT.scala 8:20]
  wire  op_O_9; // @[MapT.scala 8:20]
  wire  op_O_10; // @[MapT.scala 8:20]
  wire  op_O_11; // @[MapT.scala 8:20]
  wire  op_O_12; // @[MapT.scala 8:20]
  wire  op_O_13; // @[MapT.scala 8:20]
  wire  op_O_14; // @[MapT.scala 8:20]
  wire  op_O_15; // @[MapT.scala 8:20]
  MapS_4 op ( // @[MapT.scala 8:20]
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .I_3(op_I_3),
    .I_4(op_I_4),
    .I_5(op_I_5),
    .I_6(op_I_6),
    .I_7(op_I_7),
    .I_8(op_I_8),
    .I_9(op_I_9),
    .I_10(op_I_10),
    .I_11(op_I_11),
    .I_12(op_I_12),
    .I_13(op_I_13),
    .I_14(op_I_14),
    .I_15(op_I_15),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7),
    .O_8(op_O_8),
    .O_9(op_O_9),
    .O_10(op_O_10),
    .O_11(op_O_11),
    .O_12(op_O_12),
    .O_13(op_O_13),
    .O_14(op_O_14),
    .O_15(op_O_15)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign O_8 = op_O_8; // @[MapT.scala 15:7]
  assign O_9 = op_O_9; // @[MapT.scala 15:7]
  assign O_10 = op_O_10; // @[MapT.scala 15:7]
  assign O_11 = op_O_11; // @[MapT.scala 15:7]
  assign O_12 = op_O_12; // @[MapT.scala 15:7]
  assign O_13 = op_O_13; // @[MapT.scala 15:7]
  assign O_14 = op_O_14; // @[MapT.scala 15:7]
  assign O_15 = op_O_15; // @[MapT.scala 15:7]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
  assign op_I_3 = I_3; // @[MapT.scala 14:10]
  assign op_I_4 = I_4; // @[MapT.scala 14:10]
  assign op_I_5 = I_5; // @[MapT.scala 14:10]
  assign op_I_6 = I_6; // @[MapT.scala 14:10]
  assign op_I_7 = I_7; // @[MapT.scala 14:10]
  assign op_I_8 = I_8; // @[MapT.scala 14:10]
  assign op_I_9 = I_9; // @[MapT.scala 14:10]
  assign op_I_10 = I_10; // @[MapT.scala 14:10]
  assign op_I_11 = I_11; // @[MapT.scala 14:10]
  assign op_I_12 = I_12; // @[MapT.scala 14:10]
  assign op_I_13 = I_13; // @[MapT.scala 14:10]
  assign op_I_14 = I_14; // @[MapT.scala 14:10]
  assign op_I_15 = I_15; // @[MapT.scala 14:10]
endmodule
module AtomTuple_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [7:0]  I1,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module RShift(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [7:0]  I_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 402:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 400:7]
endmodule
module LShift(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [7:0]  I_t1b,
  output [31:0] O
);
  wire [286:0] _GEN_0; // @[Arithmetic.scala 431:25]
  wire [286:0] _T; // @[Arithmetic.scala 431:25]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 431:25]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 431:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 433:14]
  assign O = _T[31:0]; // @[Arithmetic.scala 431:7]
endmodule
module Eq(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  wire  _T; // @[Arithmetic.scala 494:25]
  assign _T = I_t0b == I_t1b; // @[Arithmetic.scala 494:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 496:14]
  assign O = {{31'd0}, _T}; // @[Arithmetic.scala 494:7]
endmodule
module Module_1(
  output        valid_down,
  input  [31:0] I,
  output        O
);
  wire  n120_valid_up; // @[Top.scala 36:22]
  wire  n120_valid_down; // @[Top.scala 36:22]
  wire [31:0] n120_I0; // @[Top.scala 36:22]
  wire [7:0] n120_I1; // @[Top.scala 36:22]
  wire [31:0] n120_O_t0b; // @[Top.scala 36:22]
  wire [7:0] n120_O_t1b; // @[Top.scala 36:22]
  wire  n121_valid_up; // @[Top.scala 40:22]
  wire  n121_valid_down; // @[Top.scala 40:22]
  wire [31:0] n121_I_t0b; // @[Top.scala 40:22]
  wire [7:0] n121_I_t1b; // @[Top.scala 40:22]
  wire [31:0] n121_O; // @[Top.scala 40:22]
  wire  n122_valid_up; // @[Top.scala 43:22]
  wire  n122_valid_down; // @[Top.scala 43:22]
  wire [31:0] n122_I0; // @[Top.scala 43:22]
  wire [7:0] n122_I1; // @[Top.scala 43:22]
  wire [31:0] n122_O_t0b; // @[Top.scala 43:22]
  wire [7:0] n122_O_t1b; // @[Top.scala 43:22]
  wire  n123_valid_up; // @[Top.scala 47:22]
  wire  n123_valid_down; // @[Top.scala 47:22]
  wire [31:0] n123_I_t0b; // @[Top.scala 47:22]
  wire [7:0] n123_I_t1b; // @[Top.scala 47:22]
  wire [31:0] n123_O; // @[Top.scala 47:22]
  wire  n124_valid_up; // @[Top.scala 50:22]
  wire  n124_valid_down; // @[Top.scala 50:22]
  wire [31:0] n124_I0; // @[Top.scala 50:22]
  wire [31:0] n124_I1; // @[Top.scala 50:22]
  wire [31:0] n124_O_t0b; // @[Top.scala 50:22]
  wire [31:0] n124_O_t1b; // @[Top.scala 50:22]
  wire  n125_valid_up; // @[Top.scala 54:22]
  wire  n125_valid_down; // @[Top.scala 54:22]
  wire [31:0] n125_I_t0b; // @[Top.scala 54:22]
  wire [31:0] n125_I_t1b; // @[Top.scala 54:22]
  wire [31:0] n125_O; // @[Top.scala 54:22]
  wire  n126_valid_up; // @[Top.scala 57:22]
  wire  n126_valid_down; // @[Top.scala 57:22]
  wire  n126_I; // @[Top.scala 57:22]
  wire  n126_O; // @[Top.scala 57:22]
  AtomTuple_1 n120 ( // @[Top.scala 36:22]
    .valid_up(n120_valid_up),
    .valid_down(n120_valid_down),
    .I0(n120_I0),
    .I1(n120_I1),
    .O_t0b(n120_O_t0b),
    .O_t1b(n120_O_t1b)
  );
  RShift n121 ( // @[Top.scala 40:22]
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_t0b(n121_I_t0b),
    .I_t1b(n121_I_t1b),
    .O(n121_O)
  );
  AtomTuple_1 n122 ( // @[Top.scala 43:22]
    .valid_up(n122_valid_up),
    .valid_down(n122_valid_down),
    .I0(n122_I0),
    .I1(n122_I1),
    .O_t0b(n122_O_t0b),
    .O_t1b(n122_O_t1b)
  );
  LShift n123 ( // @[Top.scala 47:22]
    .valid_up(n123_valid_up),
    .valid_down(n123_valid_down),
    .I_t0b(n123_I_t0b),
    .I_t1b(n123_I_t1b),
    .O(n123_O)
  );
  AtomTuple n124 ( // @[Top.scala 50:22]
    .valid_up(n124_valid_up),
    .valid_down(n124_valid_down),
    .I0(n124_I0),
    .I1(n124_I1),
    .O_t0b(n124_O_t0b),
    .O_t1b(n124_O_t1b)
  );
  Eq n125 ( // @[Top.scala 54:22]
    .valid_up(n125_valid_up),
    .valid_down(n125_valid_down),
    .I_t0b(n125_I_t0b),
    .I_t1b(n125_I_t1b),
    .O(n125_O)
  );
  Not n126 ( // @[Top.scala 57:22]
    .valid_up(n126_valid_up),
    .valid_down(n126_valid_down),
    .I(n126_I),
    .O(n126_O)
  );
  assign valid_down = n126_valid_down; // @[Top.scala 61:16]
  assign O = n126_O; // @[Top.scala 60:7]
  assign n120_valid_up = 1'h1; // @[Top.scala 39:19]
  assign n120_I0 = I; // @[Top.scala 37:13]
  assign n120_I1 = 8'h1; // @[Top.scala 38:13]
  assign n121_valid_up = n120_valid_down; // @[Top.scala 42:19]
  assign n121_I_t0b = n120_O_t0b; // @[Top.scala 41:12]
  assign n121_I_t1b = n120_O_t1b; // @[Top.scala 41:12]
  assign n122_valid_up = n121_valid_down; // @[Top.scala 46:19]
  assign n122_I0 = n121_O; // @[Top.scala 44:13]
  assign n122_I1 = 8'h1; // @[Top.scala 45:13]
  assign n123_valid_up = n122_valid_down; // @[Top.scala 49:19]
  assign n123_I_t0b = n122_O_t0b; // @[Top.scala 48:12]
  assign n123_I_t1b = n122_O_t1b; // @[Top.scala 48:12]
  assign n124_valid_up = n123_valid_down; // @[Top.scala 53:19]
  assign n124_I0 = I; // @[Top.scala 51:13]
  assign n124_I1 = n123_O; // @[Top.scala 52:13]
  assign n125_valid_up = n124_valid_down; // @[Top.scala 56:19]
  assign n125_I_t0b = n124_O_t0b; // @[Top.scala 55:12]
  assign n125_I_t1b = n124_O_t1b; // @[Top.scala 55:12]
  assign n126_valid_up = n125_valid_down; // @[Top.scala 59:19]
  assign n126_I = n125_O[0]; // @[Top.scala 58:12]
endmodule
module MapS_5(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7,
  output        O_8,
  output        O_9,
  output        O_10,
  output        O_11,
  output        O_12,
  output        O_13,
  output        O_14,
  output        O_15
);
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire  other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire  other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_2_I; // @[MapS.scala 10:86]
  wire  other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_3_I; // @[MapS.scala 10:86]
  wire  other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_4_I; // @[MapS.scala 10:86]
  wire  other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_5_I; // @[MapS.scala 10:86]
  wire  other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_6_I; // @[MapS.scala 10:86]
  wire  other_ops_6_O; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_7_I; // @[MapS.scala 10:86]
  wire  other_ops_7_O; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_8_I; // @[MapS.scala 10:86]
  wire  other_ops_8_O; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_9_I; // @[MapS.scala 10:86]
  wire  other_ops_9_O; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_10_I; // @[MapS.scala 10:86]
  wire  other_ops_10_O; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_11_I; // @[MapS.scala 10:86]
  wire  other_ops_11_O; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_12_I; // @[MapS.scala 10:86]
  wire  other_ops_12_O; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_13_I; // @[MapS.scala 10:86]
  wire  other_ops_13_O; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [31:0] other_ops_14_I; // @[MapS.scala 10:86]
  wire  other_ops_14_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_1 fst_op ( // @[MapS.scala 9:22]
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  Module_1 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  Module_1 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  Module_1 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_2_valid_down),
    .I(other_ops_2_I),
    .O(other_ops_2_O)
  );
  Module_1 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_3_valid_down),
    .I(other_ops_3_I),
    .O(other_ops_3_O)
  );
  Module_1 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_4_valid_down),
    .I(other_ops_4_I),
    .O(other_ops_4_O)
  );
  Module_1 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_5_valid_down),
    .I(other_ops_5_I),
    .O(other_ops_5_O)
  );
  Module_1 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_6_valid_down),
    .I(other_ops_6_I),
    .O(other_ops_6_O)
  );
  Module_1 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_7_valid_down),
    .I(other_ops_7_I),
    .O(other_ops_7_O)
  );
  Module_1 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_8_valid_down),
    .I(other_ops_8_I),
    .O(other_ops_8_O)
  );
  Module_1 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_9_valid_down),
    .I(other_ops_9_I),
    .O(other_ops_9_O)
  );
  Module_1 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_10_valid_down),
    .I(other_ops_10_I),
    .O(other_ops_10_O)
  );
  Module_1 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_11_valid_down),
    .I(other_ops_11_I),
    .O(other_ops_11_O)
  );
  Module_1 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_12_valid_down),
    .I(other_ops_12_I),
    .O(other_ops_12_O)
  );
  Module_1 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_13_valid_down),
    .I(other_ops_13_I),
    .O(other_ops_13_O)
  );
  Module_1 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_down(other_ops_14_valid_down),
    .I(other_ops_14_I),
    .O(other_ops_14_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign O_8 = other_ops_7_O; // @[MapS.scala 21:12]
  assign O_9 = other_ops_8_O; // @[MapS.scala 21:12]
  assign O_10 = other_ops_9_O; // @[MapS.scala 21:12]
  assign O_11 = other_ops_10_O; // @[MapS.scala 21:12]
  assign O_12 = other_ops_11_O; // @[MapS.scala 21:12]
  assign O_13 = other_ops_12_O; // @[MapS.scala 21:12]
  assign O_14 = other_ops_13_O; // @[MapS.scala 21:12]
  assign O_15 = other_ops_14_O; // @[MapS.scala 21:12]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
  assign other_ops_2_I = I_3; // @[MapS.scala 20:41]
  assign other_ops_3_I = I_4; // @[MapS.scala 20:41]
  assign other_ops_4_I = I_5; // @[MapS.scala 20:41]
  assign other_ops_5_I = I_6; // @[MapS.scala 20:41]
  assign other_ops_6_I = I_7; // @[MapS.scala 20:41]
  assign other_ops_7_I = I_8; // @[MapS.scala 20:41]
  assign other_ops_8_I = I_9; // @[MapS.scala 20:41]
  assign other_ops_9_I = I_10; // @[MapS.scala 20:41]
  assign other_ops_10_I = I_11; // @[MapS.scala 20:41]
  assign other_ops_11_I = I_12; // @[MapS.scala 20:41]
  assign other_ops_12_I = I_13; // @[MapS.scala 20:41]
  assign other_ops_13_I = I_14; // @[MapS.scala 20:41]
  assign other_ops_14_I = I_15; // @[MapS.scala 20:41]
endmodule
module MapT_9(
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output        O_0,
  output        O_1,
  output        O_2,
  output        O_3,
  output        O_4,
  output        O_5,
  output        O_6,
  output        O_7,
  output        O_8,
  output        O_9,
  output        O_10,
  output        O_11,
  output        O_12,
  output        O_13,
  output        O_14,
  output        O_15
);
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3; // @[MapT.scala 8:20]
  wire [31:0] op_I_4; // @[MapT.scala 8:20]
  wire [31:0] op_I_5; // @[MapT.scala 8:20]
  wire [31:0] op_I_6; // @[MapT.scala 8:20]
  wire [31:0] op_I_7; // @[MapT.scala 8:20]
  wire [31:0] op_I_8; // @[MapT.scala 8:20]
  wire [31:0] op_I_9; // @[MapT.scala 8:20]
  wire [31:0] op_I_10; // @[MapT.scala 8:20]
  wire [31:0] op_I_11; // @[MapT.scala 8:20]
  wire [31:0] op_I_12; // @[MapT.scala 8:20]
  wire [31:0] op_I_13; // @[MapT.scala 8:20]
  wire [31:0] op_I_14; // @[MapT.scala 8:20]
  wire [31:0] op_I_15; // @[MapT.scala 8:20]
  wire  op_O_0; // @[MapT.scala 8:20]
  wire  op_O_1; // @[MapT.scala 8:20]
  wire  op_O_2; // @[MapT.scala 8:20]
  wire  op_O_3; // @[MapT.scala 8:20]
  wire  op_O_4; // @[MapT.scala 8:20]
  wire  op_O_5; // @[MapT.scala 8:20]
  wire  op_O_6; // @[MapT.scala 8:20]
  wire  op_O_7; // @[MapT.scala 8:20]
  wire  op_O_8; // @[MapT.scala 8:20]
  wire  op_O_9; // @[MapT.scala 8:20]
  wire  op_O_10; // @[MapT.scala 8:20]
  wire  op_O_11; // @[MapT.scala 8:20]
  wire  op_O_12; // @[MapT.scala 8:20]
  wire  op_O_13; // @[MapT.scala 8:20]
  wire  op_O_14; // @[MapT.scala 8:20]
  wire  op_O_15; // @[MapT.scala 8:20]
  MapS_5 op ( // @[MapT.scala 8:20]
    .valid_down(op_valid_down),
    .I_0(op_I_0),
    .I_1(op_I_1),
    .I_2(op_I_2),
    .I_3(op_I_3),
    .I_4(op_I_4),
    .I_5(op_I_5),
    .I_6(op_I_6),
    .I_7(op_I_7),
    .I_8(op_I_8),
    .I_9(op_I_9),
    .I_10(op_I_10),
    .I_11(op_I_11),
    .I_12(op_I_12),
    .I_13(op_I_13),
    .I_14(op_I_14),
    .I_15(op_I_15),
    .O_0(op_O_0),
    .O_1(op_O_1),
    .O_2(op_O_2),
    .O_3(op_O_3),
    .O_4(op_O_4),
    .O_5(op_O_5),
    .O_6(op_O_6),
    .O_7(op_O_7),
    .O_8(op_O_8),
    .O_9(op_O_9),
    .O_10(op_O_10),
    .O_11(op_O_11),
    .O_12(op_O_12),
    .O_13(op_O_13),
    .O_14(op_O_14),
    .O_15(op_O_15)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0 = op_O_0; // @[MapT.scala 15:7]
  assign O_1 = op_O_1; // @[MapT.scala 15:7]
  assign O_2 = op_O_2; // @[MapT.scala 15:7]
  assign O_3 = op_O_3; // @[MapT.scala 15:7]
  assign O_4 = op_O_4; // @[MapT.scala 15:7]
  assign O_5 = op_O_5; // @[MapT.scala 15:7]
  assign O_6 = op_O_6; // @[MapT.scala 15:7]
  assign O_7 = op_O_7; // @[MapT.scala 15:7]
  assign O_8 = op_O_8; // @[MapT.scala 15:7]
  assign O_9 = op_O_9; // @[MapT.scala 15:7]
  assign O_10 = op_O_10; // @[MapT.scala 15:7]
  assign O_11 = op_O_11; // @[MapT.scala 15:7]
  assign O_12 = op_O_12; // @[MapT.scala 15:7]
  assign O_13 = op_O_13; // @[MapT.scala 15:7]
  assign O_14 = op_O_14; // @[MapT.scala 15:7]
  assign O_15 = op_O_15; // @[MapT.scala 15:7]
  assign op_I_0 = I_0; // @[MapT.scala 14:10]
  assign op_I_1 = I_1; // @[MapT.scala 14:10]
  assign op_I_2 = I_2; // @[MapT.scala 14:10]
  assign op_I_3 = I_3; // @[MapT.scala 14:10]
  assign op_I_4 = I_4; // @[MapT.scala 14:10]
  assign op_I_5 = I_5; // @[MapT.scala 14:10]
  assign op_I_6 = I_6; // @[MapT.scala 14:10]
  assign op_I_7 = I_7; // @[MapT.scala 14:10]
  assign op_I_8 = I_8; // @[MapT.scala 14:10]
  assign op_I_9 = I_9; // @[MapT.scala 14:10]
  assign op_I_10 = I_10; // @[MapT.scala 14:10]
  assign op_I_11 = I_11; // @[MapT.scala 14:10]
  assign op_I_12 = I_12; // @[MapT.scala 14:10]
  assign op_I_13 = I_13; // @[MapT.scala 14:10]
  assign op_I_14 = I_14; // @[MapT.scala 14:10]
  assign op_I_15 = I_15; // @[MapT.scala 14:10]
endmodule
module AtomTuple_4(
  input   valid_up,
  output  valid_down,
  input   I0,
  input   I1,
  output  O_t0b,
  output  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input   valid_up,
  output  valid_down,
  input   I0_0,
  input   I0_1,
  input   I0_2,
  input   I0_3,
  input   I0_4,
  input   I0_5,
  input   I0_6,
  input   I0_7,
  input   I0_8,
  input   I0_9,
  input   I0_10,
  input   I0_11,
  input   I0_12,
  input   I0_13,
  input   I0_14,
  input   I0_15,
  input   I1_0,
  input   I1_1,
  input   I1_2,
  input   I1_3,
  input   I1_4,
  input   I1_5,
  input   I1_6,
  input   I1_7,
  input   I1_8,
  input   I1_9,
  input   I1_10,
  input   I1_11,
  input   I1_12,
  input   I1_13,
  input   I1_14,
  input   I1_15,
  output  O_0_t0b,
  output  O_0_t1b,
  output  O_1_t0b,
  output  O_1_t1b,
  output  O_2_t0b,
  output  O_2_t1b,
  output  O_3_t0b,
  output  O_3_t1b,
  output  O_4_t0b,
  output  O_4_t1b,
  output  O_5_t0b,
  output  O_5_t1b,
  output  O_6_t0b,
  output  O_6_t1b,
  output  O_7_t0b,
  output  O_7_t1b,
  output  O_8_t0b,
  output  O_8_t1b,
  output  O_9_t0b,
  output  O_9_t1b,
  output  O_10_t0b,
  output  O_10_t1b,
  output  O_11_t0b,
  output  O_11_t1b,
  output  O_12_t0b,
  output  O_12_t1b,
  output  O_13_t0b,
  output  O_13_t1b,
  output  O_14_t0b,
  output  O_14_t1b,
  output  O_15_t0b,
  output  O_15_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire  fst_op_I0; // @[Map2S.scala 9:22]
  wire  fst_op_I1; // @[Map2S.scala 9:22]
  wire  fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire  fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_0_I0; // @[Map2S.scala 10:86]
  wire  other_ops_0_I1; // @[Map2S.scala 10:86]
  wire  other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_1_I0; // @[Map2S.scala 10:86]
  wire  other_ops_1_I1; // @[Map2S.scala 10:86]
  wire  other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_2_I0; // @[Map2S.scala 10:86]
  wire  other_ops_2_I1; // @[Map2S.scala 10:86]
  wire  other_ops_2_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_2_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_3_I0; // @[Map2S.scala 10:86]
  wire  other_ops_3_I1; // @[Map2S.scala 10:86]
  wire  other_ops_3_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_3_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_4_I0; // @[Map2S.scala 10:86]
  wire  other_ops_4_I1; // @[Map2S.scala 10:86]
  wire  other_ops_4_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_4_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_5_I0; // @[Map2S.scala 10:86]
  wire  other_ops_5_I1; // @[Map2S.scala 10:86]
  wire  other_ops_5_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_5_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_6_I0; // @[Map2S.scala 10:86]
  wire  other_ops_6_I1; // @[Map2S.scala 10:86]
  wire  other_ops_6_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_6_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_7_I0; // @[Map2S.scala 10:86]
  wire  other_ops_7_I1; // @[Map2S.scala 10:86]
  wire  other_ops_7_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_7_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_8_I0; // @[Map2S.scala 10:86]
  wire  other_ops_8_I1; // @[Map2S.scala 10:86]
  wire  other_ops_8_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_8_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_9_I0; // @[Map2S.scala 10:86]
  wire  other_ops_9_I1; // @[Map2S.scala 10:86]
  wire  other_ops_9_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_9_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_10_I0; // @[Map2S.scala 10:86]
  wire  other_ops_10_I1; // @[Map2S.scala 10:86]
  wire  other_ops_10_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_10_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_11_I0; // @[Map2S.scala 10:86]
  wire  other_ops_11_I1; // @[Map2S.scala 10:86]
  wire  other_ops_11_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_11_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_12_I0; // @[Map2S.scala 10:86]
  wire  other_ops_12_I1; // @[Map2S.scala 10:86]
  wire  other_ops_12_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_12_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_13_I0; // @[Map2S.scala 10:86]
  wire  other_ops_13_I1; // @[Map2S.scala 10:86]
  wire  other_ops_13_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_13_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire  other_ops_14_I0; // @[Map2S.scala 10:86]
  wire  other_ops_14_I1; // @[Map2S.scala 10:86]
  wire  other_ops_14_O_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_14_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  AtomTuple_4 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple_4 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple_4 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  AtomTuple_4 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_t0b(other_ops_2_O_t0b),
    .O_t1b(other_ops_2_O_t1b)
  );
  AtomTuple_4 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_t0b(other_ops_3_O_t0b),
    .O_t1b(other_ops_3_O_t1b)
  );
  AtomTuple_4 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_t0b(other_ops_4_O_t0b),
    .O_t1b(other_ops_4_O_t1b)
  );
  AtomTuple_4 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_t0b(other_ops_5_O_t0b),
    .O_t1b(other_ops_5_O_t1b)
  );
  AtomTuple_4 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_t0b(other_ops_6_O_t0b),
    .O_t1b(other_ops_6_O_t1b)
  );
  AtomTuple_4 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0(other_ops_7_I0),
    .I1(other_ops_7_I1),
    .O_t0b(other_ops_7_O_t0b),
    .O_t1b(other_ops_7_O_t1b)
  );
  AtomTuple_4 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0(other_ops_8_I0),
    .I1(other_ops_8_I1),
    .O_t0b(other_ops_8_O_t0b),
    .O_t1b(other_ops_8_O_t1b)
  );
  AtomTuple_4 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0(other_ops_9_I0),
    .I1(other_ops_9_I1),
    .O_t0b(other_ops_9_O_t0b),
    .O_t1b(other_ops_9_O_t1b)
  );
  AtomTuple_4 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0(other_ops_10_I0),
    .I1(other_ops_10_I1),
    .O_t0b(other_ops_10_O_t0b),
    .O_t1b(other_ops_10_O_t1b)
  );
  AtomTuple_4 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0(other_ops_11_I0),
    .I1(other_ops_11_I1),
    .O_t0b(other_ops_11_O_t0b),
    .O_t1b(other_ops_11_O_t1b)
  );
  AtomTuple_4 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0(other_ops_12_I0),
    .I1(other_ops_12_I1),
    .O_t0b(other_ops_12_O_t0b),
    .O_t1b(other_ops_12_O_t1b)
  );
  AtomTuple_4 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0(other_ops_13_I0),
    .I1(other_ops_13_I1),
    .O_t0b(other_ops_13_O_t0b),
    .O_t1b(other_ops_13_O_t1b)
  );
  AtomTuple_4 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0(other_ops_14_I0),
    .I1(other_ops_14_I1),
    .O_t0b(other_ops_14_O_t0b),
    .O_t1b(other_ops_14_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign O_3_t0b = other_ops_2_O_t0b; // @[Map2S.scala 24:12]
  assign O_3_t1b = other_ops_2_O_t1b; // @[Map2S.scala 24:12]
  assign O_4_t0b = other_ops_3_O_t0b; // @[Map2S.scala 24:12]
  assign O_4_t1b = other_ops_3_O_t1b; // @[Map2S.scala 24:12]
  assign O_5_t0b = other_ops_4_O_t0b; // @[Map2S.scala 24:12]
  assign O_5_t1b = other_ops_4_O_t1b; // @[Map2S.scala 24:12]
  assign O_6_t0b = other_ops_5_O_t0b; // @[Map2S.scala 24:12]
  assign O_6_t1b = other_ops_5_O_t1b; // @[Map2S.scala 24:12]
  assign O_7_t0b = other_ops_6_O_t0b; // @[Map2S.scala 24:12]
  assign O_7_t1b = other_ops_6_O_t1b; // @[Map2S.scala 24:12]
  assign O_8_t0b = other_ops_7_O_t0b; // @[Map2S.scala 24:12]
  assign O_8_t1b = other_ops_7_O_t1b; // @[Map2S.scala 24:12]
  assign O_9_t0b = other_ops_8_O_t0b; // @[Map2S.scala 24:12]
  assign O_9_t1b = other_ops_8_O_t1b; // @[Map2S.scala 24:12]
  assign O_10_t0b = other_ops_9_O_t0b; // @[Map2S.scala 24:12]
  assign O_10_t1b = other_ops_9_O_t1b; // @[Map2S.scala 24:12]
  assign O_11_t0b = other_ops_10_O_t0b; // @[Map2S.scala 24:12]
  assign O_11_t1b = other_ops_10_O_t1b; // @[Map2S.scala 24:12]
  assign O_12_t0b = other_ops_11_O_t0b; // @[Map2S.scala 24:12]
  assign O_12_t1b = other_ops_11_O_t1b; // @[Map2S.scala 24:12]
  assign O_13_t0b = other_ops_12_O_t0b; // @[Map2S.scala 24:12]
  assign O_13_t1b = other_ops_12_O_t1b; // @[Map2S.scala 24:12]
  assign O_14_t0b = other_ops_13_O_t0b; // @[Map2S.scala 24:12]
  assign O_14_t1b = other_ops_13_O_t1b; // @[Map2S.scala 24:12]
  assign O_15_t0b = other_ops_14_O_t0b; // @[Map2S.scala 24:12]
  assign O_15_t1b = other_ops_14_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0 = I0_8; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0 = I0_9; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0 = I0_10; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0 = I0_11; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0 = I0_12; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0 = I0_13; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0 = I0_14; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0 = I0_15; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T_8(
  input   valid_up,
  output  valid_down,
  input   I0_0,
  input   I0_1,
  input   I0_2,
  input   I0_3,
  input   I0_4,
  input   I0_5,
  input   I0_6,
  input   I0_7,
  input   I0_8,
  input   I0_9,
  input   I0_10,
  input   I0_11,
  input   I0_12,
  input   I0_13,
  input   I0_14,
  input   I0_15,
  input   I1_0,
  input   I1_1,
  input   I1_2,
  input   I1_3,
  input   I1_4,
  input   I1_5,
  input   I1_6,
  input   I1_7,
  input   I1_8,
  input   I1_9,
  input   I1_10,
  input   I1_11,
  input   I1_12,
  input   I1_13,
  input   I1_14,
  input   I1_15,
  output  O_0_t0b,
  output  O_0_t1b,
  output  O_1_t0b,
  output  O_1_t1b,
  output  O_2_t0b,
  output  O_2_t1b,
  output  O_3_t0b,
  output  O_3_t1b,
  output  O_4_t0b,
  output  O_4_t1b,
  output  O_5_t0b,
  output  O_5_t1b,
  output  O_6_t0b,
  output  O_6_t1b,
  output  O_7_t0b,
  output  O_7_t1b,
  output  O_8_t0b,
  output  O_8_t1b,
  output  O_9_t0b,
  output  O_9_t1b,
  output  O_10_t0b,
  output  O_10_t1b,
  output  O_11_t0b,
  output  O_11_t1b,
  output  O_12_t0b,
  output  O_12_t1b,
  output  O_13_t0b,
  output  O_13_t1b,
  output  O_14_t0b,
  output  O_14_t1b,
  output  O_15_t0b,
  output  O_15_t1b
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire  op_I0_0; // @[Map2T.scala 8:20]
  wire  op_I0_1; // @[Map2T.scala 8:20]
  wire  op_I0_2; // @[Map2T.scala 8:20]
  wire  op_I0_3; // @[Map2T.scala 8:20]
  wire  op_I0_4; // @[Map2T.scala 8:20]
  wire  op_I0_5; // @[Map2T.scala 8:20]
  wire  op_I0_6; // @[Map2T.scala 8:20]
  wire  op_I0_7; // @[Map2T.scala 8:20]
  wire  op_I0_8; // @[Map2T.scala 8:20]
  wire  op_I0_9; // @[Map2T.scala 8:20]
  wire  op_I0_10; // @[Map2T.scala 8:20]
  wire  op_I0_11; // @[Map2T.scala 8:20]
  wire  op_I0_12; // @[Map2T.scala 8:20]
  wire  op_I0_13; // @[Map2T.scala 8:20]
  wire  op_I0_14; // @[Map2T.scala 8:20]
  wire  op_I0_15; // @[Map2T.scala 8:20]
  wire  op_I1_0; // @[Map2T.scala 8:20]
  wire  op_I1_1; // @[Map2T.scala 8:20]
  wire  op_I1_2; // @[Map2T.scala 8:20]
  wire  op_I1_3; // @[Map2T.scala 8:20]
  wire  op_I1_4; // @[Map2T.scala 8:20]
  wire  op_I1_5; // @[Map2T.scala 8:20]
  wire  op_I1_6; // @[Map2T.scala 8:20]
  wire  op_I1_7; // @[Map2T.scala 8:20]
  wire  op_I1_8; // @[Map2T.scala 8:20]
  wire  op_I1_9; // @[Map2T.scala 8:20]
  wire  op_I1_10; // @[Map2T.scala 8:20]
  wire  op_I1_11; // @[Map2T.scala 8:20]
  wire  op_I1_12; // @[Map2T.scala 8:20]
  wire  op_I1_13; // @[Map2T.scala 8:20]
  wire  op_I1_14; // @[Map2T.scala 8:20]
  wire  op_I1_15; // @[Map2T.scala 8:20]
  wire  op_O_0_t0b; // @[Map2T.scala 8:20]
  wire  op_O_0_t1b; // @[Map2T.scala 8:20]
  wire  op_O_1_t0b; // @[Map2T.scala 8:20]
  wire  op_O_1_t1b; // @[Map2T.scala 8:20]
  wire  op_O_2_t0b; // @[Map2T.scala 8:20]
  wire  op_O_2_t1b; // @[Map2T.scala 8:20]
  wire  op_O_3_t0b; // @[Map2T.scala 8:20]
  wire  op_O_3_t1b; // @[Map2T.scala 8:20]
  wire  op_O_4_t0b; // @[Map2T.scala 8:20]
  wire  op_O_4_t1b; // @[Map2T.scala 8:20]
  wire  op_O_5_t0b; // @[Map2T.scala 8:20]
  wire  op_O_5_t1b; // @[Map2T.scala 8:20]
  wire  op_O_6_t0b; // @[Map2T.scala 8:20]
  wire  op_O_6_t1b; // @[Map2T.scala 8:20]
  wire  op_O_7_t0b; // @[Map2T.scala 8:20]
  wire  op_O_7_t1b; // @[Map2T.scala 8:20]
  wire  op_O_8_t0b; // @[Map2T.scala 8:20]
  wire  op_O_8_t1b; // @[Map2T.scala 8:20]
  wire  op_O_9_t0b; // @[Map2T.scala 8:20]
  wire  op_O_9_t1b; // @[Map2T.scala 8:20]
  wire  op_O_10_t0b; // @[Map2T.scala 8:20]
  wire  op_O_10_t1b; // @[Map2T.scala 8:20]
  wire  op_O_11_t0b; // @[Map2T.scala 8:20]
  wire  op_O_11_t1b; // @[Map2T.scala 8:20]
  wire  op_O_12_t0b; // @[Map2T.scala 8:20]
  wire  op_O_12_t1b; // @[Map2T.scala 8:20]
  wire  op_O_13_t0b; // @[Map2T.scala 8:20]
  wire  op_O_13_t1b; // @[Map2T.scala 8:20]
  wire  op_O_14_t0b; // @[Map2T.scala 8:20]
  wire  op_O_14_t1b; // @[Map2T.scala 8:20]
  wire  op_O_15_t0b; // @[Map2T.scala 8:20]
  wire  op_O_15_t1b; // @[Map2T.scala 8:20]
  Map2S_8 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I0_8(op_I0_8),
    .I0_9(op_I0_9),
    .I0_10(op_I0_10),
    .I0_11(op_I0_11),
    .I0_12(op_I0_12),
    .I0_13(op_I0_13),
    .I0_14(op_I0_14),
    .I0_15(op_I0_15),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_t0b(op_O_0_t0b),
    .O_0_t1b(op_O_0_t1b),
    .O_1_t0b(op_O_1_t0b),
    .O_1_t1b(op_O_1_t1b),
    .O_2_t0b(op_O_2_t0b),
    .O_2_t1b(op_O_2_t1b),
    .O_3_t0b(op_O_3_t0b),
    .O_3_t1b(op_O_3_t1b),
    .O_4_t0b(op_O_4_t0b),
    .O_4_t1b(op_O_4_t1b),
    .O_5_t0b(op_O_5_t0b),
    .O_5_t1b(op_O_5_t1b),
    .O_6_t0b(op_O_6_t0b),
    .O_6_t1b(op_O_6_t1b),
    .O_7_t0b(op_O_7_t0b),
    .O_7_t1b(op_O_7_t1b),
    .O_8_t0b(op_O_8_t0b),
    .O_8_t1b(op_O_8_t1b),
    .O_9_t0b(op_O_9_t0b),
    .O_9_t1b(op_O_9_t1b),
    .O_10_t0b(op_O_10_t0b),
    .O_10_t1b(op_O_10_t1b),
    .O_11_t0b(op_O_11_t0b),
    .O_11_t1b(op_O_11_t1b),
    .O_12_t0b(op_O_12_t0b),
    .O_12_t1b(op_O_12_t1b),
    .O_13_t0b(op_O_13_t0b),
    .O_13_t1b(op_O_13_t1b),
    .O_14_t0b(op_O_14_t0b),
    .O_14_t1b(op_O_14_t1b),
    .O_15_t0b(op_O_15_t0b),
    .O_15_t1b(op_O_15_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_t0b = op_O_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_t1b = op_O_0_t1b; // @[Map2T.scala 17:7]
  assign O_1_t0b = op_O_1_t0b; // @[Map2T.scala 17:7]
  assign O_1_t1b = op_O_1_t1b; // @[Map2T.scala 17:7]
  assign O_2_t0b = op_O_2_t0b; // @[Map2T.scala 17:7]
  assign O_2_t1b = op_O_2_t1b; // @[Map2T.scala 17:7]
  assign O_3_t0b = op_O_3_t0b; // @[Map2T.scala 17:7]
  assign O_3_t1b = op_O_3_t1b; // @[Map2T.scala 17:7]
  assign O_4_t0b = op_O_4_t0b; // @[Map2T.scala 17:7]
  assign O_4_t1b = op_O_4_t1b; // @[Map2T.scala 17:7]
  assign O_5_t0b = op_O_5_t0b; // @[Map2T.scala 17:7]
  assign O_5_t1b = op_O_5_t1b; // @[Map2T.scala 17:7]
  assign O_6_t0b = op_O_6_t0b; // @[Map2T.scala 17:7]
  assign O_6_t1b = op_O_6_t1b; // @[Map2T.scala 17:7]
  assign O_7_t0b = op_O_7_t0b; // @[Map2T.scala 17:7]
  assign O_7_t1b = op_O_7_t1b; // @[Map2T.scala 17:7]
  assign O_8_t0b = op_O_8_t0b; // @[Map2T.scala 17:7]
  assign O_8_t1b = op_O_8_t1b; // @[Map2T.scala 17:7]
  assign O_9_t0b = op_O_9_t0b; // @[Map2T.scala 17:7]
  assign O_9_t1b = op_O_9_t1b; // @[Map2T.scala 17:7]
  assign O_10_t0b = op_O_10_t0b; // @[Map2T.scala 17:7]
  assign O_10_t1b = op_O_10_t1b; // @[Map2T.scala 17:7]
  assign O_11_t0b = op_O_11_t0b; // @[Map2T.scala 17:7]
  assign O_11_t1b = op_O_11_t1b; // @[Map2T.scala 17:7]
  assign O_12_t0b = op_O_12_t0b; // @[Map2T.scala 17:7]
  assign O_12_t1b = op_O_12_t1b; // @[Map2T.scala 17:7]
  assign O_13_t0b = op_O_13_t0b; // @[Map2T.scala 17:7]
  assign O_13_t1b = op_O_13_t1b; // @[Map2T.scala 17:7]
  assign O_14_t0b = op_O_14_t0b; // @[Map2T.scala 17:7]
  assign O_14_t1b = op_O_14_t1b; // @[Map2T.scala 17:7]
  assign O_15_t0b = op_O_15_t0b; // @[Map2T.scala 17:7]
  assign O_15_t1b = op_O_15_t1b; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I0_8 = I0_8; // @[Map2T.scala 15:11]
  assign op_I0_9 = I0_9; // @[Map2T.scala 15:11]
  assign op_I0_10 = I0_10; // @[Map2T.scala 15:11]
  assign op_I0_11 = I0_11; // @[Map2T.scala 15:11]
  assign op_I0_12 = I0_12; // @[Map2T.scala 15:11]
  assign op_I0_13 = I0_13; // @[Map2T.scala 15:11]
  assign op_I0_14 = I0_14; // @[Map2T.scala 15:11]
  assign op_I0_15 = I0_15; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module PartitionS_4(
  input   valid_up,
  output  valid_down,
  input   I_0_t0b,
  input   I_0_t1b,
  input   I_1_t0b,
  input   I_1_t1b,
  input   I_2_t0b,
  input   I_2_t1b,
  input   I_3_t0b,
  input   I_3_t1b,
  input   I_4_t0b,
  input   I_4_t1b,
  input   I_5_t0b,
  input   I_5_t1b,
  input   I_6_t0b,
  input   I_6_t1b,
  input   I_7_t0b,
  input   I_7_t1b,
  input   I_8_t0b,
  input   I_8_t1b,
  input   I_9_t0b,
  input   I_9_t1b,
  input   I_10_t0b,
  input   I_10_t1b,
  input   I_11_t0b,
  input   I_11_t1b,
  input   I_12_t0b,
  input   I_12_t1b,
  input   I_13_t0b,
  input   I_13_t1b,
  input   I_14_t0b,
  input   I_14_t1b,
  input   I_15_t0b,
  input   I_15_t1b,
  output  O_0_0_t0b,
  output  O_0_0_t1b,
  output  O_1_0_t0b,
  output  O_1_0_t1b,
  output  O_2_0_t0b,
  output  O_2_0_t1b,
  output  O_3_0_t0b,
  output  O_3_0_t1b,
  output  O_4_0_t0b,
  output  O_4_0_t1b,
  output  O_5_0_t0b,
  output  O_5_0_t1b,
  output  O_6_0_t0b,
  output  O_6_0_t1b,
  output  O_7_0_t0b,
  output  O_7_0_t1b,
  output  O_8_0_t0b,
  output  O_8_0_t1b,
  output  O_9_0_t0b,
  output  O_9_0_t1b,
  output  O_10_0_t0b,
  output  O_10_0_t1b,
  output  O_11_0_t0b,
  output  O_11_0_t1b,
  output  O_12_0_t0b,
  output  O_12_0_t1b,
  output  O_13_0_t0b,
  output  O_13_0_t1b,
  output  O_14_0_t0b,
  output  O_14_0_t1b,
  output  O_15_0_t0b,
  output  O_15_0_t1b
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_t0b = I_0_t0b; // @[Partition.scala 15:39]
  assign O_0_0_t1b = I_0_t1b; // @[Partition.scala 15:39]
  assign O_1_0_t0b = I_1_t0b; // @[Partition.scala 15:39]
  assign O_1_0_t1b = I_1_t1b; // @[Partition.scala 15:39]
  assign O_2_0_t0b = I_2_t0b; // @[Partition.scala 15:39]
  assign O_2_0_t1b = I_2_t1b; // @[Partition.scala 15:39]
  assign O_3_0_t0b = I_3_t0b; // @[Partition.scala 15:39]
  assign O_3_0_t1b = I_3_t1b; // @[Partition.scala 15:39]
  assign O_4_0_t0b = I_4_t0b; // @[Partition.scala 15:39]
  assign O_4_0_t1b = I_4_t1b; // @[Partition.scala 15:39]
  assign O_5_0_t0b = I_5_t0b; // @[Partition.scala 15:39]
  assign O_5_0_t1b = I_5_t1b; // @[Partition.scala 15:39]
  assign O_6_0_t0b = I_6_t0b; // @[Partition.scala 15:39]
  assign O_6_0_t1b = I_6_t1b; // @[Partition.scala 15:39]
  assign O_7_0_t0b = I_7_t0b; // @[Partition.scala 15:39]
  assign O_7_0_t1b = I_7_t1b; // @[Partition.scala 15:39]
  assign O_8_0_t0b = I_8_t0b; // @[Partition.scala 15:39]
  assign O_8_0_t1b = I_8_t1b; // @[Partition.scala 15:39]
  assign O_9_0_t0b = I_9_t0b; // @[Partition.scala 15:39]
  assign O_9_0_t1b = I_9_t1b; // @[Partition.scala 15:39]
  assign O_10_0_t0b = I_10_t0b; // @[Partition.scala 15:39]
  assign O_10_0_t1b = I_10_t1b; // @[Partition.scala 15:39]
  assign O_11_0_t0b = I_11_t0b; // @[Partition.scala 15:39]
  assign O_11_0_t1b = I_11_t1b; // @[Partition.scala 15:39]
  assign O_12_0_t0b = I_12_t0b; // @[Partition.scala 15:39]
  assign O_12_0_t1b = I_12_t1b; // @[Partition.scala 15:39]
  assign O_13_0_t0b = I_13_t0b; // @[Partition.scala 15:39]
  assign O_13_0_t1b = I_13_t1b; // @[Partition.scala 15:39]
  assign O_14_0_t0b = I_14_t0b; // @[Partition.scala 15:39]
  assign O_14_0_t1b = I_14_t1b; // @[Partition.scala 15:39]
  assign O_15_0_t0b = I_15_t0b; // @[Partition.scala 15:39]
  assign O_15_0_t1b = I_15_t1b; // @[Partition.scala 15:39]
endmodule
module MapT_10(
  input   valid_up,
  output  valid_down,
  input   I_0_t0b,
  input   I_0_t1b,
  input   I_1_t0b,
  input   I_1_t1b,
  input   I_2_t0b,
  input   I_2_t1b,
  input   I_3_t0b,
  input   I_3_t1b,
  input   I_4_t0b,
  input   I_4_t1b,
  input   I_5_t0b,
  input   I_5_t1b,
  input   I_6_t0b,
  input   I_6_t1b,
  input   I_7_t0b,
  input   I_7_t1b,
  input   I_8_t0b,
  input   I_8_t1b,
  input   I_9_t0b,
  input   I_9_t1b,
  input   I_10_t0b,
  input   I_10_t1b,
  input   I_11_t0b,
  input   I_11_t1b,
  input   I_12_t0b,
  input   I_12_t1b,
  input   I_13_t0b,
  input   I_13_t1b,
  input   I_14_t0b,
  input   I_14_t1b,
  input   I_15_t0b,
  input   I_15_t1b,
  output  O_0_0_t0b,
  output  O_0_0_t1b,
  output  O_1_0_t0b,
  output  O_1_0_t1b,
  output  O_2_0_t0b,
  output  O_2_0_t1b,
  output  O_3_0_t0b,
  output  O_3_0_t1b,
  output  O_4_0_t0b,
  output  O_4_0_t1b,
  output  O_5_0_t0b,
  output  O_5_0_t1b,
  output  O_6_0_t0b,
  output  O_6_0_t1b,
  output  O_7_0_t0b,
  output  O_7_0_t1b,
  output  O_8_0_t0b,
  output  O_8_0_t1b,
  output  O_9_0_t0b,
  output  O_9_0_t1b,
  output  O_10_0_t0b,
  output  O_10_0_t1b,
  output  O_11_0_t0b,
  output  O_11_0_t1b,
  output  O_12_0_t0b,
  output  O_12_0_t1b,
  output  O_13_0_t0b,
  output  O_13_0_t1b,
  output  O_14_0_t0b,
  output  O_14_0_t1b,
  output  O_15_0_t0b,
  output  O_15_0_t1b
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire  op_I_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_1_t0b; // @[MapT.scala 8:20]
  wire  op_I_1_t1b; // @[MapT.scala 8:20]
  wire  op_I_2_t0b; // @[MapT.scala 8:20]
  wire  op_I_2_t1b; // @[MapT.scala 8:20]
  wire  op_I_3_t0b; // @[MapT.scala 8:20]
  wire  op_I_3_t1b; // @[MapT.scala 8:20]
  wire  op_I_4_t0b; // @[MapT.scala 8:20]
  wire  op_I_4_t1b; // @[MapT.scala 8:20]
  wire  op_I_5_t0b; // @[MapT.scala 8:20]
  wire  op_I_5_t1b; // @[MapT.scala 8:20]
  wire  op_I_6_t0b; // @[MapT.scala 8:20]
  wire  op_I_6_t1b; // @[MapT.scala 8:20]
  wire  op_I_7_t0b; // @[MapT.scala 8:20]
  wire  op_I_7_t1b; // @[MapT.scala 8:20]
  wire  op_I_8_t0b; // @[MapT.scala 8:20]
  wire  op_I_8_t1b; // @[MapT.scala 8:20]
  wire  op_I_9_t0b; // @[MapT.scala 8:20]
  wire  op_I_9_t1b; // @[MapT.scala 8:20]
  wire  op_I_10_t0b; // @[MapT.scala 8:20]
  wire  op_I_10_t1b; // @[MapT.scala 8:20]
  wire  op_I_11_t0b; // @[MapT.scala 8:20]
  wire  op_I_11_t1b; // @[MapT.scala 8:20]
  wire  op_I_12_t0b; // @[MapT.scala 8:20]
  wire  op_I_12_t1b; // @[MapT.scala 8:20]
  wire  op_I_13_t0b; // @[MapT.scala 8:20]
  wire  op_I_13_t1b; // @[MapT.scala 8:20]
  wire  op_I_14_t0b; // @[MapT.scala 8:20]
  wire  op_I_14_t1b; // @[MapT.scala 8:20]
  wire  op_I_15_t0b; // @[MapT.scala 8:20]
  wire  op_I_15_t1b; // @[MapT.scala 8:20]
  wire  op_O_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_1_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_1_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_2_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_2_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_3_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_3_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_4_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_4_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_5_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_5_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_6_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_6_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_7_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_7_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_8_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_8_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_9_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_9_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_10_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_10_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_11_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_11_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_12_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_12_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_13_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_13_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_14_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_14_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_15_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_15_0_t1b; // @[MapT.scala 8:20]
  PartitionS_4 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_t0b(op_I_0_t0b),
    .I_0_t1b(op_I_0_t1b),
    .I_1_t0b(op_I_1_t0b),
    .I_1_t1b(op_I_1_t1b),
    .I_2_t0b(op_I_2_t0b),
    .I_2_t1b(op_I_2_t1b),
    .I_3_t0b(op_I_3_t0b),
    .I_3_t1b(op_I_3_t1b),
    .I_4_t0b(op_I_4_t0b),
    .I_4_t1b(op_I_4_t1b),
    .I_5_t0b(op_I_5_t0b),
    .I_5_t1b(op_I_5_t1b),
    .I_6_t0b(op_I_6_t0b),
    .I_6_t1b(op_I_6_t1b),
    .I_7_t0b(op_I_7_t0b),
    .I_7_t1b(op_I_7_t1b),
    .I_8_t0b(op_I_8_t0b),
    .I_8_t1b(op_I_8_t1b),
    .I_9_t0b(op_I_9_t0b),
    .I_9_t1b(op_I_9_t1b),
    .I_10_t0b(op_I_10_t0b),
    .I_10_t1b(op_I_10_t1b),
    .I_11_t0b(op_I_11_t0b),
    .I_11_t1b(op_I_11_t1b),
    .I_12_t0b(op_I_12_t0b),
    .I_12_t1b(op_I_12_t1b),
    .I_13_t0b(op_I_13_t0b),
    .I_13_t1b(op_I_13_t1b),
    .I_14_t0b(op_I_14_t0b),
    .I_14_t1b(op_I_14_t1b),
    .I_15_t0b(op_I_15_t0b),
    .I_15_t1b(op_I_15_t1b),
    .O_0_0_t0b(op_O_0_0_t0b),
    .O_0_0_t1b(op_O_0_0_t1b),
    .O_1_0_t0b(op_O_1_0_t0b),
    .O_1_0_t1b(op_O_1_0_t1b),
    .O_2_0_t0b(op_O_2_0_t0b),
    .O_2_0_t1b(op_O_2_0_t1b),
    .O_3_0_t0b(op_O_3_0_t0b),
    .O_3_0_t1b(op_O_3_0_t1b),
    .O_4_0_t0b(op_O_4_0_t0b),
    .O_4_0_t1b(op_O_4_0_t1b),
    .O_5_0_t0b(op_O_5_0_t0b),
    .O_5_0_t1b(op_O_5_0_t1b),
    .O_6_0_t0b(op_O_6_0_t0b),
    .O_6_0_t1b(op_O_6_0_t1b),
    .O_7_0_t0b(op_O_7_0_t0b),
    .O_7_0_t1b(op_O_7_0_t1b),
    .O_8_0_t0b(op_O_8_0_t0b),
    .O_8_0_t1b(op_O_8_0_t1b),
    .O_9_0_t0b(op_O_9_0_t0b),
    .O_9_0_t1b(op_O_9_0_t1b),
    .O_10_0_t0b(op_O_10_0_t0b),
    .O_10_0_t1b(op_O_10_0_t1b),
    .O_11_0_t0b(op_O_11_0_t0b),
    .O_11_0_t1b(op_O_11_0_t1b),
    .O_12_0_t0b(op_O_12_0_t0b),
    .O_12_0_t1b(op_O_12_0_t1b),
    .O_13_0_t0b(op_O_13_0_t0b),
    .O_13_0_t1b(op_O_13_0_t1b),
    .O_14_0_t0b(op_O_14_0_t0b),
    .O_14_0_t1b(op_O_14_0_t1b),
    .O_15_0_t0b(op_O_15_0_t0b),
    .O_15_0_t1b(op_O_15_0_t1b)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_t0b = op_O_0_0_t0b; // @[MapT.scala 15:7]
  assign O_0_0_t1b = op_O_0_0_t1b; // @[MapT.scala 15:7]
  assign O_1_0_t0b = op_O_1_0_t0b; // @[MapT.scala 15:7]
  assign O_1_0_t1b = op_O_1_0_t1b; // @[MapT.scala 15:7]
  assign O_2_0_t0b = op_O_2_0_t0b; // @[MapT.scala 15:7]
  assign O_2_0_t1b = op_O_2_0_t1b; // @[MapT.scala 15:7]
  assign O_3_0_t0b = op_O_3_0_t0b; // @[MapT.scala 15:7]
  assign O_3_0_t1b = op_O_3_0_t1b; // @[MapT.scala 15:7]
  assign O_4_0_t0b = op_O_4_0_t0b; // @[MapT.scala 15:7]
  assign O_4_0_t1b = op_O_4_0_t1b; // @[MapT.scala 15:7]
  assign O_5_0_t0b = op_O_5_0_t0b; // @[MapT.scala 15:7]
  assign O_5_0_t1b = op_O_5_0_t1b; // @[MapT.scala 15:7]
  assign O_6_0_t0b = op_O_6_0_t0b; // @[MapT.scala 15:7]
  assign O_6_0_t1b = op_O_6_0_t1b; // @[MapT.scala 15:7]
  assign O_7_0_t0b = op_O_7_0_t0b; // @[MapT.scala 15:7]
  assign O_7_0_t1b = op_O_7_0_t1b; // @[MapT.scala 15:7]
  assign O_8_0_t0b = op_O_8_0_t0b; // @[MapT.scala 15:7]
  assign O_8_0_t1b = op_O_8_0_t1b; // @[MapT.scala 15:7]
  assign O_9_0_t0b = op_O_9_0_t0b; // @[MapT.scala 15:7]
  assign O_9_0_t1b = op_O_9_0_t1b; // @[MapT.scala 15:7]
  assign O_10_0_t0b = op_O_10_0_t0b; // @[MapT.scala 15:7]
  assign O_10_0_t1b = op_O_10_0_t1b; // @[MapT.scala 15:7]
  assign O_11_0_t0b = op_O_11_0_t0b; // @[MapT.scala 15:7]
  assign O_11_0_t1b = op_O_11_0_t1b; // @[MapT.scala 15:7]
  assign O_12_0_t0b = op_O_12_0_t0b; // @[MapT.scala 15:7]
  assign O_12_0_t1b = op_O_12_0_t1b; // @[MapT.scala 15:7]
  assign O_13_0_t0b = op_O_13_0_t0b; // @[MapT.scala 15:7]
  assign O_13_0_t1b = op_O_13_0_t1b; // @[MapT.scala 15:7]
  assign O_14_0_t0b = op_O_14_0_t0b; // @[MapT.scala 15:7]
  assign O_14_0_t1b = op_O_14_0_t1b; // @[MapT.scala 15:7]
  assign O_15_0_t0b = op_O_15_0_t0b; // @[MapT.scala 15:7]
  assign O_15_0_t1b = op_O_15_0_t1b; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_t0b = I_0_t0b; // @[MapT.scala 14:10]
  assign op_I_0_t1b = I_0_t1b; // @[MapT.scala 14:10]
  assign op_I_1_t0b = I_1_t0b; // @[MapT.scala 14:10]
  assign op_I_1_t1b = I_1_t1b; // @[MapT.scala 14:10]
  assign op_I_2_t0b = I_2_t0b; // @[MapT.scala 14:10]
  assign op_I_2_t1b = I_2_t1b; // @[MapT.scala 14:10]
  assign op_I_3_t0b = I_3_t0b; // @[MapT.scala 14:10]
  assign op_I_3_t1b = I_3_t1b; // @[MapT.scala 14:10]
  assign op_I_4_t0b = I_4_t0b; // @[MapT.scala 14:10]
  assign op_I_4_t1b = I_4_t1b; // @[MapT.scala 14:10]
  assign op_I_5_t0b = I_5_t0b; // @[MapT.scala 14:10]
  assign op_I_5_t1b = I_5_t1b; // @[MapT.scala 14:10]
  assign op_I_6_t0b = I_6_t0b; // @[MapT.scala 14:10]
  assign op_I_6_t1b = I_6_t1b; // @[MapT.scala 14:10]
  assign op_I_7_t0b = I_7_t0b; // @[MapT.scala 14:10]
  assign op_I_7_t1b = I_7_t1b; // @[MapT.scala 14:10]
  assign op_I_8_t0b = I_8_t0b; // @[MapT.scala 14:10]
  assign op_I_8_t1b = I_8_t1b; // @[MapT.scala 14:10]
  assign op_I_9_t0b = I_9_t0b; // @[MapT.scala 14:10]
  assign op_I_9_t1b = I_9_t1b; // @[MapT.scala 14:10]
  assign op_I_10_t0b = I_10_t0b; // @[MapT.scala 14:10]
  assign op_I_10_t1b = I_10_t1b; // @[MapT.scala 14:10]
  assign op_I_11_t0b = I_11_t0b; // @[MapT.scala 14:10]
  assign op_I_11_t1b = I_11_t1b; // @[MapT.scala 14:10]
  assign op_I_12_t0b = I_12_t0b; // @[MapT.scala 14:10]
  assign op_I_12_t1b = I_12_t1b; // @[MapT.scala 14:10]
  assign op_I_13_t0b = I_13_t0b; // @[MapT.scala 14:10]
  assign op_I_13_t1b = I_13_t1b; // @[MapT.scala 14:10]
  assign op_I_14_t0b = I_14_t0b; // @[MapT.scala 14:10]
  assign op_I_14_t1b = I_14_t1b; // @[MapT.scala 14:10]
  assign op_I_15_t0b = I_15_t0b; // @[MapT.scala 14:10]
  assign op_I_15_t1b = I_15_t1b; // @[MapT.scala 14:10]
endmodule
module PartitionS_5(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t0b,
  input   I_0_0_t1b,
  input   I_1_0_t0b,
  input   I_1_0_t1b,
  input   I_2_0_t0b,
  input   I_2_0_t1b,
  input   I_3_0_t0b,
  input   I_3_0_t1b,
  input   I_4_0_t0b,
  input   I_4_0_t1b,
  input   I_5_0_t0b,
  input   I_5_0_t1b,
  input   I_6_0_t0b,
  input   I_6_0_t1b,
  input   I_7_0_t0b,
  input   I_7_0_t1b,
  input   I_8_0_t0b,
  input   I_8_0_t1b,
  input   I_9_0_t0b,
  input   I_9_0_t1b,
  input   I_10_0_t0b,
  input   I_10_0_t1b,
  input   I_11_0_t0b,
  input   I_11_0_t1b,
  input   I_12_0_t0b,
  input   I_12_0_t1b,
  input   I_13_0_t0b,
  input   I_13_0_t1b,
  input   I_14_0_t0b,
  input   I_14_0_t1b,
  input   I_15_0_t0b,
  input   I_15_0_t1b,
  output  O_0_0_0_t0b,
  output  O_0_0_0_t1b,
  output  O_1_0_0_t0b,
  output  O_1_0_0_t1b,
  output  O_2_0_0_t0b,
  output  O_2_0_0_t1b,
  output  O_3_0_0_t0b,
  output  O_3_0_0_t1b,
  output  O_4_0_0_t0b,
  output  O_4_0_0_t1b,
  output  O_5_0_0_t0b,
  output  O_5_0_0_t1b,
  output  O_6_0_0_t0b,
  output  O_6_0_0_t1b,
  output  O_7_0_0_t0b,
  output  O_7_0_0_t1b,
  output  O_8_0_0_t0b,
  output  O_8_0_0_t1b,
  output  O_9_0_0_t0b,
  output  O_9_0_0_t1b,
  output  O_10_0_0_t0b,
  output  O_10_0_0_t1b,
  output  O_11_0_0_t0b,
  output  O_11_0_0_t1b,
  output  O_12_0_0_t0b,
  output  O_12_0_0_t1b,
  output  O_13_0_0_t0b,
  output  O_13_0_0_t1b,
  output  O_14_0_0_t0b,
  output  O_14_0_0_t1b,
  output  O_15_0_0_t0b,
  output  O_15_0_0_t1b
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_t0b = I_0_0_t0b; // @[Partition.scala 15:39]
  assign O_0_0_0_t1b = I_0_0_t1b; // @[Partition.scala 15:39]
  assign O_1_0_0_t0b = I_1_0_t0b; // @[Partition.scala 15:39]
  assign O_1_0_0_t1b = I_1_0_t1b; // @[Partition.scala 15:39]
  assign O_2_0_0_t0b = I_2_0_t0b; // @[Partition.scala 15:39]
  assign O_2_0_0_t1b = I_2_0_t1b; // @[Partition.scala 15:39]
  assign O_3_0_0_t0b = I_3_0_t0b; // @[Partition.scala 15:39]
  assign O_3_0_0_t1b = I_3_0_t1b; // @[Partition.scala 15:39]
  assign O_4_0_0_t0b = I_4_0_t0b; // @[Partition.scala 15:39]
  assign O_4_0_0_t1b = I_4_0_t1b; // @[Partition.scala 15:39]
  assign O_5_0_0_t0b = I_5_0_t0b; // @[Partition.scala 15:39]
  assign O_5_0_0_t1b = I_5_0_t1b; // @[Partition.scala 15:39]
  assign O_6_0_0_t0b = I_6_0_t0b; // @[Partition.scala 15:39]
  assign O_6_0_0_t1b = I_6_0_t1b; // @[Partition.scala 15:39]
  assign O_7_0_0_t0b = I_7_0_t0b; // @[Partition.scala 15:39]
  assign O_7_0_0_t1b = I_7_0_t1b; // @[Partition.scala 15:39]
  assign O_8_0_0_t0b = I_8_0_t0b; // @[Partition.scala 15:39]
  assign O_8_0_0_t1b = I_8_0_t1b; // @[Partition.scala 15:39]
  assign O_9_0_0_t0b = I_9_0_t0b; // @[Partition.scala 15:39]
  assign O_9_0_0_t1b = I_9_0_t1b; // @[Partition.scala 15:39]
  assign O_10_0_0_t0b = I_10_0_t0b; // @[Partition.scala 15:39]
  assign O_10_0_0_t1b = I_10_0_t1b; // @[Partition.scala 15:39]
  assign O_11_0_0_t0b = I_11_0_t0b; // @[Partition.scala 15:39]
  assign O_11_0_0_t1b = I_11_0_t1b; // @[Partition.scala 15:39]
  assign O_12_0_0_t0b = I_12_0_t0b; // @[Partition.scala 15:39]
  assign O_12_0_0_t1b = I_12_0_t1b; // @[Partition.scala 15:39]
  assign O_13_0_0_t0b = I_13_0_t0b; // @[Partition.scala 15:39]
  assign O_13_0_0_t1b = I_13_0_t1b; // @[Partition.scala 15:39]
  assign O_14_0_0_t0b = I_14_0_t0b; // @[Partition.scala 15:39]
  assign O_14_0_0_t1b = I_14_0_t1b; // @[Partition.scala 15:39]
  assign O_15_0_0_t0b = I_15_0_t0b; // @[Partition.scala 15:39]
  assign O_15_0_0_t1b = I_15_0_t1b; // @[Partition.scala 15:39]
endmodule
module MapT_11(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t0b,
  input   I_0_0_t1b,
  input   I_1_0_t0b,
  input   I_1_0_t1b,
  input   I_2_0_t0b,
  input   I_2_0_t1b,
  input   I_3_0_t0b,
  input   I_3_0_t1b,
  input   I_4_0_t0b,
  input   I_4_0_t1b,
  input   I_5_0_t0b,
  input   I_5_0_t1b,
  input   I_6_0_t0b,
  input   I_6_0_t1b,
  input   I_7_0_t0b,
  input   I_7_0_t1b,
  input   I_8_0_t0b,
  input   I_8_0_t1b,
  input   I_9_0_t0b,
  input   I_9_0_t1b,
  input   I_10_0_t0b,
  input   I_10_0_t1b,
  input   I_11_0_t0b,
  input   I_11_0_t1b,
  input   I_12_0_t0b,
  input   I_12_0_t1b,
  input   I_13_0_t0b,
  input   I_13_0_t1b,
  input   I_14_0_t0b,
  input   I_14_0_t1b,
  input   I_15_0_t0b,
  input   I_15_0_t1b,
  output  O_0_0_0_t0b,
  output  O_0_0_0_t1b,
  output  O_1_0_0_t0b,
  output  O_1_0_0_t1b,
  output  O_2_0_0_t0b,
  output  O_2_0_0_t1b,
  output  O_3_0_0_t0b,
  output  O_3_0_0_t1b,
  output  O_4_0_0_t0b,
  output  O_4_0_0_t1b,
  output  O_5_0_0_t0b,
  output  O_5_0_0_t1b,
  output  O_6_0_0_t0b,
  output  O_6_0_0_t1b,
  output  O_7_0_0_t0b,
  output  O_7_0_0_t1b,
  output  O_8_0_0_t0b,
  output  O_8_0_0_t1b,
  output  O_9_0_0_t0b,
  output  O_9_0_0_t1b,
  output  O_10_0_0_t0b,
  output  O_10_0_0_t1b,
  output  O_11_0_0_t0b,
  output  O_11_0_0_t1b,
  output  O_12_0_0_t0b,
  output  O_12_0_0_t1b,
  output  O_13_0_0_t0b,
  output  O_13_0_0_t1b,
  output  O_14_0_0_t0b,
  output  O_14_0_0_t1b,
  output  O_15_0_0_t0b,
  output  O_15_0_0_t1b
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire  op_I_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_1_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_1_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_2_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_2_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_3_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_3_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_4_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_4_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_5_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_5_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_6_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_6_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_7_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_7_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_8_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_8_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_9_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_9_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_10_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_10_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_11_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_11_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_12_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_12_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_13_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_13_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_14_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_14_0_t1b; // @[MapT.scala 8:20]
  wire  op_I_15_0_t0b; // @[MapT.scala 8:20]
  wire  op_I_15_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_0_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_0_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_1_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_1_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_2_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_2_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_3_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_3_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_4_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_4_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_5_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_5_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_6_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_6_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_7_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_7_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_8_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_8_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_9_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_9_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_10_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_10_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_11_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_11_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_12_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_12_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_13_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_13_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_14_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_14_0_0_t1b; // @[MapT.scala 8:20]
  wire  op_O_15_0_0_t0b; // @[MapT.scala 8:20]
  wire  op_O_15_0_0_t1b; // @[MapT.scala 8:20]
  PartitionS_5 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_t0b(op_I_0_0_t0b),
    .I_0_0_t1b(op_I_0_0_t1b),
    .I_1_0_t0b(op_I_1_0_t0b),
    .I_1_0_t1b(op_I_1_0_t1b),
    .I_2_0_t0b(op_I_2_0_t0b),
    .I_2_0_t1b(op_I_2_0_t1b),
    .I_3_0_t0b(op_I_3_0_t0b),
    .I_3_0_t1b(op_I_3_0_t1b),
    .I_4_0_t0b(op_I_4_0_t0b),
    .I_4_0_t1b(op_I_4_0_t1b),
    .I_5_0_t0b(op_I_5_0_t0b),
    .I_5_0_t1b(op_I_5_0_t1b),
    .I_6_0_t0b(op_I_6_0_t0b),
    .I_6_0_t1b(op_I_6_0_t1b),
    .I_7_0_t0b(op_I_7_0_t0b),
    .I_7_0_t1b(op_I_7_0_t1b),
    .I_8_0_t0b(op_I_8_0_t0b),
    .I_8_0_t1b(op_I_8_0_t1b),
    .I_9_0_t0b(op_I_9_0_t0b),
    .I_9_0_t1b(op_I_9_0_t1b),
    .I_10_0_t0b(op_I_10_0_t0b),
    .I_10_0_t1b(op_I_10_0_t1b),
    .I_11_0_t0b(op_I_11_0_t0b),
    .I_11_0_t1b(op_I_11_0_t1b),
    .I_12_0_t0b(op_I_12_0_t0b),
    .I_12_0_t1b(op_I_12_0_t1b),
    .I_13_0_t0b(op_I_13_0_t0b),
    .I_13_0_t1b(op_I_13_0_t1b),
    .I_14_0_t0b(op_I_14_0_t0b),
    .I_14_0_t1b(op_I_14_0_t1b),
    .I_15_0_t0b(op_I_15_0_t0b),
    .I_15_0_t1b(op_I_15_0_t1b),
    .O_0_0_0_t0b(op_O_0_0_0_t0b),
    .O_0_0_0_t1b(op_O_0_0_0_t1b),
    .O_1_0_0_t0b(op_O_1_0_0_t0b),
    .O_1_0_0_t1b(op_O_1_0_0_t1b),
    .O_2_0_0_t0b(op_O_2_0_0_t0b),
    .O_2_0_0_t1b(op_O_2_0_0_t1b),
    .O_3_0_0_t0b(op_O_3_0_0_t0b),
    .O_3_0_0_t1b(op_O_3_0_0_t1b),
    .O_4_0_0_t0b(op_O_4_0_0_t0b),
    .O_4_0_0_t1b(op_O_4_0_0_t1b),
    .O_5_0_0_t0b(op_O_5_0_0_t0b),
    .O_5_0_0_t1b(op_O_5_0_0_t1b),
    .O_6_0_0_t0b(op_O_6_0_0_t0b),
    .O_6_0_0_t1b(op_O_6_0_0_t1b),
    .O_7_0_0_t0b(op_O_7_0_0_t0b),
    .O_7_0_0_t1b(op_O_7_0_0_t1b),
    .O_8_0_0_t0b(op_O_8_0_0_t0b),
    .O_8_0_0_t1b(op_O_8_0_0_t1b),
    .O_9_0_0_t0b(op_O_9_0_0_t0b),
    .O_9_0_0_t1b(op_O_9_0_0_t1b),
    .O_10_0_0_t0b(op_O_10_0_0_t0b),
    .O_10_0_0_t1b(op_O_10_0_0_t1b),
    .O_11_0_0_t0b(op_O_11_0_0_t0b),
    .O_11_0_0_t1b(op_O_11_0_0_t1b),
    .O_12_0_0_t0b(op_O_12_0_0_t0b),
    .O_12_0_0_t1b(op_O_12_0_0_t1b),
    .O_13_0_0_t0b(op_O_13_0_0_t0b),
    .O_13_0_0_t1b(op_O_13_0_0_t1b),
    .O_14_0_0_t0b(op_O_14_0_0_t0b),
    .O_14_0_0_t1b(op_O_14_0_0_t1b),
    .O_15_0_0_t0b(op_O_15_0_0_t0b),
    .O_15_0_0_t1b(op_O_15_0_0_t1b)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_t0b = op_O_0_0_0_t0b; // @[MapT.scala 15:7]
  assign O_0_0_0_t1b = op_O_0_0_0_t1b; // @[MapT.scala 15:7]
  assign O_1_0_0_t0b = op_O_1_0_0_t0b; // @[MapT.scala 15:7]
  assign O_1_0_0_t1b = op_O_1_0_0_t1b; // @[MapT.scala 15:7]
  assign O_2_0_0_t0b = op_O_2_0_0_t0b; // @[MapT.scala 15:7]
  assign O_2_0_0_t1b = op_O_2_0_0_t1b; // @[MapT.scala 15:7]
  assign O_3_0_0_t0b = op_O_3_0_0_t0b; // @[MapT.scala 15:7]
  assign O_3_0_0_t1b = op_O_3_0_0_t1b; // @[MapT.scala 15:7]
  assign O_4_0_0_t0b = op_O_4_0_0_t0b; // @[MapT.scala 15:7]
  assign O_4_0_0_t1b = op_O_4_0_0_t1b; // @[MapT.scala 15:7]
  assign O_5_0_0_t0b = op_O_5_0_0_t0b; // @[MapT.scala 15:7]
  assign O_5_0_0_t1b = op_O_5_0_0_t1b; // @[MapT.scala 15:7]
  assign O_6_0_0_t0b = op_O_6_0_0_t0b; // @[MapT.scala 15:7]
  assign O_6_0_0_t1b = op_O_6_0_0_t1b; // @[MapT.scala 15:7]
  assign O_7_0_0_t0b = op_O_7_0_0_t0b; // @[MapT.scala 15:7]
  assign O_7_0_0_t1b = op_O_7_0_0_t1b; // @[MapT.scala 15:7]
  assign O_8_0_0_t0b = op_O_8_0_0_t0b; // @[MapT.scala 15:7]
  assign O_8_0_0_t1b = op_O_8_0_0_t1b; // @[MapT.scala 15:7]
  assign O_9_0_0_t0b = op_O_9_0_0_t0b; // @[MapT.scala 15:7]
  assign O_9_0_0_t1b = op_O_9_0_0_t1b; // @[MapT.scala 15:7]
  assign O_10_0_0_t0b = op_O_10_0_0_t0b; // @[MapT.scala 15:7]
  assign O_10_0_0_t1b = op_O_10_0_0_t1b; // @[MapT.scala 15:7]
  assign O_11_0_0_t0b = op_O_11_0_0_t0b; // @[MapT.scala 15:7]
  assign O_11_0_0_t1b = op_O_11_0_0_t1b; // @[MapT.scala 15:7]
  assign O_12_0_0_t0b = op_O_12_0_0_t0b; // @[MapT.scala 15:7]
  assign O_12_0_0_t1b = op_O_12_0_0_t1b; // @[MapT.scala 15:7]
  assign O_13_0_0_t0b = op_O_13_0_0_t0b; // @[MapT.scala 15:7]
  assign O_13_0_0_t1b = op_O_13_0_0_t1b; // @[MapT.scala 15:7]
  assign O_14_0_0_t0b = op_O_14_0_0_t0b; // @[MapT.scala 15:7]
  assign O_14_0_0_t1b = op_O_14_0_0_t1b; // @[MapT.scala 15:7]
  assign O_15_0_0_t0b = op_O_15_0_0_t0b; // @[MapT.scala 15:7]
  assign O_15_0_0_t1b = op_O_15_0_0_t1b; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_t0b = I_0_0_t0b; // @[MapT.scala 14:10]
  assign op_I_0_0_t1b = I_0_0_t1b; // @[MapT.scala 14:10]
  assign op_I_1_0_t0b = I_1_0_t0b; // @[MapT.scala 14:10]
  assign op_I_1_0_t1b = I_1_0_t1b; // @[MapT.scala 14:10]
  assign op_I_2_0_t0b = I_2_0_t0b; // @[MapT.scala 14:10]
  assign op_I_2_0_t1b = I_2_0_t1b; // @[MapT.scala 14:10]
  assign op_I_3_0_t0b = I_3_0_t0b; // @[MapT.scala 14:10]
  assign op_I_3_0_t1b = I_3_0_t1b; // @[MapT.scala 14:10]
  assign op_I_4_0_t0b = I_4_0_t0b; // @[MapT.scala 14:10]
  assign op_I_4_0_t1b = I_4_0_t1b; // @[MapT.scala 14:10]
  assign op_I_5_0_t0b = I_5_0_t0b; // @[MapT.scala 14:10]
  assign op_I_5_0_t1b = I_5_0_t1b; // @[MapT.scala 14:10]
  assign op_I_6_0_t0b = I_6_0_t0b; // @[MapT.scala 14:10]
  assign op_I_6_0_t1b = I_6_0_t1b; // @[MapT.scala 14:10]
  assign op_I_7_0_t0b = I_7_0_t0b; // @[MapT.scala 14:10]
  assign op_I_7_0_t1b = I_7_0_t1b; // @[MapT.scala 14:10]
  assign op_I_8_0_t0b = I_8_0_t0b; // @[MapT.scala 14:10]
  assign op_I_8_0_t1b = I_8_0_t1b; // @[MapT.scala 14:10]
  assign op_I_9_0_t0b = I_9_0_t0b; // @[MapT.scala 14:10]
  assign op_I_9_0_t1b = I_9_0_t1b; // @[MapT.scala 14:10]
  assign op_I_10_0_t0b = I_10_0_t0b; // @[MapT.scala 14:10]
  assign op_I_10_0_t1b = I_10_0_t1b; // @[MapT.scala 14:10]
  assign op_I_11_0_t0b = I_11_0_t0b; // @[MapT.scala 14:10]
  assign op_I_11_0_t1b = I_11_0_t1b; // @[MapT.scala 14:10]
  assign op_I_12_0_t0b = I_12_0_t0b; // @[MapT.scala 14:10]
  assign op_I_12_0_t1b = I_12_0_t1b; // @[MapT.scala 14:10]
  assign op_I_13_0_t0b = I_13_0_t0b; // @[MapT.scala 14:10]
  assign op_I_13_0_t1b = I_13_0_t1b; // @[MapT.scala 14:10]
  assign op_I_14_0_t0b = I_14_0_t0b; // @[MapT.scala 14:10]
  assign op_I_14_0_t1b = I_14_0_t1b; // @[MapT.scala 14:10]
  assign op_I_15_0_t0b = I_15_0_t0b; // @[MapT.scala 14:10]
  assign op_I_15_0_t1b = I_15_0_t1b; // @[MapT.scala 14:10]
endmodule
module FIFO_1(
  input   clock,
  input   reset,
  input   valid_up,
  output  valid_down,
  input   I_0_0_0_t0b,
  input   I_0_0_0_t1b,
  input   I_1_0_0_t0b,
  input   I_1_0_0_t1b,
  input   I_2_0_0_t0b,
  input   I_2_0_0_t1b,
  input   I_3_0_0_t0b,
  input   I_3_0_0_t1b,
  input   I_4_0_0_t0b,
  input   I_4_0_0_t1b,
  input   I_5_0_0_t0b,
  input   I_5_0_0_t1b,
  input   I_6_0_0_t0b,
  input   I_6_0_0_t1b,
  input   I_7_0_0_t0b,
  input   I_7_0_0_t1b,
  input   I_8_0_0_t0b,
  input   I_8_0_0_t1b,
  input   I_9_0_0_t0b,
  input   I_9_0_0_t1b,
  input   I_10_0_0_t0b,
  input   I_10_0_0_t1b,
  input   I_11_0_0_t0b,
  input   I_11_0_0_t1b,
  input   I_12_0_0_t0b,
  input   I_12_0_0_t1b,
  input   I_13_0_0_t0b,
  input   I_13_0_0_t1b,
  input   I_14_0_0_t0b,
  input   I_14_0_0_t1b,
  input   I_15_0_0_t0b,
  input   I_15_0_0_t1b,
  output  O_0_0_0_t0b,
  output  O_0_0_0_t1b,
  output  O_1_0_0_t0b,
  output  O_1_0_0_t1b,
  output  O_2_0_0_t0b,
  output  O_2_0_0_t1b,
  output  O_3_0_0_t0b,
  output  O_3_0_0_t1b,
  output  O_4_0_0_t0b,
  output  O_4_0_0_t1b,
  output  O_5_0_0_t0b,
  output  O_5_0_0_t1b,
  output  O_6_0_0_t0b,
  output  O_6_0_0_t1b,
  output  O_7_0_0_t0b,
  output  O_7_0_0_t1b,
  output  O_8_0_0_t0b,
  output  O_8_0_0_t1b,
  output  O_9_0_0_t0b,
  output  O_9_0_0_t1b,
  output  O_10_0_0_t0b,
  output  O_10_0_0_t1b,
  output  O_11_0_0_t0b,
  output  O_11_0_0_t1b,
  output  O_12_0_0_t0b,
  output  O_12_0_0_t1b,
  output  O_13_0_0_t0b,
  output  O_13_0_0_t1b,
  output  O_14_0_0_t0b,
  output  O_14_0_0_t1b,
  output  O_15_0_0_t0b,
  output  O_15_0_0_t1b
);
  reg  _T__0_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg  _T__0_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg  _T__1_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg  _T__1_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg  _T__2_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg  _T__2_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg  _T__3_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg  _T__3_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg  _T__4_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg  _T__4_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg  _T__5_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg  _T__5_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg  _T__6_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg  _T__6_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg  _T__7_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg  _T__7_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T__8_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_16;
  reg  _T__8_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_17;
  reg  _T__9_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_18;
  reg  _T__9_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_19;
  reg  _T__10_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_20;
  reg  _T__10_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_21;
  reg  _T__11_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_22;
  reg  _T__11_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_23;
  reg  _T__12_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_24;
  reg  _T__12_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_25;
  reg  _T__13_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_26;
  reg  _T__13_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_27;
  reg  _T__14_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_28;
  reg  _T__14_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_29;
  reg  _T__15_0_0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_30;
  reg  _T__15_0_0_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_31;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_32;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_0_0_t0b = _T__0_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_0_0_0_t1b = _T__0_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_1_0_0_t0b = _T__1_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_1_0_0_t1b = _T__1_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_2_0_0_t0b = _T__2_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_2_0_0_t1b = _T__2_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_3_0_0_t0b = _T__3_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_3_0_0_t1b = _T__3_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_4_0_0_t0b = _T__4_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_4_0_0_t1b = _T__4_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_5_0_0_t0b = _T__5_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_5_0_0_t1b = _T__5_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_6_0_0_t0b = _T__6_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_6_0_0_t1b = _T__6_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_7_0_0_t0b = _T__7_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_7_0_0_t1b = _T__7_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_8_0_0_t0b = _T__8_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_8_0_0_t1b = _T__8_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_9_0_0_t0b = _T__9_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_9_0_0_t1b = _T__9_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_10_0_0_t0b = _T__10_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_10_0_0_t1b = _T__10_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_11_0_0_t0b = _T__11_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_11_0_0_t1b = _T__11_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_12_0_0_t0b = _T__12_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_12_0_0_t1b = _T__12_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_13_0_0_t0b = _T__13_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_13_0_0_t1b = _T__13_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_14_0_0_t0b = _T__14_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_14_0_0_t1b = _T__14_0_0_t1b; // @[FIFO.scala 14:7]
  assign O_15_0_0_t0b = _T__15_0_0_t0b; // @[FIFO.scala 14:7]
  assign O_15_0_0_t1b = _T__15_0_0_t1b; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_0_0_t0b = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__0_0_0_t1b = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__1_0_0_t0b = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__1_0_0_t1b = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__2_0_0_t0b = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__2_0_0_t1b = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__3_0_0_t0b = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__3_0_0_t1b = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__4_0_0_t0b = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__4_0_0_t1b = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__5_0_0_t0b = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__5_0_0_t1b = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__6_0_0_t0b = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__6_0_0_t1b = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__7_0_0_t0b = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__7_0_0_t1b = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T__8_0_0_t0b = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T__8_0_0_t1b = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__9_0_0_t0b = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__9_0_0_t1b = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T__10_0_0_t0b = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T__10_0_0_t1b = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__11_0_0_t0b = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__11_0_0_t1b = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T__12_0_0_t0b = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T__12_0_0_t1b = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__13_0_0_t0b = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__13_0_0_t1b = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T__14_0_0_t0b = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T__14_0_0_t1b = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__15_0_0_t0b = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__15_0_0_t1b = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_0_0_t0b <= I_0_0_0_t0b;
    _T__0_0_0_t1b <= I_0_0_0_t1b;
    _T__1_0_0_t0b <= I_1_0_0_t0b;
    _T__1_0_0_t1b <= I_1_0_0_t1b;
    _T__2_0_0_t0b <= I_2_0_0_t0b;
    _T__2_0_0_t1b <= I_2_0_0_t1b;
    _T__3_0_0_t0b <= I_3_0_0_t0b;
    _T__3_0_0_t1b <= I_3_0_0_t1b;
    _T__4_0_0_t0b <= I_4_0_0_t0b;
    _T__4_0_0_t1b <= I_4_0_0_t1b;
    _T__5_0_0_t0b <= I_5_0_0_t0b;
    _T__5_0_0_t1b <= I_5_0_0_t1b;
    _T__6_0_0_t0b <= I_6_0_0_t0b;
    _T__6_0_0_t1b <= I_6_0_0_t1b;
    _T__7_0_0_t0b <= I_7_0_0_t0b;
    _T__7_0_0_t1b <= I_7_0_0_t1b;
    _T__8_0_0_t0b <= I_8_0_0_t0b;
    _T__8_0_0_t1b <= I_8_0_0_t1b;
    _T__9_0_0_t0b <= I_9_0_0_t0b;
    _T__9_0_0_t1b <= I_9_0_0_t1b;
    _T__10_0_0_t0b <= I_10_0_0_t0b;
    _T__10_0_0_t1b <= I_10_0_0_t1b;
    _T__11_0_0_t0b <= I_11_0_0_t0b;
    _T__11_0_0_t1b <= I_11_0_0_t1b;
    _T__12_0_0_t0b <= I_12_0_0_t0b;
    _T__12_0_0_t1b <= I_12_0_0_t1b;
    _T__13_0_0_t0b <= I_13_0_0_t0b;
    _T__13_0_0_t1b <= I_13_0_0_t1b;
    _T__14_0_0_t0b <= I_14_0_0_t0b;
    _T__14_0_0_t1b <= I_14_0_0_t1b;
    _T__15_0_0_t0b <= I_15_0_0_t0b;
    _T__15_0_0_t1b <= I_15_0_0_t1b;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module Fst(
  input   valid_up,
  output  valid_down,
  input   I_t0b,
  output  O
);
  assign valid_down = valid_up; // @[Tuple.scala 59:14]
  assign O = I_t0b; // @[Tuple.scala 58:5]
endmodule
module MapS_6(
  input   valid_up,
  output  valid_down,
  input   I_0_t0b,
  output  O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_t0b; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  Fst fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
endmodule
module MapS_7(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t0b,
  output  O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire  fst_op_O_0; // @[MapS.scala 9:22]
  MapS_6 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
endmodule
module FIFO_2(
  input   clock,
  input   reset,
  input   valid_up,
  output  valid_down,
  input   I_0_0,
  output  O_0_0
);
  reg  _T_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire  _T_0_0__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire  _T_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T_0_0__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [1:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T_0_0__T_15_addr = _T_0_0__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_15_data = _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0__T_15_data = _T_0_0__T_15_addr >= 2'h3 ? _RAND_1[0:0] : _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_5_data = I_0_0;
  assign _T_0_0__T_5_addr = value_2;
  assign _T_0_0__T_5_mask = 1'h1;
  assign _T_0_0__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_9 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0 = _T_0_0__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_0_0__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_0_0__T_15_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_2 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_0_0__T_5_en & _T_0_0__T_5_mask) begin
      _T_0_0[_T_0_0__T_5_addr] <= _T_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module Snd(
  input   valid_up,
  output  valid_down,
  input   I_t1b,
  output  O
);
  assign valid_down = valid_up; // @[Tuple.scala 67:14]
  assign O = I_t1b; // @[Tuple.scala 66:5]
endmodule
module MapS_8(
  input   valid_up,
  output  valid_down,
  input   I_0_t1b,
  output  O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_t1b; // @[MapS.scala 9:22]
  wire  fst_op_O; // @[MapS.scala 9:22]
  Snd fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_9(
  input   valid_up,
  output  valid_down,
  input   I_0_0_t1b,
  output  O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire  fst_op_O_0; // @[MapS.scala 9:22]
  MapS_8 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module DownS(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_1_0,
  input  [31:0] I_1_1,
  input  [31:0] I_1_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0_0 = I_1_0; // @[Downsample.scala 12:8]
  assign O_0_1 = I_1_1; // @[Downsample.scala 12:8]
  assign O_0_2 = I_1_2; // @[Downsample.scala 12:8]
endmodule
module DownS_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  output [31:0] O_0
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0 = I_0; // @[Downsample.scala 12:8]
endmodule
module MapS_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  DownS_1 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
endmodule
module DownS_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_2,
  output [31:0] O_0
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0 = I_2; // @[Downsample.scala 12:8]
endmodule
module MapS_11(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_2,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  DownS_2 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
endmodule
module Map2S_9(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I1_0,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_9 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Add(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 108:14]
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 106:7]
endmodule
module MapS_12(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_0_t1b,
  output [31:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  Add fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_13(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_12 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_2(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n182_valid_up; // @[Top.scala 68:22]
  wire  n182_valid_down; // @[Top.scala 68:22]
  wire [31:0] n182_I0; // @[Top.scala 68:22]
  wire [7:0] n182_I1; // @[Top.scala 68:22]
  wire [31:0] n182_O_t0b; // @[Top.scala 68:22]
  wire [7:0] n182_O_t1b; // @[Top.scala 68:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple_1 n182 ( // @[Top.scala 68:22]
    .valid_up(n182_valid_up),
    .valid_down(n182_valid_down),
    .I0(n182_I0),
    .I1(n182_I1),
    .O_t0b(n182_O_t0b),
    .O_t1b(n182_O_t1b)
  );
  assign valid_down = n182_valid_down; // @[Top.scala 73:16]
  assign O_t0b = n182_O_t0b; // @[Top.scala 72:7]
  assign O_t1b = n182_O_t1b; // @[Top.scala 72:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n182_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 71:19]
  assign n182_I0 = I; // @[Top.scala 69:13]
  assign n182_I1 = 8'h1; // @[Top.scala 70:13]
endmodule
module MapS_14(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  output [31:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[MapS.scala 9:22]
  Module_2 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_t0b = fst_op_O_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b = fst_op_O_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
endmodule
module MapS_15(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[MapS.scala 9:22]
  MapS_14 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
endmodule
module MapS_16(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [7:0]  I_0_t1b,
  output [31:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_17(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [7:0]  I_0_0_t1b,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_16 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module DownS_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_1,
  output [31:0] O_0
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0 = I_1; // @[Downsample.scala 12:8]
endmodule
module MapS_18(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_1,
  output [31:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  DownS_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_1(fst_op_I_1),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
endmodule
module DownS_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0_0 = I_0_0; // @[Downsample.scala 12:8]
  assign O_0_1 = I_0_1; // @[Downsample.scala 12:8]
  assign O_0_2 = I_0_2; // @[Downsample.scala 12:8]
endmodule
module DownS_6(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_2_0,
  input  [31:0] I_2_1,
  input  [31:0] I_2_2,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  assign valid_down = valid_up; // @[Downsample.scala 13:14]
  assign O_0_0 = I_2_0; // @[Downsample.scala 12:8]
  assign O_0_1 = I_2_1; // @[Downsample.scala 12:8]
  assign O_0_2 = I_2_2; // @[Downsample.scala 12:8]
endmodule
module AtomTuple_10(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0,
  input  [31:0] I1_t0b,
  input  [31:0] I1_t1b,
  output [31:0] O_t0b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b = I1_t1b; // @[Tuple.scala 50:9]
endmodule
module Map2S_15(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I1_0_t0b,
  input  [31:0] I1_0_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b; // @[Map2S.scala 9:22]
  AtomTuple_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1_t0b(fst_op_I1_t0b),
    .I1_t1b(fst_op_I1_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b(fst_op_O_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b = fst_op_O_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b = I1_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b = I1_0_t1b; // @[Map2S.scala 18:13]
endmodule
module Map2S_16(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I1_0_0_t0b,
  input  [31:0] I1_0_0_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b; // @[Map2S.scala 9:22]
  Map2S_15 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0_t0b(fst_op_I1_0_t0b),
    .I1_0_t1b(fst_op_I1_0_t1b),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b_t0b(fst_op_O_0_t1b_t0b),
    .O_0_t1b_t1b(fst_op_O_0_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b = fst_op_O_0_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b = fst_op_O_0_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_t0b = I1_0_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b = I1_0_0_t1b; // @[Map2S.scala 18:13]
endmodule
module FIFO_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  reg [31:0] _T_0_0_t0b [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [31:0] _T_0_0_t0b__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t0b__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [31:0] _T_0_0_t0b__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t0b__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0_t0b__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0_t0b__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0_t0b__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T_0_0_t0b__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [31:0] _T_0_0_t1b_t0b [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [31:0] _T_0_0_t1b_t0b__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t0b__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [31:0] _T_0_0_t1b_t0b__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t0b__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t0b__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t0b__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0_t1b_t0b__T_15_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [1:0] _T_0_0_t1b_t0b__T_15_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [31:0] _T_0_0_t1b_t1b [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [31:0] _T_0_0_t1b_t1b__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t1b__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [31:0] _T_0_0_t1b_t1b__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0_t1b_t1b__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t1b__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0_t1b_t1b__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0_t1b_t1b__T_15_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [1:0] _T_0_0_t1b_t1b__T_15_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_12;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_13;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_14;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [1:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T_0_0_t0b__T_15_addr = _T_0_0_t0b__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t0b__T_15_data = _T_0_0_t0b[_T_0_0_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0_t0b__T_15_data = _T_0_0_t0b__T_15_addr >= 2'h3 ? _RAND_1[31:0] : _T_0_0_t0b[_T_0_0_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t0b__T_5_data = I_0_0_t0b;
  assign _T_0_0_t0b__T_5_addr = value_2;
  assign _T_0_0_t0b__T_5_mask = 1'h1;
  assign _T_0_0_t0b__T_5_en = valid_up;
  assign _T_0_0_t1b_t0b__T_15_addr = _T_0_0_t1b_t0b__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t0b__T_15_data = _T_0_0_t1b_t0b[_T_0_0_t1b_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0_t1b_t0b__T_15_data = _T_0_0_t1b_t0b__T_15_addr >= 2'h3 ? _RAND_5[31:0] : _T_0_0_t1b_t0b[_T_0_0_t1b_t0b__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t0b__T_5_data = I_0_0_t1b_t0b;
  assign _T_0_0_t1b_t0b__T_5_addr = value_2;
  assign _T_0_0_t1b_t0b__T_5_mask = 1'h1;
  assign _T_0_0_t1b_t0b__T_5_en = valid_up;
  assign _T_0_0_t1b_t1b__T_15_addr = _T_0_0_t1b_t1b__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t1b__T_15_data = _T_0_0_t1b_t1b[_T_0_0_t1b_t1b__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0_t1b_t1b__T_15_data = _T_0_0_t1b_t1b__T_15_addr >= 2'h3 ? _RAND_9[31:0] : _T_0_0_t1b_t1b[_T_0_0_t1b_t1b__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0_t1b_t1b__T_5_data = I_0_0_t1b_t1b;
  assign _T_0_0_t1b_t1b__T_5_addr = value_2;
  assign _T_0_0_t1b_t1b__T_5_mask = 1'h1;
  assign _T_0_0_t1b_t1b__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_9 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0_t0b = _T_0_0_t0b__T_15_data; // @[FIFO.scala 43:11]
  assign O_0_0_t1b_t0b = _T_0_0_t1b_t0b__T_15_data; // @[FIFO.scala 43:11]
  assign O_0_0_t1b_t1b = _T_0_0_t1b_t1b__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0_t0b[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_0_0_t0b__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_0_0_t0b__T_15_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0_t1b_t0b[initvar] = _RAND_4[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_0_0_t1b_t0b__T_15_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_0_0_t1b_t0b__T_15_addr_pipe_0 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0_t1b_t1b[initvar] = _RAND_8[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_0_0_t1b_t1b__T_15_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_0_0_t1b_t1b__T_15_addr_pipe_0 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  value = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  value_1 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  value_2 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_0_0_t0b__T_5_en & _T_0_0_t0b__T_5_mask) begin
      _T_0_0_t0b[_T_0_0_t0b__T_5_addr] <= _T_0_0_t0b__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0_t0b__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0_t0b__T_15_addr_pipe_0 <= value_1;
    end
    if(_T_0_0_t1b_t0b__T_5_en & _T_0_0_t1b_t0b__T_5_mask) begin
      _T_0_0_t1b_t0b[_T_0_0_t1b_t0b__T_5_addr] <= _T_0_0_t1b_t0b__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0_t1b_t0b__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0_t1b_t0b__T_15_addr_pipe_0 <= value_1;
    end
    if(_T_0_0_t1b_t1b__T_5_en & _T_0_0_t1b_t1b__T_5_mask) begin
      _T_0_0_t1b_t1b[_T_0_0_t1b_t1b__T_5_addr] <= _T_0_0_t1b_t1b__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0_t1b_t1b__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0_t1b_t1b__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module FIFO_5(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0
);
  reg [31:0] _T_0_0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [31:0] _T_0_0__T_15_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_15_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [31:0] _T_0_0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T_0_0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T_0_0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T_0_0__T_15_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T_0_0__T_15_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_4;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_9; // @[Counter.scala 38:22]
  wire  _T_10; // @[FIFO.scala 42:39]
  wire  _T_16; // @[Counter.scala 37:24]
  wire [1:0] _T_18; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  assign _T_0_0__T_15_addr = _T_0_0__T_15_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_15_data = _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T_0_0__T_15_data = _T_0_0__T_15_addr >= 2'h3 ? _RAND_1[31:0] : _T_0_0[_T_0_0__T_15_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_0_0__T_5_data = I_0_0;
  assign _T_0_0__T_5_addr = value_2;
  assign _T_0_0__T_5_mask = 1'h1;
  assign _T_0_0__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_9 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_10 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_16 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_18 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_10 & _T_10; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0_0 = _T_0_0__T_15_data; // @[FIFO.scala 43:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T_0_0[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_0_0__T_15_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_0_0__T_15_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  value = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value_1 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  value_2 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_0_0__T_5_en & _T_0_0__T_5_mask) begin
      _T_0_0[_T_0_0__T_5_addr] <= _T_0_0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T_0_0__T_15_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T_0_0__T_15_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_9;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_10) begin
        if (_T_16) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
  end
endmodule
module Map2S_17(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I1_0,
  output [31:0] O_0_0,
  output [31:0] O_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_18(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  Map2S_17 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_19(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I1_0,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2; // @[Map2S.scala 9:22]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_20(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  Map2S_19 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module SSeqTupleAppender_5(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0,
  input  [31:0] I0_1,
  input  [31:0] I0_2,
  input  [31:0] I1,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I0_2; // @[Tuple.scala 24:34]
  assign O_3 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_21(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I1_0,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_0_3
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_3; // @[Map2S.scala 9:22]
  SSeqTupleAppender_5 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2),
    .O_3(fst_op_O_3)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_0_3 = fst_op_O_3; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_22(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I1_0_0,
  output [31:0] O_0_0_0,
  output [31:0] O_0_0_1,
  output [31:0] O_0_0_2,
  output [31:0] O_0_0_3
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_3; // @[Map2S.scala 9:22]
  Map2S_21 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I1_0(fst_op_I1_0),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_0_3(fst_op_O_0_3)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_0_3 = fst_op_O_0_3; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module SSeqTupleToSSeq_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
  assign O_3 = I_3; // @[Tuple.scala 41:5]
endmodule
module Remove1S_4(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_0_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_I_3; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  wire [31:0] op_inst_O_3; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_4 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .I_3(op_inst_I_3),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2),
    .O_3(op_inst_O_3)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign O_3 = op_inst_O_3; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_3 = I_0_3; // @[Remove1S.scala 13:13]
endmodule
module MapS_27(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_0_3,
  output [31:0] O_0_0,
  output [31:0] O_0_1,
  output [31:0] O_0_2,
  output [31:0] O_0_3
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_3; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_3; // @[MapS.scala 9:22]
  Remove1S_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_0_3(fst_op_I_0_3),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2),
    .O_3(fst_op_O_3)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_0_3 = fst_op_O_3; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_3 = I_0_0_3; // @[MapS.scala 16:12]
endmodule
module AddNoValid(
  input  [31:0] I_t0b,
  input  [31:0] I_t1b,
  output [31:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg [31:0] _T_4; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_5;
  reg  _T_6; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_6;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  AddNoValid AddNoValid_2 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_2_I_t0b),
    .I_t1b(AddNoValid_2_I_t1b),
    .O(AddNoValid_2_O)
  );
  assign valid_down = _T_6; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = AddNoValid_2_O; // @[ReduceS.scala 31:18]
  assign AddNoValid_1_I_t1b = _T_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t0b = _T_4; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t1b = _T_3; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    _T_4 <= I_3;
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= valid_up;
    end
    _T_6 <= _T_5;
  end
endmodule
module MapS_28(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_0_3,
  output [31:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_3; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .I_3(fst_op_I_3),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_3 = I_0_3; // @[MapS.scala 16:12]
endmodule
module InitialDelayCounter_2(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h3; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h3; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_4(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I,
  output [31:0] O_t0b,
  output [7:0]  O_t1b
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n274_valid_up; // @[Top.scala 92:22]
  wire  n274_valid_down; // @[Top.scala 92:22]
  wire [31:0] n274_I0; // @[Top.scala 92:22]
  wire [7:0] n274_I1; // @[Top.scala 92:22]
  wire [31:0] n274_O_t0b; // @[Top.scala 92:22]
  wire [7:0] n274_O_t1b; // @[Top.scala 92:22]
  InitialDelayCounter_2 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple_1 n274 ( // @[Top.scala 92:22]
    .valid_up(n274_valid_up),
    .valid_down(n274_valid_down),
    .I0(n274_I0),
    .I1(n274_I1),
    .O_t0b(n274_O_t0b),
    .O_t1b(n274_O_t1b)
  );
  assign valid_down = n274_valid_down; // @[Top.scala 97:16]
  assign O_t0b = n274_O_t0b; // @[Top.scala 96:7]
  assign O_t1b = n274_O_t1b; // @[Top.scala 96:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n274_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 95:19]
  assign n274_I0 = I; // @[Top.scala 93:13]
  assign n274_I1 = 8'h2; // @[Top.scala 94:13]
endmodule
module MapS_29(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  output [31:0] O_0_t0b,
  output [7:0]  O_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[MapS.scala 9:22]
  Module_4 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_t0b = fst_op_O_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b = fst_op_O_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
endmodule
module MapS_30(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  output [31:0] O_0_0_t0b,
  output [7:0]  O_0_0_t1b
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[MapS.scala 9:22]
  MapS_29 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
endmodule
module ReduceS_1(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0
);
  wire [31:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t0b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_I_t1b; // @[ReduceS.scala 20:43]
  wire [31:0] AddNoValid_2_O; // @[ReduceS.scala 20:43]
  reg [31:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [31:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [31:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [31:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg [31:0] _T_4; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_5;
  reg  _T_6; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_6;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  AddNoValid AddNoValid_2 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_2_I_t0b),
    .I_t1b(AddNoValid_2_I_t1b),
    .O(AddNoValid_2_O)
  );
  assign valid_down = _T_6; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = AddNoValid_2_O; // @[ReduceS.scala 31:18]
  assign AddNoValid_1_I_t1b = _T_4; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_2_I_t1b = _T_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    _T_4 <= I_3;
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= valid_up;
    end
    _T_6 <= _T_5;
  end
endmodule
module MapS_38(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0,
  input  [31:0] I_0_1,
  input  [31:0] I_0_2,
  input  [31:0] I_0_3,
  output [31:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_3; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0; // @[MapS.scala 9:22]
  ReduceS_1 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .I_3(fst_op_I_3),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_3 = I_0_3; // @[MapS.scala 16:12]
endmodule
module AtomTuple_15(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_t0b,
  input  [31:0] I0_t1b_t0b,
  input  [31:0] I0_t1b_t1b,
  input  [31:0] I1_t0b,
  input  [31:0] I1_t1b_t0b,
  input  [31:0] I1_t1b_t1b,
  output [31:0] O_t0b_t0b,
  output [31:0] O_t0b_t1b_t0b,
  output [31:0] O_t0b_t1b_t1b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b_t0b,
  output [31:0] O_t1b_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b_t0b = I0_t0b; // @[Tuple.scala 49:9]
  assign O_t0b_t1b_t0b = I0_t1b_t0b; // @[Tuple.scala 49:9]
  assign O_t0b_t1b_t1b = I0_t1b_t1b; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t0b = I1_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t1b = I1_t1b_t1b; // @[Tuple.scala 50:9]
endmodule
module Map2S_33(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_t0b,
  input  [31:0] I0_0_t1b_t0b,
  input  [31:0] I0_0_t1b_t1b,
  input  [31:0] I1_0_t0b,
  input  [31:0] I1_0_t1b_t0b,
  input  [31:0] I1_0_t1b_t1b,
  output [31:0] O_0_t0b_t0b,
  output [31:0] O_0_t0b_t1b_t0b,
  output [31:0] O_0_t0b_t1b_t1b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  AtomTuple_15 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_t0b(fst_op_I0_t0b),
    .I0_t1b_t0b(fst_op_I0_t1b_t0b),
    .I0_t1b_t1b(fst_op_I0_t1b_t1b),
    .I1_t0b(fst_op_I1_t0b),
    .I1_t1b_t0b(fst_op_I1_t1b_t0b),
    .I1_t1b_t1b(fst_op_I1_t1b_t1b),
    .O_t0b_t0b(fst_op_O_t0b_t0b),
    .O_t0b_t1b_t0b(fst_op_O_t0b_t1b_t0b),
    .O_t0b_t1b_t1b(fst_op_O_t0b_t1b_t1b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b_t0b(fst_op_O_t1b_t1b_t0b),
    .O_t1b_t1b_t1b(fst_op_O_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b_t0b = fst_op_O_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t0b_t1b_t0b = fst_op_O_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t0b_t1b_t1b = fst_op_O_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t0b = fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t1b = fst_op_O_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_t0b = I0_0_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_t1b_t0b = I0_0_t1b_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_t1b_t1b = I0_0_t1b_t1b; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b = I1_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t0b = I1_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t1b = I1_0_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module Map2S_34(
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_t0b,
  input  [31:0] I0_0_0_t1b_t0b,
  input  [31:0] I0_0_0_t1b_t1b,
  input  [31:0] I1_0_0_t0b,
  input  [31:0] I1_0_0_t1b_t0b,
  input  [31:0] I1_0_0_t1b_t1b,
  output [31:0] O_0_0_t0b_t0b,
  output [31:0] O_0_0_t0b_t1b_t0b,
  output [31:0] O_0_0_t0b_t1b_t1b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  Map2S_33 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_t0b(fst_op_I0_0_t0b),
    .I0_0_t1b_t0b(fst_op_I0_0_t1b_t0b),
    .I0_0_t1b_t1b(fst_op_I0_0_t1b_t1b),
    .I1_0_t0b(fst_op_I1_0_t0b),
    .I1_0_t1b_t0b(fst_op_I1_0_t1b_t0b),
    .I1_0_t1b_t1b(fst_op_I1_0_t1b_t1b),
    .O_0_t0b_t0b(fst_op_O_0_t0b_t0b),
    .O_0_t0b_t1b_t0b(fst_op_O_0_t0b_t1b_t0b),
    .O_0_t0b_t1b_t1b(fst_op_O_0_t0b_t1b_t1b),
    .O_0_t1b_t0b(fst_op_O_0_t1b_t0b),
    .O_0_t1b_t1b_t0b(fst_op_O_0_t1b_t1b_t0b),
    .O_0_t1b_t1b_t1b(fst_op_O_0_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b_t0b = fst_op_O_0_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t0b_t1b_t0b = fst_op_O_0_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t0b_t1b_t1b = fst_op_O_0_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b = fst_op_O_0_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t0b = fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t1b = fst_op_O_0_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_t0b = I0_0_0_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_t1b_t0b = I0_0_0_t1b_t0b; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_t1b_t1b = I0_0_0_t1b_t1b; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_t0b = I1_0_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t0b = I1_0_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t1b = I1_0_0_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module AtomTuple_16(
  input         valid_up,
  output        valid_down,
  input         I0,
  input  [31:0] I1_t0b_t0b,
  input  [31:0] I1_t0b_t1b_t0b,
  input  [31:0] I1_t0b_t1b_t1b,
  input  [31:0] I1_t1b_t0b,
  input  [31:0] I1_t1b_t1b_t0b,
  input  [31:0] I1_t1b_t1b_t1b,
  output        O_t0b,
  output [31:0] O_t1b_t0b_t0b,
  output [31:0] O_t1b_t0b_t1b_t0b,
  output [31:0] O_t1b_t0b_t1b_t1b,
  output [31:0] O_t1b_t1b_t0b,
  output [31:0] O_t1b_t1b_t1b_t0b,
  output [31:0] O_t1b_t1b_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b_t0b = I1_t0b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t0b_t1b_t0b = I1_t0b_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t0b_t1b_t1b = I1_t0b_t1b_t1b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t0b = I1_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t1b_t0b = I1_t1b_t1b_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b_t1b_t1b = I1_t1b_t1b_t1b; // @[Tuple.scala 50:9]
endmodule
module Map2S_35(
  input         valid_up,
  output        valid_down,
  input         I0_0,
  input  [31:0] I1_0_t0b_t0b,
  input  [31:0] I1_0_t0b_t1b_t0b,
  input  [31:0] I1_0_t0b_t1b_t1b,
  input  [31:0] I1_0_t1b_t0b,
  input  [31:0] I1_0_t1b_t1b_t0b,
  input  [31:0] I1_0_t1b_t1b_t1b,
  output        O_0_t0b,
  output [31:0] O_0_t1b_t0b_t0b,
  output [31:0] O_0_t1b_t0b_t1b_t0b,
  output [31:0] O_0_t1b_t0b_t1b_t1b,
  output [31:0] O_0_t1b_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t1b_t0b,
  output [31:0] O_0_t1b_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire  fst_op_I0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  wire  fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  AtomTuple_16 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1_t0b_t0b(fst_op_I1_t0b_t0b),
    .I1_t0b_t1b_t0b(fst_op_I1_t0b_t1b_t0b),
    .I1_t0b_t1b_t1b(fst_op_I1_t0b_t1b_t1b),
    .I1_t1b_t0b(fst_op_I1_t1b_t0b),
    .I1_t1b_t1b_t0b(fst_op_I1_t1b_t1b_t0b),
    .I1_t1b_t1b_t1b(fst_op_I1_t1b_t1b_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b_t0b(fst_op_O_t1b_t0b_t0b),
    .O_t1b_t0b_t1b_t0b(fst_op_O_t1b_t0b_t1b_t0b),
    .O_t1b_t0b_t1b_t1b(fst_op_O_t1b_t0b_t1b_t1b),
    .O_t1b_t1b_t0b(fst_op_O_t1b_t1b_t0b),
    .O_t1b_t1b_t1b_t0b(fst_op_O_t1b_t1b_t1b_t0b),
    .O_t1b_t1b_t1b_t1b(fst_op_O_t1b_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b_t0b = fst_op_O_t1b_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b_t1b_t0b = fst_op_O_t1b_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t0b_t1b_t1b = fst_op_O_t1b_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t0b = fst_op_O_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t1b_t0b = fst_op_O_t1b_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b_t1b_t1b_t1b = fst_op_O_t1b_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_t0b_t0b = I1_0_t0b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t0b_t1b_t0b = I1_0_t0b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t0b_t1b_t1b = I1_0_t0b_t1b_t1b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t0b = I1_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t1b_t0b = I1_0_t1b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_t1b_t1b_t1b = I1_0_t1b_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module Map2S_36(
  input         valid_up,
  output        valid_down,
  input         I0_0_0,
  input  [31:0] I1_0_0_t0b_t0b,
  input  [31:0] I1_0_0_t0b_t1b_t0b,
  input  [31:0] I1_0_0_t0b_t1b_t1b,
  input  [31:0] I1_0_0_t1b_t0b,
  input  [31:0] I1_0_0_t1b_t1b_t0b,
  input  [31:0] I1_0_0_t1b_t1b_t1b,
  output        O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b_t0b,
  output [31:0] O_0_0_t1b_t0b_t1b_t0b,
  output [31:0] O_0_0_t1b_t0b_t1b_t1b,
  output [31:0] O_0_0_t1b_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b_t1b_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire  fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I1_0_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  wire  fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b_t1b_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b_t1b_t1b; // @[Map2S.scala 9:22]
  Map2S_35 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0_t0b_t0b(fst_op_I1_0_t0b_t0b),
    .I1_0_t0b_t1b_t0b(fst_op_I1_0_t0b_t1b_t0b),
    .I1_0_t0b_t1b_t1b(fst_op_I1_0_t0b_t1b_t1b),
    .I1_0_t1b_t0b(fst_op_I1_0_t1b_t0b),
    .I1_0_t1b_t1b_t0b(fst_op_I1_0_t1b_t1b_t0b),
    .I1_0_t1b_t1b_t1b(fst_op_I1_0_t1b_t1b_t1b),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b_t0b_t0b(fst_op_O_0_t1b_t0b_t0b),
    .O_0_t1b_t0b_t1b_t0b(fst_op_O_0_t1b_t0b_t1b_t0b),
    .O_0_t1b_t0b_t1b_t1b(fst_op_O_0_t1b_t0b_t1b_t1b),
    .O_0_t1b_t1b_t0b(fst_op_O_0_t1b_t1b_t0b),
    .O_0_t1b_t1b_t1b_t0b(fst_op_O_0_t1b_t1b_t1b_t0b),
    .O_0_t1b_t1b_t1b_t1b(fst_op_O_0_t1b_t1b_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b_t0b = fst_op_O_0_t1b_t0b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b_t1b_t0b = fst_op_O_0_t1b_t0b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t0b_t1b_t1b = fst_op_O_0_t1b_t0b_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t0b = fst_op_O_0_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t1b_t0b = fst_op_O_0_t1b_t1b_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b_t1b_t1b_t1b = fst_op_O_0_t1b_t1b_t1b_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_t0b_t0b = I1_0_0_t0b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t0b_t1b_t0b = I1_0_0_t0b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t0b_t1b_t1b = I1_0_0_t0b_t1b_t1b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t0b = I1_0_0_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t1b_t0b = I1_0_0_t1b_t1b_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_t1b_t1b_t1b = I1_0_0_t1b_t1b_t1b; // @[Map2S.scala 18:13]
endmodule
module If(
  input         valid_up,
  output        valid_down,
  input         I_t0b,
  input  [31:0] I_t1b_t0b_t0b,
  input  [31:0] I_t1b_t0b_t1b_t0b,
  input  [31:0] I_t1b_t0b_t1b_t1b,
  input  [31:0] I_t1b_t1b_t0b,
  input  [31:0] I_t1b_t1b_t1b_t0b,
  input  [31:0] I_t1b_t1b_t1b_t1b,
  output [31:0] O_t0b,
  output [31:0] O_t1b_t0b,
  output [31:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Arithmetic.scala 525:14]
  assign O_t0b = I_t0b ? I_t1b_t0b_t0b : I_t1b_t1b_t0b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
  assign O_t1b_t0b = I_t0b ? I_t1b_t0b_t1b_t0b : I_t1b_t1b_t1b_t0b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
  assign O_t1b_t1b = I_t0b ? I_t1b_t0b_t1b_t1b : I_t1b_t1b_t1b_t1b; // @[Arithmetic.scala 523:9 Arithmetic.scala 524:20]
endmodule
module MapS_43(
  input         valid_up,
  output        valid_down,
  input         I_0_t0b,
  input  [31:0] I_0_t1b_t0b_t0b,
  input  [31:0] I_0_t1b_t0b_t1b_t0b,
  input  [31:0] I_0_t1b_t0b_t1b_t1b,
  input  [31:0] I_0_t1b_t1b_t0b,
  input  [31:0] I_0_t1b_t1b_t1b_t0b,
  input  [31:0] I_0_t1b_t1b_t1b_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t0b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_t1b_t1b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_t1b_t1b; // @[MapS.scala 9:22]
  If fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b_t0b_t0b(fst_op_I_t1b_t0b_t0b),
    .I_t1b_t0b_t1b_t0b(fst_op_I_t1b_t0b_t1b_t0b),
    .I_t1b_t0b_t1b_t1b(fst_op_I_t1b_t0b_t1b_t1b),
    .I_t1b_t1b_t0b(fst_op_I_t1b_t1b_t0b),
    .I_t1b_t1b_t1b_t0b(fst_op_I_t1b_t1b_t1b_t0b),
    .I_t1b_t1b_t1b_t1b(fst_op_I_t1b_t1b_t1b_t1b),
    .O_t0b(fst_op_O_t0b),
    .O_t1b_t0b(fst_op_O_t1b_t0b),
    .O_t1b_t1b(fst_op_O_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_t0b = fst_op_O_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b_t0b = fst_op_O_t1b_t0b; // @[MapS.scala 17:8]
  assign O_0_t1b_t1b = fst_op_O_t1b_t1b; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t0b_t0b = I_0_t1b_t0b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t0b_t1b_t0b = I_0_t1b_t0b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t0b_t1b_t1b = I_0_t1b_t0b_t1b_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b_t0b = I_0_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b_t1b_t0b = I_0_t1b_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b_t1b_t1b_t1b = I_0_t1b_t1b_t1b_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_44(
  input         valid_up,
  output        valid_down,
  input         I_0_0_t0b,
  input  [31:0] I_0_0_t1b_t0b_t0b,
  input  [31:0] I_0_0_t1b_t0b_t1b_t0b,
  input  [31:0] I_0_0_t1b_t0b_t1b_t1b,
  input  [31:0] I_0_0_t1b_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b_t1b_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire  fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t0b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t0b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t0b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t1b_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_I_0_t1b_t1b_t1b_t1b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t0b; // @[MapS.scala 9:22]
  wire [31:0] fst_op_O_0_t1b_t1b; // @[MapS.scala 9:22]
  MapS_43 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b_t0b_t0b(fst_op_I_0_t1b_t0b_t0b),
    .I_0_t1b_t0b_t1b_t0b(fst_op_I_0_t1b_t0b_t1b_t0b),
    .I_0_t1b_t0b_t1b_t1b(fst_op_I_0_t1b_t0b_t1b_t1b),
    .I_0_t1b_t1b_t0b(fst_op_I_0_t1b_t1b_t0b),
    .I_0_t1b_t1b_t1b_t0b(fst_op_I_0_t1b_t1b_t1b_t0b),
    .I_0_t1b_t1b_t1b_t1b(fst_op_I_0_t1b_t1b_t1b_t1b),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b_t0b(fst_op_O_0_t1b_t0b),
    .O_0_t1b_t1b(fst_op_O_0_t1b_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b_t0b = fst_op_O_0_t1b_t0b; // @[MapS.scala 17:8]
  assign O_0_0_t1b_t1b = fst_op_O_0_t1b_t1b; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t0b_t0b = I_0_0_t1b_t0b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t0b_t1b_t0b = I_0_0_t1b_t0b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t0b_t1b_t1b = I_0_0_t1b_t0b_t1b_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t1b_t0b = I_0_0_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t1b_t1b_t0b = I_0_0_t1b_t1b_t1b_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b_t1b_t1b_t1b = I_0_0_t1b_t1b_t1b_t1b; // @[MapS.scala 16:12]
endmodule
module Module_6(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0,
  input  [31:0] I0_0_1,
  input  [31:0] I0_0_2,
  input  [31:0] I0_1_0,
  input  [31:0] I0_1_1,
  input  [31:0] I0_1_2,
  input  [31:0] I0_2_0,
  input  [31:0] I0_2_1,
  input  [31:0] I0_2_2,
  input         I1_0_0_t0b,
  input         I1_0_0_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b
);
  wire  n152_valid_up; // @[Top.scala 116:22]
  wire  n152_valid_down; // @[Top.scala 116:22]
  wire  n152_I_0_0_t0b; // @[Top.scala 116:22]
  wire  n152_O_0_0; // @[Top.scala 116:22]
  wire  n430_clock; // @[Top.scala 119:22]
  wire  n430_reset; // @[Top.scala 119:22]
  wire  n430_valid_up; // @[Top.scala 119:22]
  wire  n430_valid_down; // @[Top.scala 119:22]
  wire  n430_I_0_0; // @[Top.scala 119:22]
  wire  n430_O_0_0; // @[Top.scala 119:22]
  wire  n157_valid_up; // @[Top.scala 122:22]
  wire  n157_valid_down; // @[Top.scala 122:22]
  wire  n157_I_0_0_t1b; // @[Top.scala 122:22]
  wire  n157_O_0_0; // @[Top.scala 122:22]
  wire  n360_clock; // @[Top.scala 125:22]
  wire  n360_reset; // @[Top.scala 125:22]
  wire  n360_valid_up; // @[Top.scala 125:22]
  wire  n360_valid_down; // @[Top.scala 125:22]
  wire  n360_I_0_0; // @[Top.scala 125:22]
  wire  n360_O_0_0; // @[Top.scala 125:22]
  wire  n159_valid_up; // @[Top.scala 128:22]
  wire  n159_valid_down; // @[Top.scala 128:22]
  wire [31:0] n159_I_1_0; // @[Top.scala 128:22]
  wire [31:0] n159_I_1_1; // @[Top.scala 128:22]
  wire [31:0] n159_I_1_2; // @[Top.scala 128:22]
  wire [31:0] n159_O_0_0; // @[Top.scala 128:22]
  wire [31:0] n159_O_0_1; // @[Top.scala 128:22]
  wire [31:0] n159_O_0_2; // @[Top.scala 128:22]
  wire  n162_valid_up; // @[Top.scala 131:22]
  wire  n162_valid_down; // @[Top.scala 131:22]
  wire [31:0] n162_I_0_0; // @[Top.scala 131:22]
  wire [31:0] n162_O_0_0; // @[Top.scala 131:22]
  wire  n165_valid_up; // @[Top.scala 134:22]
  wire  n165_valid_down; // @[Top.scala 134:22]
  wire [31:0] n165_I_0_2; // @[Top.scala 134:22]
  wire [31:0] n165_O_0_0; // @[Top.scala 134:22]
  wire  n166_valid_up; // @[Top.scala 137:22]
  wire  n166_valid_down; // @[Top.scala 137:22]
  wire [31:0] n166_I0_0_0; // @[Top.scala 137:22]
  wire [31:0] n166_I1_0_0; // @[Top.scala 137:22]
  wire [31:0] n166_O_0_0_t0b; // @[Top.scala 137:22]
  wire [31:0] n166_O_0_0_t1b; // @[Top.scala 137:22]
  wire  n177_valid_up; // @[Top.scala 141:22]
  wire  n177_valid_down; // @[Top.scala 141:22]
  wire [31:0] n177_I_0_0_t0b; // @[Top.scala 141:22]
  wire [31:0] n177_I_0_0_t1b; // @[Top.scala 141:22]
  wire [31:0] n177_O_0_0; // @[Top.scala 141:22]
  wire  n184_clock; // @[Top.scala 144:22]
  wire  n184_reset; // @[Top.scala 144:22]
  wire  n184_valid_up; // @[Top.scala 144:22]
  wire  n184_valid_down; // @[Top.scala 144:22]
  wire [31:0] n184_I_0_0; // @[Top.scala 144:22]
  wire [31:0] n184_O_0_0_t0b; // @[Top.scala 144:22]
  wire [7:0] n184_O_0_0_t1b; // @[Top.scala 144:22]
  wire  n189_valid_up; // @[Top.scala 147:22]
  wire  n189_valid_down; // @[Top.scala 147:22]
  wire [31:0] n189_I_0_0_t0b; // @[Top.scala 147:22]
  wire [7:0] n189_I_0_0_t1b; // @[Top.scala 147:22]
  wire [31:0] n189_O_0_0; // @[Top.scala 147:22]
  wire  n192_valid_up; // @[Top.scala 150:22]
  wire  n192_valid_down; // @[Top.scala 150:22]
  wire [31:0] n192_I_0_1; // @[Top.scala 150:22]
  wire [31:0] n192_O_0_0; // @[Top.scala 150:22]
  wire  n193_valid_up; // @[Top.scala 153:22]
  wire  n193_valid_down; // @[Top.scala 153:22]
  wire [31:0] n193_I_0_0; // @[Top.scala 153:22]
  wire [31:0] n193_I_0_1; // @[Top.scala 153:22]
  wire [31:0] n193_I_0_2; // @[Top.scala 153:22]
  wire [31:0] n193_O_0_0; // @[Top.scala 153:22]
  wire [31:0] n193_O_0_1; // @[Top.scala 153:22]
  wire [31:0] n193_O_0_2; // @[Top.scala 153:22]
  wire  n196_valid_up; // @[Top.scala 156:22]
  wire  n196_valid_down; // @[Top.scala 156:22]
  wire [31:0] n196_I_0_1; // @[Top.scala 156:22]
  wire [31:0] n196_O_0_0; // @[Top.scala 156:22]
  wire  n197_valid_up; // @[Top.scala 159:22]
  wire  n197_valid_down; // @[Top.scala 159:22]
  wire [31:0] n197_I_2_0; // @[Top.scala 159:22]
  wire [31:0] n197_I_2_1; // @[Top.scala 159:22]
  wire [31:0] n197_I_2_2; // @[Top.scala 159:22]
  wire [31:0] n197_O_0_0; // @[Top.scala 159:22]
  wire [31:0] n197_O_0_1; // @[Top.scala 159:22]
  wire [31:0] n197_O_0_2; // @[Top.scala 159:22]
  wire  n200_valid_up; // @[Top.scala 162:22]
  wire  n200_valid_down; // @[Top.scala 162:22]
  wire [31:0] n200_I_0_1; // @[Top.scala 162:22]
  wire [31:0] n200_O_0_0; // @[Top.scala 162:22]
  wire  n201_valid_up; // @[Top.scala 165:22]
  wire  n201_valid_down; // @[Top.scala 165:22]
  wire [31:0] n201_I0_0_0; // @[Top.scala 165:22]
  wire [31:0] n201_I1_0_0; // @[Top.scala 165:22]
  wire [31:0] n201_O_0_0_t0b; // @[Top.scala 165:22]
  wire [31:0] n201_O_0_0_t1b; // @[Top.scala 165:22]
  wire  n212_valid_up; // @[Top.scala 169:22]
  wire  n212_valid_down; // @[Top.scala 169:22]
  wire [31:0] n212_I_0_0_t0b; // @[Top.scala 169:22]
  wire [31:0] n212_I_0_0_t1b; // @[Top.scala 169:22]
  wire [31:0] n212_O_0_0; // @[Top.scala 169:22]
  wire  n219_clock; // @[Top.scala 172:22]
  wire  n219_reset; // @[Top.scala 172:22]
  wire  n219_valid_up; // @[Top.scala 172:22]
  wire  n219_valid_down; // @[Top.scala 172:22]
  wire [31:0] n219_I_0_0; // @[Top.scala 172:22]
  wire [31:0] n219_O_0_0_t0b; // @[Top.scala 172:22]
  wire [7:0] n219_O_0_0_t1b; // @[Top.scala 172:22]
  wire  n224_valid_up; // @[Top.scala 175:22]
  wire  n224_valid_down; // @[Top.scala 175:22]
  wire [31:0] n224_I_0_0_t0b; // @[Top.scala 175:22]
  wire [7:0] n224_I_0_0_t1b; // @[Top.scala 175:22]
  wire [31:0] n224_O_0_0; // @[Top.scala 175:22]
  wire  n225_valid_up; // @[Top.scala 178:22]
  wire  n225_valid_down; // @[Top.scala 178:22]
  wire [31:0] n225_I0_0_0; // @[Top.scala 178:22]
  wire [31:0] n225_I1_0_0; // @[Top.scala 178:22]
  wire [31:0] n225_O_0_0_t0b; // @[Top.scala 178:22]
  wire [31:0] n225_O_0_0_t1b; // @[Top.scala 178:22]
  wire  n232_valid_up; // @[Top.scala 182:22]
  wire  n232_valid_down; // @[Top.scala 182:22]
  wire [31:0] n232_I0_0_0; // @[Top.scala 182:22]
  wire [31:0] n232_I1_0_0_t0b; // @[Top.scala 182:22]
  wire [31:0] n232_I1_0_0_t1b; // @[Top.scala 182:22]
  wire [31:0] n232_O_0_0_t0b; // @[Top.scala 182:22]
  wire [31:0] n232_O_0_0_t1b_t0b; // @[Top.scala 182:22]
  wire [31:0] n232_O_0_0_t1b_t1b; // @[Top.scala 182:22]
  wire  n352_clock; // @[Top.scala 186:22]
  wire  n352_reset; // @[Top.scala 186:22]
  wire  n352_valid_up; // @[Top.scala 186:22]
  wire  n352_valid_down; // @[Top.scala 186:22]
  wire [31:0] n352_I_0_0_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_I_0_0_t1b_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_I_0_0_t1b_t1b; // @[Top.scala 186:22]
  wire [31:0] n352_O_0_0_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_O_0_0_t1b_t0b; // @[Top.scala 186:22]
  wire [31:0] n352_O_0_0_t1b_t1b; // @[Top.scala 186:22]
  wire  n344_clock; // @[Top.scala 189:22]
  wire  n344_reset; // @[Top.scala 189:22]
  wire  n344_valid_up; // @[Top.scala 189:22]
  wire  n344_valid_down; // @[Top.scala 189:22]
  wire [31:0] n344_I_0_0; // @[Top.scala 189:22]
  wire [31:0] n344_O_0_0; // @[Top.scala 189:22]
  wire  n239_valid_up; // @[Top.scala 192:22]
  wire  n239_valid_down; // @[Top.scala 192:22]
  wire [31:0] n239_I0_0_0; // @[Top.scala 192:22]
  wire [31:0] n239_I1_0_0; // @[Top.scala 192:22]
  wire [31:0] n239_O_0_0_0; // @[Top.scala 192:22]
  wire [31:0] n239_O_0_0_1; // @[Top.scala 192:22]
  wire  n246_valid_up; // @[Top.scala 196:22]
  wire  n246_valid_down; // @[Top.scala 196:22]
  wire [31:0] n246_I0_0_0_0; // @[Top.scala 196:22]
  wire [31:0] n246_I0_0_0_1; // @[Top.scala 196:22]
  wire [31:0] n246_I1_0_0; // @[Top.scala 196:22]
  wire [31:0] n246_O_0_0_0; // @[Top.scala 196:22]
  wire [31:0] n246_O_0_0_1; // @[Top.scala 196:22]
  wire [31:0] n246_O_0_0_2; // @[Top.scala 196:22]
  wire  n253_valid_up; // @[Top.scala 200:22]
  wire  n253_valid_down; // @[Top.scala 200:22]
  wire [31:0] n253_I0_0_0_0; // @[Top.scala 200:22]
  wire [31:0] n253_I0_0_0_1; // @[Top.scala 200:22]
  wire [31:0] n253_I0_0_0_2; // @[Top.scala 200:22]
  wire [31:0] n253_I1_0_0; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_0; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_1; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_2; // @[Top.scala 200:22]
  wire [31:0] n253_O_0_0_3; // @[Top.scala 200:22]
  wire  n264_valid_up; // @[Top.scala 204:22]
  wire  n264_valid_down; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_0; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_1; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_2; // @[Top.scala 204:22]
  wire [31:0] n264_I_0_0_3; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_0; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_1; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_2; // @[Top.scala 204:22]
  wire [31:0] n264_O_0_3; // @[Top.scala 204:22]
  wire  n269_clock; // @[Top.scala 207:22]
  wire  n269_reset; // @[Top.scala 207:22]
  wire  n269_valid_up; // @[Top.scala 207:22]
  wire  n269_valid_down; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_0; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_1; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_2; // @[Top.scala 207:22]
  wire [31:0] n269_I_0_3; // @[Top.scala 207:22]
  wire [31:0] n269_O_0_0; // @[Top.scala 207:22]
  wire  n276_clock; // @[Top.scala 210:22]
  wire  n276_reset; // @[Top.scala 210:22]
  wire  n276_valid_up; // @[Top.scala 210:22]
  wire  n276_valid_down; // @[Top.scala 210:22]
  wire [31:0] n276_I_0_0; // @[Top.scala 210:22]
  wire [31:0] n276_O_0_0_t0b; // @[Top.scala 210:22]
  wire [7:0] n276_O_0_0_t1b; // @[Top.scala 210:22]
  wire  n281_valid_up; // @[Top.scala 213:22]
  wire  n281_valid_down; // @[Top.scala 213:22]
  wire [31:0] n281_I_0_0_t0b; // @[Top.scala 213:22]
  wire [7:0] n281_I_0_0_t1b; // @[Top.scala 213:22]
  wire [31:0] n281_O_0_0; // @[Top.scala 213:22]
  wire  n284_valid_up; // @[Top.scala 216:22]
  wire  n284_valid_down; // @[Top.scala 216:22]
  wire [31:0] n284_I_0_0; // @[Top.scala 216:22]
  wire [31:0] n284_O_0_0; // @[Top.scala 216:22]
  wire  n287_valid_up; // @[Top.scala 219:22]
  wire  n287_valid_down; // @[Top.scala 219:22]
  wire [31:0] n287_I_0_2; // @[Top.scala 219:22]
  wire [31:0] n287_O_0_0; // @[Top.scala 219:22]
  wire  n288_valid_up; // @[Top.scala 222:22]
  wire  n288_valid_down; // @[Top.scala 222:22]
  wire [31:0] n288_I0_0_0; // @[Top.scala 222:22]
  wire [31:0] n288_I1_0_0; // @[Top.scala 222:22]
  wire [31:0] n288_O_0_0_0; // @[Top.scala 222:22]
  wire [31:0] n288_O_0_0_1; // @[Top.scala 222:22]
  wire  n297_valid_up; // @[Top.scala 226:22]
  wire  n297_valid_down; // @[Top.scala 226:22]
  wire [31:0] n297_I_0_0; // @[Top.scala 226:22]
  wire [31:0] n297_O_0_0; // @[Top.scala 226:22]
  wire  n298_valid_up; // @[Top.scala 229:22]
  wire  n298_valid_down; // @[Top.scala 229:22]
  wire [31:0] n298_I0_0_0_0; // @[Top.scala 229:22]
  wire [31:0] n298_I0_0_0_1; // @[Top.scala 229:22]
  wire [31:0] n298_I1_0_0; // @[Top.scala 229:22]
  wire [31:0] n298_O_0_0_0; // @[Top.scala 229:22]
  wire [31:0] n298_O_0_0_1; // @[Top.scala 229:22]
  wire [31:0] n298_O_0_0_2; // @[Top.scala 229:22]
  wire  n307_valid_up; // @[Top.scala 233:22]
  wire  n307_valid_down; // @[Top.scala 233:22]
  wire [31:0] n307_I_0_2; // @[Top.scala 233:22]
  wire [31:0] n307_O_0_0; // @[Top.scala 233:22]
  wire  n308_valid_up; // @[Top.scala 236:22]
  wire  n308_valid_down; // @[Top.scala 236:22]
  wire [31:0] n308_I0_0_0_0; // @[Top.scala 236:22]
  wire [31:0] n308_I0_0_0_1; // @[Top.scala 236:22]
  wire [31:0] n308_I0_0_0_2; // @[Top.scala 236:22]
  wire [31:0] n308_I1_0_0; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_0; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_1; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_2; // @[Top.scala 236:22]
  wire [31:0] n308_O_0_0_3; // @[Top.scala 236:22]
  wire  n319_valid_up; // @[Top.scala 240:22]
  wire  n319_valid_down; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_0; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_1; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_2; // @[Top.scala 240:22]
  wire [31:0] n319_I_0_0_3; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_0; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_1; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_2; // @[Top.scala 240:22]
  wire [31:0] n319_O_0_3; // @[Top.scala 240:22]
  wire  n324_clock; // @[Top.scala 243:22]
  wire  n324_reset; // @[Top.scala 243:22]
  wire  n324_valid_up; // @[Top.scala 243:22]
  wire  n324_valid_down; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_0; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_1; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_2; // @[Top.scala 243:22]
  wire [31:0] n324_I_0_3; // @[Top.scala 243:22]
  wire [31:0] n324_O_0_0; // @[Top.scala 243:22]
  wire  n331_clock; // @[Top.scala 246:22]
  wire  n331_reset; // @[Top.scala 246:22]
  wire  n331_valid_up; // @[Top.scala 246:22]
  wire  n331_valid_down; // @[Top.scala 246:22]
  wire [31:0] n331_I_0_0; // @[Top.scala 246:22]
  wire [31:0] n331_O_0_0_t0b; // @[Top.scala 246:22]
  wire [7:0] n331_O_0_0_t1b; // @[Top.scala 246:22]
  wire  n336_valid_up; // @[Top.scala 249:22]
  wire  n336_valid_down; // @[Top.scala 249:22]
  wire [31:0] n336_I_0_0_t0b; // @[Top.scala 249:22]
  wire [7:0] n336_I_0_0_t1b; // @[Top.scala 249:22]
  wire [31:0] n336_O_0_0; // @[Top.scala 249:22]
  wire  n337_valid_up; // @[Top.scala 252:22]
  wire  n337_valid_down; // @[Top.scala 252:22]
  wire [31:0] n337_I0_0_0; // @[Top.scala 252:22]
  wire [31:0] n337_I1_0_0; // @[Top.scala 252:22]
  wire [31:0] n337_O_0_0_t0b; // @[Top.scala 252:22]
  wire [31:0] n337_O_0_0_t1b; // @[Top.scala 252:22]
  wire  n345_valid_up; // @[Top.scala 256:22]
  wire  n345_valid_down; // @[Top.scala 256:22]
  wire [31:0] n345_I0_0_0; // @[Top.scala 256:22]
  wire [31:0] n345_I1_0_0_t0b; // @[Top.scala 256:22]
  wire [31:0] n345_I1_0_0_t1b; // @[Top.scala 256:22]
  wire [31:0] n345_O_0_0_t0b; // @[Top.scala 256:22]
  wire [31:0] n345_O_0_0_t1b_t0b; // @[Top.scala 256:22]
  wire [31:0] n345_O_0_0_t1b_t1b; // @[Top.scala 256:22]
  wire  n353_valid_up; // @[Top.scala 260:22]
  wire  n353_valid_down; // @[Top.scala 260:22]
  wire [31:0] n353_I0_0_0_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I0_0_0_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I0_0_0_t1b_t1b; // @[Top.scala 260:22]
  wire [31:0] n353_I1_0_0_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I1_0_0_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_I1_0_0_t1b_t1b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t0b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t0b_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t0b_t1b_t1b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t1b_t1b_t0b; // @[Top.scala 260:22]
  wire [31:0] n353_O_0_0_t1b_t1b_t1b; // @[Top.scala 260:22]
  wire  n361_valid_up; // @[Top.scala 264:22]
  wire  n361_valid_down; // @[Top.scala 264:22]
  wire  n361_I0_0_0; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t0b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t0b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t0b_t1b_t1b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t1b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_I1_0_0_t1b_t1b_t1b; // @[Top.scala 264:22]
  wire  n361_O_0_0_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t0b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 264:22]
  wire [31:0] n361_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 264:22]
  wire  n372_valid_up; // @[Top.scala 268:22]
  wire  n372_valid_down; // @[Top.scala 268:22]
  wire  n372_I_0_0_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t0b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_I_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 268:22]
  wire [31:0] n372_O_0_0_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_O_0_0_t1b_t0b; // @[Top.scala 268:22]
  wire [31:0] n372_O_0_0_t1b_t1b; // @[Top.scala 268:22]
  wire  n410_clock; // @[Top.scala 271:22]
  wire  n410_reset; // @[Top.scala 271:22]
  wire  n410_valid_up; // @[Top.scala 271:22]
  wire  n410_valid_down; // @[Top.scala 271:22]
  wire  n410_I_0_0; // @[Top.scala 271:22]
  wire  n410_O_0_0; // @[Top.scala 271:22]
  wire  n373_clock; // @[Top.scala 274:22]
  wire  n373_reset; // @[Top.scala 274:22]
  wire  n373_valid_up; // @[Top.scala 274:22]
  wire  n373_valid_down; // @[Top.scala 274:22]
  wire [31:0] n373_I_0_0; // @[Top.scala 274:22]
  wire [31:0] n373_O_0_0; // @[Top.scala 274:22]
  wire  n374_valid_up; // @[Top.scala 277:22]
  wire  n374_valid_down; // @[Top.scala 277:22]
  wire [31:0] n374_I0_0_0; // @[Top.scala 277:22]
  wire [31:0] n374_I1_0_0; // @[Top.scala 277:22]
  wire [31:0] n374_O_0_0_t0b; // @[Top.scala 277:22]
  wire [31:0] n374_O_0_0_t1b; // @[Top.scala 277:22]
  wire  n381_valid_up; // @[Top.scala 281:22]
  wire  n381_valid_down; // @[Top.scala 281:22]
  wire [31:0] n381_I0_0_0; // @[Top.scala 281:22]
  wire [31:0] n381_I1_0_0_t0b; // @[Top.scala 281:22]
  wire [31:0] n381_I1_0_0_t1b; // @[Top.scala 281:22]
  wire [31:0] n381_O_0_0_t0b; // @[Top.scala 281:22]
  wire [31:0] n381_O_0_0_t1b_t0b; // @[Top.scala 281:22]
  wire [31:0] n381_O_0_0_t1b_t1b; // @[Top.scala 281:22]
  wire  n388_valid_up; // @[Top.scala 285:22]
  wire  n388_valid_down; // @[Top.scala 285:22]
  wire [31:0] n388_I0_0_0; // @[Top.scala 285:22]
  wire [31:0] n388_I1_0_0; // @[Top.scala 285:22]
  wire [31:0] n388_O_0_0_t0b; // @[Top.scala 285:22]
  wire [31:0] n388_O_0_0_t1b; // @[Top.scala 285:22]
  wire  n395_valid_up; // @[Top.scala 289:22]
  wire  n395_valid_down; // @[Top.scala 289:22]
  wire [31:0] n395_I0_0_0; // @[Top.scala 289:22]
  wire [31:0] n395_I1_0_0_t0b; // @[Top.scala 289:22]
  wire [31:0] n395_I1_0_0_t1b; // @[Top.scala 289:22]
  wire [31:0] n395_O_0_0_t0b; // @[Top.scala 289:22]
  wire [31:0] n395_O_0_0_t1b_t0b; // @[Top.scala 289:22]
  wire [31:0] n395_O_0_0_t1b_t1b; // @[Top.scala 289:22]
  wire  n402_clock; // @[Top.scala 293:22]
  wire  n402_reset; // @[Top.scala 293:22]
  wire  n402_valid_up; // @[Top.scala 293:22]
  wire  n402_valid_down; // @[Top.scala 293:22]
  wire [31:0] n402_I_0_0_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_I_0_0_t1b_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_I_0_0_t1b_t1b; // @[Top.scala 293:22]
  wire [31:0] n402_O_0_0_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_O_0_0_t1b_t0b; // @[Top.scala 293:22]
  wire [31:0] n402_O_0_0_t1b_t1b; // @[Top.scala 293:22]
  wire  n403_valid_up; // @[Top.scala 296:22]
  wire  n403_valid_down; // @[Top.scala 296:22]
  wire [31:0] n403_I0_0_0_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I0_0_0_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I0_0_0_t1b_t1b; // @[Top.scala 296:22]
  wire [31:0] n403_I1_0_0_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I1_0_0_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_I1_0_0_t1b_t1b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t0b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t0b_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t0b_t1b_t1b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t1b_t1b_t0b; // @[Top.scala 296:22]
  wire [31:0] n403_O_0_0_t1b_t1b_t1b; // @[Top.scala 296:22]
  wire  n411_valid_up; // @[Top.scala 300:22]
  wire  n411_valid_down; // @[Top.scala 300:22]
  wire  n411_I0_0_0; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t0b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t0b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t0b_t1b_t1b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t1b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_I1_0_0_t1b_t1b_t1b; // @[Top.scala 300:22]
  wire  n411_O_0_0_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t0b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 300:22]
  wire [31:0] n411_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 300:22]
  wire  n422_valid_up; // @[Top.scala 304:22]
  wire  n422_valid_down; // @[Top.scala 304:22]
  wire  n422_I_0_0_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t0b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_I_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 304:22]
  wire [31:0] n422_O_0_0_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_O_0_0_t1b_t0b; // @[Top.scala 304:22]
  wire [31:0] n422_O_0_0_t1b_t1b; // @[Top.scala 304:22]
  wire  n423_valid_up; // @[Top.scala 307:22]
  wire  n423_valid_down; // @[Top.scala 307:22]
  wire [31:0] n423_I0_0_0_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I0_0_0_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I0_0_0_t1b_t1b; // @[Top.scala 307:22]
  wire [31:0] n423_I1_0_0_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I1_0_0_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_I1_0_0_t1b_t1b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t0b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t0b_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t0b_t1b_t1b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t1b_t1b_t0b; // @[Top.scala 307:22]
  wire [31:0] n423_O_0_0_t1b_t1b_t1b; // @[Top.scala 307:22]
  wire  n431_valid_up; // @[Top.scala 311:22]
  wire  n431_valid_down; // @[Top.scala 311:22]
  wire  n431_I0_0_0; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t0b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t0b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t0b_t1b_t1b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t1b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_I1_0_0_t1b_t1b_t1b; // @[Top.scala 311:22]
  wire  n431_O_0_0_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t0b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 311:22]
  wire [31:0] n431_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 311:22]
  wire  n442_valid_up; // @[Top.scala 315:22]
  wire  n442_valid_down; // @[Top.scala 315:22]
  wire  n442_I_0_0_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t0b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_I_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 315:22]
  wire [31:0] n442_O_0_0_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_O_0_0_t1b_t0b; // @[Top.scala 315:22]
  wire [31:0] n442_O_0_0_t1b_t1b; // @[Top.scala 315:22]
  MapS_7 n152 ( // @[Top.scala 116:22]
    .valid_up(n152_valid_up),
    .valid_down(n152_valid_down),
    .I_0_0_t0b(n152_I_0_0_t0b),
    .O_0_0(n152_O_0_0)
  );
  FIFO_2 n430 ( // @[Top.scala 119:22]
    .clock(n430_clock),
    .reset(n430_reset),
    .valid_up(n430_valid_up),
    .valid_down(n430_valid_down),
    .I_0_0(n430_I_0_0),
    .O_0_0(n430_O_0_0)
  );
  MapS_9 n157 ( // @[Top.scala 122:22]
    .valid_up(n157_valid_up),
    .valid_down(n157_valid_down),
    .I_0_0_t1b(n157_I_0_0_t1b),
    .O_0_0(n157_O_0_0)
  );
  FIFO_2 n360 ( // @[Top.scala 125:22]
    .clock(n360_clock),
    .reset(n360_reset),
    .valid_up(n360_valid_up),
    .valid_down(n360_valid_down),
    .I_0_0(n360_I_0_0),
    .O_0_0(n360_O_0_0)
  );
  DownS n159 ( // @[Top.scala 128:22]
    .valid_up(n159_valid_up),
    .valid_down(n159_valid_down),
    .I_1_0(n159_I_1_0),
    .I_1_1(n159_I_1_1),
    .I_1_2(n159_I_1_2),
    .O_0_0(n159_O_0_0),
    .O_0_1(n159_O_0_1),
    .O_0_2(n159_O_0_2)
  );
  MapS_10 n162 ( // @[Top.scala 131:22]
    .valid_up(n162_valid_up),
    .valid_down(n162_valid_down),
    .I_0_0(n162_I_0_0),
    .O_0_0(n162_O_0_0)
  );
  MapS_11 n165 ( // @[Top.scala 134:22]
    .valid_up(n165_valid_up),
    .valid_down(n165_valid_down),
    .I_0_2(n165_I_0_2),
    .O_0_0(n165_O_0_0)
  );
  Map2S_10 n166 ( // @[Top.scala 137:22]
    .valid_up(n166_valid_up),
    .valid_down(n166_valid_down),
    .I0_0_0(n166_I0_0_0),
    .I1_0_0(n166_I1_0_0),
    .O_0_0_t0b(n166_O_0_0_t0b),
    .O_0_0_t1b(n166_O_0_0_t1b)
  );
  MapS_13 n177 ( // @[Top.scala 141:22]
    .valid_up(n177_valid_up),
    .valid_down(n177_valid_down),
    .I_0_0_t0b(n177_I_0_0_t0b),
    .I_0_0_t1b(n177_I_0_0_t1b),
    .O_0_0(n177_O_0_0)
  );
  MapS_15 n184 ( // @[Top.scala 144:22]
    .clock(n184_clock),
    .reset(n184_reset),
    .valid_up(n184_valid_up),
    .valid_down(n184_valid_down),
    .I_0_0(n184_I_0_0),
    .O_0_0_t0b(n184_O_0_0_t0b),
    .O_0_0_t1b(n184_O_0_0_t1b)
  );
  MapS_17 n189 ( // @[Top.scala 147:22]
    .valid_up(n189_valid_up),
    .valid_down(n189_valid_down),
    .I_0_0_t0b(n189_I_0_0_t0b),
    .I_0_0_t1b(n189_I_0_0_t1b),
    .O_0_0(n189_O_0_0)
  );
  MapS_18 n192 ( // @[Top.scala 150:22]
    .valid_up(n192_valid_up),
    .valid_down(n192_valid_down),
    .I_0_1(n192_I_0_1),
    .O_0_0(n192_O_0_0)
  );
  DownS_4 n193 ( // @[Top.scala 153:22]
    .valid_up(n193_valid_up),
    .valid_down(n193_valid_down),
    .I_0_0(n193_I_0_0),
    .I_0_1(n193_I_0_1),
    .I_0_2(n193_I_0_2),
    .O_0_0(n193_O_0_0),
    .O_0_1(n193_O_0_1),
    .O_0_2(n193_O_0_2)
  );
  MapS_18 n196 ( // @[Top.scala 156:22]
    .valid_up(n196_valid_up),
    .valid_down(n196_valid_down),
    .I_0_1(n196_I_0_1),
    .O_0_0(n196_O_0_0)
  );
  DownS_6 n197 ( // @[Top.scala 159:22]
    .valid_up(n197_valid_up),
    .valid_down(n197_valid_down),
    .I_2_0(n197_I_2_0),
    .I_2_1(n197_I_2_1),
    .I_2_2(n197_I_2_2),
    .O_0_0(n197_O_0_0),
    .O_0_1(n197_O_0_1),
    .O_0_2(n197_O_0_2)
  );
  MapS_18 n200 ( // @[Top.scala 162:22]
    .valid_up(n200_valid_up),
    .valid_down(n200_valid_down),
    .I_0_1(n200_I_0_1),
    .O_0_0(n200_O_0_0)
  );
  Map2S_10 n201 ( // @[Top.scala 165:22]
    .valid_up(n201_valid_up),
    .valid_down(n201_valid_down),
    .I0_0_0(n201_I0_0_0),
    .I1_0_0(n201_I1_0_0),
    .O_0_0_t0b(n201_O_0_0_t0b),
    .O_0_0_t1b(n201_O_0_0_t1b)
  );
  MapS_13 n212 ( // @[Top.scala 169:22]
    .valid_up(n212_valid_up),
    .valid_down(n212_valid_down),
    .I_0_0_t0b(n212_I_0_0_t0b),
    .I_0_0_t1b(n212_I_0_0_t1b),
    .O_0_0(n212_O_0_0)
  );
  MapS_15 n219 ( // @[Top.scala 172:22]
    .clock(n219_clock),
    .reset(n219_reset),
    .valid_up(n219_valid_up),
    .valid_down(n219_valid_down),
    .I_0_0(n219_I_0_0),
    .O_0_0_t0b(n219_O_0_0_t0b),
    .O_0_0_t1b(n219_O_0_0_t1b)
  );
  MapS_17 n224 ( // @[Top.scala 175:22]
    .valid_up(n224_valid_up),
    .valid_down(n224_valid_down),
    .I_0_0_t0b(n224_I_0_0_t0b),
    .I_0_0_t1b(n224_I_0_0_t1b),
    .O_0_0(n224_O_0_0)
  );
  Map2S_10 n225 ( // @[Top.scala 178:22]
    .valid_up(n225_valid_up),
    .valid_down(n225_valid_down),
    .I0_0_0(n225_I0_0_0),
    .I1_0_0(n225_I1_0_0),
    .O_0_0_t0b(n225_O_0_0_t0b),
    .O_0_0_t1b(n225_O_0_0_t1b)
  );
  Map2S_16 n232 ( // @[Top.scala 182:22]
    .valid_up(n232_valid_up),
    .valid_down(n232_valid_down),
    .I0_0_0(n232_I0_0_0),
    .I1_0_0_t0b(n232_I1_0_0_t0b),
    .I1_0_0_t1b(n232_I1_0_0_t1b),
    .O_0_0_t0b(n232_O_0_0_t0b),
    .O_0_0_t1b_t0b(n232_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n232_O_0_0_t1b_t1b)
  );
  FIFO_4 n352 ( // @[Top.scala 186:22]
    .clock(n352_clock),
    .reset(n352_reset),
    .valid_up(n352_valid_up),
    .valid_down(n352_valid_down),
    .I_0_0_t0b(n352_I_0_0_t0b),
    .I_0_0_t1b_t0b(n352_I_0_0_t1b_t0b),
    .I_0_0_t1b_t1b(n352_I_0_0_t1b_t1b),
    .O_0_0_t0b(n352_O_0_0_t0b),
    .O_0_0_t1b_t0b(n352_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n352_O_0_0_t1b_t1b)
  );
  FIFO_5 n344 ( // @[Top.scala 189:22]
    .clock(n344_clock),
    .reset(n344_reset),
    .valid_up(n344_valid_up),
    .valid_down(n344_valid_down),
    .I_0_0(n344_I_0_0),
    .O_0_0(n344_O_0_0)
  );
  Map2S_18 n239 ( // @[Top.scala 192:22]
    .valid_up(n239_valid_up),
    .valid_down(n239_valid_down),
    .I0_0_0(n239_I0_0_0),
    .I1_0_0(n239_I1_0_0),
    .O_0_0_0(n239_O_0_0_0),
    .O_0_0_1(n239_O_0_0_1)
  );
  Map2S_20 n246 ( // @[Top.scala 196:22]
    .valid_up(n246_valid_up),
    .valid_down(n246_valid_down),
    .I0_0_0_0(n246_I0_0_0_0),
    .I0_0_0_1(n246_I0_0_0_1),
    .I1_0_0(n246_I1_0_0),
    .O_0_0_0(n246_O_0_0_0),
    .O_0_0_1(n246_O_0_0_1),
    .O_0_0_2(n246_O_0_0_2)
  );
  Map2S_22 n253 ( // @[Top.scala 200:22]
    .valid_up(n253_valid_up),
    .valid_down(n253_valid_down),
    .I0_0_0_0(n253_I0_0_0_0),
    .I0_0_0_1(n253_I0_0_0_1),
    .I0_0_0_2(n253_I0_0_0_2),
    .I1_0_0(n253_I1_0_0),
    .O_0_0_0(n253_O_0_0_0),
    .O_0_0_1(n253_O_0_0_1),
    .O_0_0_2(n253_O_0_0_2),
    .O_0_0_3(n253_O_0_0_3)
  );
  MapS_27 n264 ( // @[Top.scala 204:22]
    .valid_up(n264_valid_up),
    .valid_down(n264_valid_down),
    .I_0_0_0(n264_I_0_0_0),
    .I_0_0_1(n264_I_0_0_1),
    .I_0_0_2(n264_I_0_0_2),
    .I_0_0_3(n264_I_0_0_3),
    .O_0_0(n264_O_0_0),
    .O_0_1(n264_O_0_1),
    .O_0_2(n264_O_0_2),
    .O_0_3(n264_O_0_3)
  );
  MapS_28 n269 ( // @[Top.scala 207:22]
    .clock(n269_clock),
    .reset(n269_reset),
    .valid_up(n269_valid_up),
    .valid_down(n269_valid_down),
    .I_0_0(n269_I_0_0),
    .I_0_1(n269_I_0_1),
    .I_0_2(n269_I_0_2),
    .I_0_3(n269_I_0_3),
    .O_0_0(n269_O_0_0)
  );
  MapS_30 n276 ( // @[Top.scala 210:22]
    .clock(n276_clock),
    .reset(n276_reset),
    .valid_up(n276_valid_up),
    .valid_down(n276_valid_down),
    .I_0_0(n276_I_0_0),
    .O_0_0_t0b(n276_O_0_0_t0b),
    .O_0_0_t1b(n276_O_0_0_t1b)
  );
  MapS_17 n281 ( // @[Top.scala 213:22]
    .valid_up(n281_valid_up),
    .valid_down(n281_valid_down),
    .I_0_0_t0b(n281_I_0_0_t0b),
    .I_0_0_t1b(n281_I_0_0_t1b),
    .O_0_0(n281_O_0_0)
  );
  MapS_10 n284 ( // @[Top.scala 216:22]
    .valid_up(n284_valid_up),
    .valid_down(n284_valid_down),
    .I_0_0(n284_I_0_0),
    .O_0_0(n284_O_0_0)
  );
  MapS_11 n287 ( // @[Top.scala 219:22]
    .valid_up(n287_valid_up),
    .valid_down(n287_valid_down),
    .I_0_2(n287_I_0_2),
    .O_0_0(n287_O_0_0)
  );
  Map2S_18 n288 ( // @[Top.scala 222:22]
    .valid_up(n288_valid_up),
    .valid_down(n288_valid_down),
    .I0_0_0(n288_I0_0_0),
    .I1_0_0(n288_I1_0_0),
    .O_0_0_0(n288_O_0_0_0),
    .O_0_0_1(n288_O_0_0_1)
  );
  MapS_10 n297 ( // @[Top.scala 226:22]
    .valid_up(n297_valid_up),
    .valid_down(n297_valid_down),
    .I_0_0(n297_I_0_0),
    .O_0_0(n297_O_0_0)
  );
  Map2S_20 n298 ( // @[Top.scala 229:22]
    .valid_up(n298_valid_up),
    .valid_down(n298_valid_down),
    .I0_0_0_0(n298_I0_0_0_0),
    .I0_0_0_1(n298_I0_0_0_1),
    .I1_0_0(n298_I1_0_0),
    .O_0_0_0(n298_O_0_0_0),
    .O_0_0_1(n298_O_0_0_1),
    .O_0_0_2(n298_O_0_0_2)
  );
  MapS_11 n307 ( // @[Top.scala 233:22]
    .valid_up(n307_valid_up),
    .valid_down(n307_valid_down),
    .I_0_2(n307_I_0_2),
    .O_0_0(n307_O_0_0)
  );
  Map2S_22 n308 ( // @[Top.scala 236:22]
    .valid_up(n308_valid_up),
    .valid_down(n308_valid_down),
    .I0_0_0_0(n308_I0_0_0_0),
    .I0_0_0_1(n308_I0_0_0_1),
    .I0_0_0_2(n308_I0_0_0_2),
    .I1_0_0(n308_I1_0_0),
    .O_0_0_0(n308_O_0_0_0),
    .O_0_0_1(n308_O_0_0_1),
    .O_0_0_2(n308_O_0_0_2),
    .O_0_0_3(n308_O_0_0_3)
  );
  MapS_27 n319 ( // @[Top.scala 240:22]
    .valid_up(n319_valid_up),
    .valid_down(n319_valid_down),
    .I_0_0_0(n319_I_0_0_0),
    .I_0_0_1(n319_I_0_0_1),
    .I_0_0_2(n319_I_0_0_2),
    .I_0_0_3(n319_I_0_0_3),
    .O_0_0(n319_O_0_0),
    .O_0_1(n319_O_0_1),
    .O_0_2(n319_O_0_2),
    .O_0_3(n319_O_0_3)
  );
  MapS_38 n324 ( // @[Top.scala 243:22]
    .clock(n324_clock),
    .reset(n324_reset),
    .valid_up(n324_valid_up),
    .valid_down(n324_valid_down),
    .I_0_0(n324_I_0_0),
    .I_0_1(n324_I_0_1),
    .I_0_2(n324_I_0_2),
    .I_0_3(n324_I_0_3),
    .O_0_0(n324_O_0_0)
  );
  MapS_30 n331 ( // @[Top.scala 246:22]
    .clock(n331_clock),
    .reset(n331_reset),
    .valid_up(n331_valid_up),
    .valid_down(n331_valid_down),
    .I_0_0(n331_I_0_0),
    .O_0_0_t0b(n331_O_0_0_t0b),
    .O_0_0_t1b(n331_O_0_0_t1b)
  );
  MapS_17 n336 ( // @[Top.scala 249:22]
    .valid_up(n336_valid_up),
    .valid_down(n336_valid_down),
    .I_0_0_t0b(n336_I_0_0_t0b),
    .I_0_0_t1b(n336_I_0_0_t1b),
    .O_0_0(n336_O_0_0)
  );
  Map2S_10 n337 ( // @[Top.scala 252:22]
    .valid_up(n337_valid_up),
    .valid_down(n337_valid_down),
    .I0_0_0(n337_I0_0_0),
    .I1_0_0(n337_I1_0_0),
    .O_0_0_t0b(n337_O_0_0_t0b),
    .O_0_0_t1b(n337_O_0_0_t1b)
  );
  Map2S_16 n345 ( // @[Top.scala 256:22]
    .valid_up(n345_valid_up),
    .valid_down(n345_valid_down),
    .I0_0_0(n345_I0_0_0),
    .I1_0_0_t0b(n345_I1_0_0_t0b),
    .I1_0_0_t1b(n345_I1_0_0_t1b),
    .O_0_0_t0b(n345_O_0_0_t0b),
    .O_0_0_t1b_t0b(n345_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n345_O_0_0_t1b_t1b)
  );
  Map2S_34 n353 ( // @[Top.scala 260:22]
    .valid_up(n353_valid_up),
    .valid_down(n353_valid_down),
    .I0_0_0_t0b(n353_I0_0_0_t0b),
    .I0_0_0_t1b_t0b(n353_I0_0_0_t1b_t0b),
    .I0_0_0_t1b_t1b(n353_I0_0_0_t1b_t1b),
    .I1_0_0_t0b(n353_I1_0_0_t0b),
    .I1_0_0_t1b_t0b(n353_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b(n353_I1_0_0_t1b_t1b),
    .O_0_0_t0b_t0b(n353_O_0_0_t0b_t0b),
    .O_0_0_t0b_t1b_t0b(n353_O_0_0_t0b_t1b_t0b),
    .O_0_0_t0b_t1b_t1b(n353_O_0_0_t0b_t1b_t1b),
    .O_0_0_t1b_t0b(n353_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b_t0b(n353_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b(n353_O_0_0_t1b_t1b_t1b)
  );
  Map2S_36 n361 ( // @[Top.scala 264:22]
    .valid_up(n361_valid_up),
    .valid_down(n361_valid_down),
    .I0_0_0(n361_I0_0_0),
    .I1_0_0_t0b_t0b(n361_I1_0_0_t0b_t0b),
    .I1_0_0_t0b_t1b_t0b(n361_I1_0_0_t0b_t1b_t0b),
    .I1_0_0_t0b_t1b_t1b(n361_I1_0_0_t0b_t1b_t1b),
    .I1_0_0_t1b_t0b(n361_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b_t0b(n361_I1_0_0_t1b_t1b_t0b),
    .I1_0_0_t1b_t1b_t1b(n361_I1_0_0_t1b_t1b_t1b),
    .O_0_0_t0b(n361_O_0_0_t0b),
    .O_0_0_t1b_t0b_t0b(n361_O_0_0_t1b_t0b_t0b),
    .O_0_0_t1b_t0b_t1b_t0b(n361_O_0_0_t1b_t0b_t1b_t0b),
    .O_0_0_t1b_t0b_t1b_t1b(n361_O_0_0_t1b_t0b_t1b_t1b),
    .O_0_0_t1b_t1b_t0b(n361_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t0b(n361_O_0_0_t1b_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t1b(n361_O_0_0_t1b_t1b_t1b_t1b)
  );
  MapS_44 n372 ( // @[Top.scala 268:22]
    .valid_up(n372_valid_up),
    .valid_down(n372_valid_down),
    .I_0_0_t0b(n372_I_0_0_t0b),
    .I_0_0_t1b_t0b_t0b(n372_I_0_0_t1b_t0b_t0b),
    .I_0_0_t1b_t0b_t1b_t0b(n372_I_0_0_t1b_t0b_t1b_t0b),
    .I_0_0_t1b_t0b_t1b_t1b(n372_I_0_0_t1b_t0b_t1b_t1b),
    .I_0_0_t1b_t1b_t0b(n372_I_0_0_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t0b(n372_I_0_0_t1b_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t1b(n372_I_0_0_t1b_t1b_t1b_t1b),
    .O_0_0_t0b(n372_O_0_0_t0b),
    .O_0_0_t1b_t0b(n372_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n372_O_0_0_t1b_t1b)
  );
  FIFO_2 n410 ( // @[Top.scala 271:22]
    .clock(n410_clock),
    .reset(n410_reset),
    .valid_up(n410_valid_up),
    .valid_down(n410_valid_down),
    .I_0_0(n410_I_0_0),
    .O_0_0(n410_O_0_0)
  );
  FIFO_5 n373 ( // @[Top.scala 274:22]
    .clock(n373_clock),
    .reset(n373_reset),
    .valid_up(n373_valid_up),
    .valid_down(n373_valid_down),
    .I_0_0(n373_I_0_0),
    .O_0_0(n373_O_0_0)
  );
  Map2S_10 n374 ( // @[Top.scala 277:22]
    .valid_up(n374_valid_up),
    .valid_down(n374_valid_down),
    .I0_0_0(n374_I0_0_0),
    .I1_0_0(n374_I1_0_0),
    .O_0_0_t0b(n374_O_0_0_t0b),
    .O_0_0_t1b(n374_O_0_0_t1b)
  );
  Map2S_16 n381 ( // @[Top.scala 281:22]
    .valid_up(n381_valid_up),
    .valid_down(n381_valid_down),
    .I0_0_0(n381_I0_0_0),
    .I1_0_0_t0b(n381_I1_0_0_t0b),
    .I1_0_0_t1b(n381_I1_0_0_t1b),
    .O_0_0_t0b(n381_O_0_0_t0b),
    .O_0_0_t1b_t0b(n381_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n381_O_0_0_t1b_t1b)
  );
  Map2S_10 n388 ( // @[Top.scala 285:22]
    .valid_up(n388_valid_up),
    .valid_down(n388_valid_down),
    .I0_0_0(n388_I0_0_0),
    .I1_0_0(n388_I1_0_0),
    .O_0_0_t0b(n388_O_0_0_t0b),
    .O_0_0_t1b(n388_O_0_0_t1b)
  );
  Map2S_16 n395 ( // @[Top.scala 289:22]
    .valid_up(n395_valid_up),
    .valid_down(n395_valid_down),
    .I0_0_0(n395_I0_0_0),
    .I1_0_0_t0b(n395_I1_0_0_t0b),
    .I1_0_0_t1b(n395_I1_0_0_t1b),
    .O_0_0_t0b(n395_O_0_0_t0b),
    .O_0_0_t1b_t0b(n395_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n395_O_0_0_t1b_t1b)
  );
  FIFO_4 n402 ( // @[Top.scala 293:22]
    .clock(n402_clock),
    .reset(n402_reset),
    .valid_up(n402_valid_up),
    .valid_down(n402_valid_down),
    .I_0_0_t0b(n402_I_0_0_t0b),
    .I_0_0_t1b_t0b(n402_I_0_0_t1b_t0b),
    .I_0_0_t1b_t1b(n402_I_0_0_t1b_t1b),
    .O_0_0_t0b(n402_O_0_0_t0b),
    .O_0_0_t1b_t0b(n402_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n402_O_0_0_t1b_t1b)
  );
  Map2S_34 n403 ( // @[Top.scala 296:22]
    .valid_up(n403_valid_up),
    .valid_down(n403_valid_down),
    .I0_0_0_t0b(n403_I0_0_0_t0b),
    .I0_0_0_t1b_t0b(n403_I0_0_0_t1b_t0b),
    .I0_0_0_t1b_t1b(n403_I0_0_0_t1b_t1b),
    .I1_0_0_t0b(n403_I1_0_0_t0b),
    .I1_0_0_t1b_t0b(n403_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b(n403_I1_0_0_t1b_t1b),
    .O_0_0_t0b_t0b(n403_O_0_0_t0b_t0b),
    .O_0_0_t0b_t1b_t0b(n403_O_0_0_t0b_t1b_t0b),
    .O_0_0_t0b_t1b_t1b(n403_O_0_0_t0b_t1b_t1b),
    .O_0_0_t1b_t0b(n403_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b_t0b(n403_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b(n403_O_0_0_t1b_t1b_t1b)
  );
  Map2S_36 n411 ( // @[Top.scala 300:22]
    .valid_up(n411_valid_up),
    .valid_down(n411_valid_down),
    .I0_0_0(n411_I0_0_0),
    .I1_0_0_t0b_t0b(n411_I1_0_0_t0b_t0b),
    .I1_0_0_t0b_t1b_t0b(n411_I1_0_0_t0b_t1b_t0b),
    .I1_0_0_t0b_t1b_t1b(n411_I1_0_0_t0b_t1b_t1b),
    .I1_0_0_t1b_t0b(n411_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b_t0b(n411_I1_0_0_t1b_t1b_t0b),
    .I1_0_0_t1b_t1b_t1b(n411_I1_0_0_t1b_t1b_t1b),
    .O_0_0_t0b(n411_O_0_0_t0b),
    .O_0_0_t1b_t0b_t0b(n411_O_0_0_t1b_t0b_t0b),
    .O_0_0_t1b_t0b_t1b_t0b(n411_O_0_0_t1b_t0b_t1b_t0b),
    .O_0_0_t1b_t0b_t1b_t1b(n411_O_0_0_t1b_t0b_t1b_t1b),
    .O_0_0_t1b_t1b_t0b(n411_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t0b(n411_O_0_0_t1b_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t1b(n411_O_0_0_t1b_t1b_t1b_t1b)
  );
  MapS_44 n422 ( // @[Top.scala 304:22]
    .valid_up(n422_valid_up),
    .valid_down(n422_valid_down),
    .I_0_0_t0b(n422_I_0_0_t0b),
    .I_0_0_t1b_t0b_t0b(n422_I_0_0_t1b_t0b_t0b),
    .I_0_0_t1b_t0b_t1b_t0b(n422_I_0_0_t1b_t0b_t1b_t0b),
    .I_0_0_t1b_t0b_t1b_t1b(n422_I_0_0_t1b_t0b_t1b_t1b),
    .I_0_0_t1b_t1b_t0b(n422_I_0_0_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t0b(n422_I_0_0_t1b_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t1b(n422_I_0_0_t1b_t1b_t1b_t1b),
    .O_0_0_t0b(n422_O_0_0_t0b),
    .O_0_0_t1b_t0b(n422_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n422_O_0_0_t1b_t1b)
  );
  Map2S_34 n423 ( // @[Top.scala 307:22]
    .valid_up(n423_valid_up),
    .valid_down(n423_valid_down),
    .I0_0_0_t0b(n423_I0_0_0_t0b),
    .I0_0_0_t1b_t0b(n423_I0_0_0_t1b_t0b),
    .I0_0_0_t1b_t1b(n423_I0_0_0_t1b_t1b),
    .I1_0_0_t0b(n423_I1_0_0_t0b),
    .I1_0_0_t1b_t0b(n423_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b(n423_I1_0_0_t1b_t1b),
    .O_0_0_t0b_t0b(n423_O_0_0_t0b_t0b),
    .O_0_0_t0b_t1b_t0b(n423_O_0_0_t0b_t1b_t0b),
    .O_0_0_t0b_t1b_t1b(n423_O_0_0_t0b_t1b_t1b),
    .O_0_0_t1b_t0b(n423_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b_t0b(n423_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b(n423_O_0_0_t1b_t1b_t1b)
  );
  Map2S_36 n431 ( // @[Top.scala 311:22]
    .valid_up(n431_valid_up),
    .valid_down(n431_valid_down),
    .I0_0_0(n431_I0_0_0),
    .I1_0_0_t0b_t0b(n431_I1_0_0_t0b_t0b),
    .I1_0_0_t0b_t1b_t0b(n431_I1_0_0_t0b_t1b_t0b),
    .I1_0_0_t0b_t1b_t1b(n431_I1_0_0_t0b_t1b_t1b),
    .I1_0_0_t1b_t0b(n431_I1_0_0_t1b_t0b),
    .I1_0_0_t1b_t1b_t0b(n431_I1_0_0_t1b_t1b_t0b),
    .I1_0_0_t1b_t1b_t1b(n431_I1_0_0_t1b_t1b_t1b),
    .O_0_0_t0b(n431_O_0_0_t0b),
    .O_0_0_t1b_t0b_t0b(n431_O_0_0_t1b_t0b_t0b),
    .O_0_0_t1b_t0b_t1b_t0b(n431_O_0_0_t1b_t0b_t1b_t0b),
    .O_0_0_t1b_t0b_t1b_t1b(n431_O_0_0_t1b_t0b_t1b_t1b),
    .O_0_0_t1b_t1b_t0b(n431_O_0_0_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t0b(n431_O_0_0_t1b_t1b_t1b_t0b),
    .O_0_0_t1b_t1b_t1b_t1b(n431_O_0_0_t1b_t1b_t1b_t1b)
  );
  MapS_44 n442 ( // @[Top.scala 315:22]
    .valid_up(n442_valid_up),
    .valid_down(n442_valid_down),
    .I_0_0_t0b(n442_I_0_0_t0b),
    .I_0_0_t1b_t0b_t0b(n442_I_0_0_t1b_t0b_t0b),
    .I_0_0_t1b_t0b_t1b_t0b(n442_I_0_0_t1b_t0b_t1b_t0b),
    .I_0_0_t1b_t0b_t1b_t1b(n442_I_0_0_t1b_t0b_t1b_t1b),
    .I_0_0_t1b_t1b_t0b(n442_I_0_0_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t0b(n442_I_0_0_t1b_t1b_t1b_t0b),
    .I_0_0_t1b_t1b_t1b_t1b(n442_I_0_0_t1b_t1b_t1b_t1b),
    .O_0_0_t0b(n442_O_0_0_t0b),
    .O_0_0_t1b_t0b(n442_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n442_O_0_0_t1b_t1b)
  );
  assign valid_down = n442_valid_down; // @[Top.scala 319:16]
  assign O_0_0_t0b = n442_O_0_0_t0b; // @[Top.scala 318:7]
  assign O_0_0_t1b_t0b = n442_O_0_0_t1b_t0b; // @[Top.scala 318:7]
  assign O_0_0_t1b_t1b = n442_O_0_0_t1b_t1b; // @[Top.scala 318:7]
  assign n152_valid_up = valid_up; // @[Top.scala 118:19]
  assign n152_I_0_0_t0b = I1_0_0_t0b; // @[Top.scala 117:12]
  assign n430_clock = clock;
  assign n430_reset = reset;
  assign n430_valid_up = n152_valid_down; // @[Top.scala 121:19]
  assign n430_I_0_0 = n152_O_0_0; // @[Top.scala 120:12]
  assign n157_valid_up = valid_up; // @[Top.scala 124:19]
  assign n157_I_0_0_t1b = I1_0_0_t1b; // @[Top.scala 123:12]
  assign n360_clock = clock;
  assign n360_reset = reset;
  assign n360_valid_up = n157_valid_down; // @[Top.scala 127:19]
  assign n360_I_0_0 = n157_O_0_0; // @[Top.scala 126:12]
  assign n159_valid_up = valid_up; // @[Top.scala 130:19]
  assign n159_I_1_0 = I0_1_0; // @[Top.scala 129:12]
  assign n159_I_1_1 = I0_1_1; // @[Top.scala 129:12]
  assign n159_I_1_2 = I0_1_2; // @[Top.scala 129:12]
  assign n162_valid_up = n159_valid_down; // @[Top.scala 133:19]
  assign n162_I_0_0 = n159_O_0_0; // @[Top.scala 132:12]
  assign n165_valid_up = n159_valid_down; // @[Top.scala 136:19]
  assign n165_I_0_2 = n159_O_0_2; // @[Top.scala 135:12]
  assign n166_valid_up = n162_valid_down & n165_valid_down; // @[Top.scala 140:19]
  assign n166_I0_0_0 = n162_O_0_0; // @[Top.scala 138:13]
  assign n166_I1_0_0 = n165_O_0_0; // @[Top.scala 139:13]
  assign n177_valid_up = n166_valid_down; // @[Top.scala 143:19]
  assign n177_I_0_0_t0b = n166_O_0_0_t0b; // @[Top.scala 142:12]
  assign n177_I_0_0_t1b = n166_O_0_0_t1b; // @[Top.scala 142:12]
  assign n184_clock = clock;
  assign n184_reset = reset;
  assign n184_valid_up = n177_valid_down; // @[Top.scala 146:19]
  assign n184_I_0_0 = n177_O_0_0; // @[Top.scala 145:12]
  assign n189_valid_up = n184_valid_down; // @[Top.scala 149:19]
  assign n189_I_0_0_t0b = n184_O_0_0_t0b; // @[Top.scala 148:12]
  assign n189_I_0_0_t1b = n184_O_0_0_t1b; // @[Top.scala 148:12]
  assign n192_valid_up = n159_valid_down; // @[Top.scala 152:19]
  assign n192_I_0_1 = n159_O_0_1; // @[Top.scala 151:12]
  assign n193_valid_up = valid_up; // @[Top.scala 155:19]
  assign n193_I_0_0 = I0_0_0; // @[Top.scala 154:12]
  assign n193_I_0_1 = I0_0_1; // @[Top.scala 154:12]
  assign n193_I_0_2 = I0_0_2; // @[Top.scala 154:12]
  assign n196_valid_up = n193_valid_down; // @[Top.scala 158:19]
  assign n196_I_0_1 = n193_O_0_1; // @[Top.scala 157:12]
  assign n197_valid_up = valid_up; // @[Top.scala 161:19]
  assign n197_I_2_0 = I0_2_0; // @[Top.scala 160:12]
  assign n197_I_2_1 = I0_2_1; // @[Top.scala 160:12]
  assign n197_I_2_2 = I0_2_2; // @[Top.scala 160:12]
  assign n200_valid_up = n197_valid_down; // @[Top.scala 164:19]
  assign n200_I_0_1 = n197_O_0_1; // @[Top.scala 163:12]
  assign n201_valid_up = n196_valid_down & n200_valid_down; // @[Top.scala 168:19]
  assign n201_I0_0_0 = n196_O_0_0; // @[Top.scala 166:13]
  assign n201_I1_0_0 = n200_O_0_0; // @[Top.scala 167:13]
  assign n212_valid_up = n201_valid_down; // @[Top.scala 171:19]
  assign n212_I_0_0_t0b = n201_O_0_0_t0b; // @[Top.scala 170:12]
  assign n212_I_0_0_t1b = n201_O_0_0_t1b; // @[Top.scala 170:12]
  assign n219_clock = clock;
  assign n219_reset = reset;
  assign n219_valid_up = n212_valid_down; // @[Top.scala 174:19]
  assign n219_I_0_0 = n212_O_0_0; // @[Top.scala 173:12]
  assign n224_valid_up = n219_valid_down; // @[Top.scala 177:19]
  assign n224_I_0_0_t0b = n219_O_0_0_t0b; // @[Top.scala 176:12]
  assign n224_I_0_0_t1b = n219_O_0_0_t1b; // @[Top.scala 176:12]
  assign n225_valid_up = n192_valid_down & n224_valid_down; // @[Top.scala 181:19]
  assign n225_I0_0_0 = n192_O_0_0; // @[Top.scala 179:13]
  assign n225_I1_0_0 = n224_O_0_0; // @[Top.scala 180:13]
  assign n232_valid_up = n189_valid_down & n225_valid_down; // @[Top.scala 185:19]
  assign n232_I0_0_0 = n189_O_0_0; // @[Top.scala 183:13]
  assign n232_I1_0_0_t0b = n225_O_0_0_t0b; // @[Top.scala 184:13]
  assign n232_I1_0_0_t1b = n225_O_0_0_t1b; // @[Top.scala 184:13]
  assign n352_clock = clock;
  assign n352_reset = reset;
  assign n352_valid_up = n232_valid_down; // @[Top.scala 188:19]
  assign n352_I_0_0_t0b = n232_O_0_0_t0b; // @[Top.scala 187:12]
  assign n352_I_0_0_t1b_t0b = n232_O_0_0_t1b_t0b; // @[Top.scala 187:12]
  assign n352_I_0_0_t1b_t1b = n232_O_0_0_t1b_t1b; // @[Top.scala 187:12]
  assign n344_clock = clock;
  assign n344_reset = reset;
  assign n344_valid_up = n192_valid_down; // @[Top.scala 191:19]
  assign n344_I_0_0 = n192_O_0_0; // @[Top.scala 190:12]
  assign n239_valid_up = n162_valid_down & n196_valid_down; // @[Top.scala 195:19]
  assign n239_I0_0_0 = n162_O_0_0; // @[Top.scala 193:13]
  assign n239_I1_0_0 = n196_O_0_0; // @[Top.scala 194:13]
  assign n246_valid_up = n239_valid_down & n165_valid_down; // @[Top.scala 199:19]
  assign n246_I0_0_0_0 = n239_O_0_0_0; // @[Top.scala 197:13]
  assign n246_I0_0_0_1 = n239_O_0_0_1; // @[Top.scala 197:13]
  assign n246_I1_0_0 = n165_O_0_0; // @[Top.scala 198:13]
  assign n253_valid_up = n246_valid_down & n200_valid_down; // @[Top.scala 203:19]
  assign n253_I0_0_0_0 = n246_O_0_0_0; // @[Top.scala 201:13]
  assign n253_I0_0_0_1 = n246_O_0_0_1; // @[Top.scala 201:13]
  assign n253_I0_0_0_2 = n246_O_0_0_2; // @[Top.scala 201:13]
  assign n253_I1_0_0 = n200_O_0_0; // @[Top.scala 202:13]
  assign n264_valid_up = n253_valid_down; // @[Top.scala 206:19]
  assign n264_I_0_0_0 = n253_O_0_0_0; // @[Top.scala 205:12]
  assign n264_I_0_0_1 = n253_O_0_0_1; // @[Top.scala 205:12]
  assign n264_I_0_0_2 = n253_O_0_0_2; // @[Top.scala 205:12]
  assign n264_I_0_0_3 = n253_O_0_0_3; // @[Top.scala 205:12]
  assign n269_clock = clock;
  assign n269_reset = reset;
  assign n269_valid_up = n264_valid_down; // @[Top.scala 209:19]
  assign n269_I_0_0 = n264_O_0_0; // @[Top.scala 208:12]
  assign n269_I_0_1 = n264_O_0_1; // @[Top.scala 208:12]
  assign n269_I_0_2 = n264_O_0_2; // @[Top.scala 208:12]
  assign n269_I_0_3 = n264_O_0_3; // @[Top.scala 208:12]
  assign n276_clock = clock;
  assign n276_reset = reset;
  assign n276_valid_up = n269_valid_down; // @[Top.scala 212:19]
  assign n276_I_0_0 = n269_O_0_0; // @[Top.scala 211:12]
  assign n281_valid_up = n276_valid_down; // @[Top.scala 215:19]
  assign n281_I_0_0_t0b = n276_O_0_0_t0b; // @[Top.scala 214:12]
  assign n281_I_0_0_t1b = n276_O_0_0_t1b; // @[Top.scala 214:12]
  assign n284_valid_up = n193_valid_down; // @[Top.scala 218:19]
  assign n284_I_0_0 = n193_O_0_0; // @[Top.scala 217:12]
  assign n287_valid_up = n193_valid_down; // @[Top.scala 221:19]
  assign n287_I_0_2 = n193_O_0_2; // @[Top.scala 220:12]
  assign n288_valid_up = n284_valid_down & n287_valid_down; // @[Top.scala 225:19]
  assign n288_I0_0_0 = n284_O_0_0; // @[Top.scala 223:13]
  assign n288_I1_0_0 = n287_O_0_0; // @[Top.scala 224:13]
  assign n297_valid_up = n197_valid_down; // @[Top.scala 228:19]
  assign n297_I_0_0 = n197_O_0_0; // @[Top.scala 227:12]
  assign n298_valid_up = n288_valid_down & n297_valid_down; // @[Top.scala 232:19]
  assign n298_I0_0_0_0 = n288_O_0_0_0; // @[Top.scala 230:13]
  assign n298_I0_0_0_1 = n288_O_0_0_1; // @[Top.scala 230:13]
  assign n298_I1_0_0 = n297_O_0_0; // @[Top.scala 231:13]
  assign n307_valid_up = n197_valid_down; // @[Top.scala 235:19]
  assign n307_I_0_2 = n197_O_0_2; // @[Top.scala 234:12]
  assign n308_valid_up = n298_valid_down & n307_valid_down; // @[Top.scala 239:19]
  assign n308_I0_0_0_0 = n298_O_0_0_0; // @[Top.scala 237:13]
  assign n308_I0_0_0_1 = n298_O_0_0_1; // @[Top.scala 237:13]
  assign n308_I0_0_0_2 = n298_O_0_0_2; // @[Top.scala 237:13]
  assign n308_I1_0_0 = n307_O_0_0; // @[Top.scala 238:13]
  assign n319_valid_up = n308_valid_down; // @[Top.scala 242:19]
  assign n319_I_0_0_0 = n308_O_0_0_0; // @[Top.scala 241:12]
  assign n319_I_0_0_1 = n308_O_0_0_1; // @[Top.scala 241:12]
  assign n319_I_0_0_2 = n308_O_0_0_2; // @[Top.scala 241:12]
  assign n319_I_0_0_3 = n308_O_0_0_3; // @[Top.scala 241:12]
  assign n324_clock = clock;
  assign n324_reset = reset;
  assign n324_valid_up = n319_valid_down; // @[Top.scala 245:19]
  assign n324_I_0_0 = n319_O_0_0; // @[Top.scala 244:12]
  assign n324_I_0_1 = n319_O_0_1; // @[Top.scala 244:12]
  assign n324_I_0_2 = n319_O_0_2; // @[Top.scala 244:12]
  assign n324_I_0_3 = n319_O_0_3; // @[Top.scala 244:12]
  assign n331_clock = clock;
  assign n331_reset = reset;
  assign n331_valid_up = n324_valid_down; // @[Top.scala 248:19]
  assign n331_I_0_0 = n324_O_0_0; // @[Top.scala 247:12]
  assign n336_valid_up = n331_valid_down; // @[Top.scala 251:19]
  assign n336_I_0_0_t0b = n331_O_0_0_t0b; // @[Top.scala 250:12]
  assign n336_I_0_0_t1b = n331_O_0_0_t1b; // @[Top.scala 250:12]
  assign n337_valid_up = n281_valid_down & n336_valid_down; // @[Top.scala 255:19]
  assign n337_I0_0_0 = n281_O_0_0; // @[Top.scala 253:13]
  assign n337_I1_0_0 = n336_O_0_0; // @[Top.scala 254:13]
  assign n345_valid_up = n344_valid_down & n337_valid_down; // @[Top.scala 259:19]
  assign n345_I0_0_0 = n344_O_0_0; // @[Top.scala 257:13]
  assign n345_I1_0_0_t0b = n337_O_0_0_t0b; // @[Top.scala 258:13]
  assign n345_I1_0_0_t1b = n337_O_0_0_t1b; // @[Top.scala 258:13]
  assign n353_valid_up = n352_valid_down & n345_valid_down; // @[Top.scala 263:19]
  assign n353_I0_0_0_t0b = n352_O_0_0_t0b; // @[Top.scala 261:13]
  assign n353_I0_0_0_t1b_t0b = n352_O_0_0_t1b_t0b; // @[Top.scala 261:13]
  assign n353_I0_0_0_t1b_t1b = n352_O_0_0_t1b_t1b; // @[Top.scala 261:13]
  assign n353_I1_0_0_t0b = n345_O_0_0_t0b; // @[Top.scala 262:13]
  assign n353_I1_0_0_t1b_t0b = n345_O_0_0_t1b_t0b; // @[Top.scala 262:13]
  assign n353_I1_0_0_t1b_t1b = n345_O_0_0_t1b_t1b; // @[Top.scala 262:13]
  assign n361_valid_up = n360_valid_down & n353_valid_down; // @[Top.scala 267:19]
  assign n361_I0_0_0 = n360_O_0_0; // @[Top.scala 265:13]
  assign n361_I1_0_0_t0b_t0b = n353_O_0_0_t0b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t0b_t1b_t0b = n353_O_0_0_t0b_t1b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t0b_t1b_t1b = n353_O_0_0_t0b_t1b_t1b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t1b_t0b = n353_O_0_0_t1b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t1b_t1b_t0b = n353_O_0_0_t1b_t1b_t0b; // @[Top.scala 266:13]
  assign n361_I1_0_0_t1b_t1b_t1b = n353_O_0_0_t1b_t1b_t1b; // @[Top.scala 266:13]
  assign n372_valid_up = n361_valid_down; // @[Top.scala 270:19]
  assign n372_I_0_0_t0b = n361_O_0_0_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t0b_t0b = n361_O_0_0_t1b_t0b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t0b_t1b_t0b = n361_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t0b_t1b_t1b = n361_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t1b_t0b = n361_O_0_0_t1b_t1b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t1b_t1b_t0b = n361_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 269:12]
  assign n372_I_0_0_t1b_t1b_t1b_t1b = n361_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 269:12]
  assign n410_clock = clock;
  assign n410_reset = reset;
  assign n410_valid_up = n157_valid_down; // @[Top.scala 273:19]
  assign n410_I_0_0 = n157_O_0_0; // @[Top.scala 272:12]
  assign n373_clock = clock;
  assign n373_reset = reset;
  assign n373_valid_up = n192_valid_down; // @[Top.scala 276:19]
  assign n373_I_0_0 = n192_O_0_0; // @[Top.scala 275:12]
  assign n374_valid_up = n281_valid_down & n373_valid_down; // @[Top.scala 280:19]
  assign n374_I0_0_0 = n281_O_0_0; // @[Top.scala 278:13]
  assign n374_I1_0_0 = n373_O_0_0; // @[Top.scala 279:13]
  assign n381_valid_up = n336_valid_down & n374_valid_down; // @[Top.scala 284:19]
  assign n381_I0_0_0 = n336_O_0_0; // @[Top.scala 282:13]
  assign n381_I1_0_0_t0b = n374_O_0_0_t0b; // @[Top.scala 283:13]
  assign n381_I1_0_0_t1b = n374_O_0_0_t1b; // @[Top.scala 283:13]
  assign n388_valid_up = n192_valid_down & n189_valid_down; // @[Top.scala 288:19]
  assign n388_I0_0_0 = n192_O_0_0; // @[Top.scala 286:13]
  assign n388_I1_0_0 = n189_O_0_0; // @[Top.scala 287:13]
  assign n395_valid_up = n224_valid_down & n388_valid_down; // @[Top.scala 292:19]
  assign n395_I0_0_0 = n224_O_0_0; // @[Top.scala 290:13]
  assign n395_I1_0_0_t0b = n388_O_0_0_t0b; // @[Top.scala 291:13]
  assign n395_I1_0_0_t1b = n388_O_0_0_t1b; // @[Top.scala 291:13]
  assign n402_clock = clock;
  assign n402_reset = reset;
  assign n402_valid_up = n395_valid_down; // @[Top.scala 295:19]
  assign n402_I_0_0_t0b = n395_O_0_0_t0b; // @[Top.scala 294:12]
  assign n402_I_0_0_t1b_t0b = n395_O_0_0_t1b_t0b; // @[Top.scala 294:12]
  assign n402_I_0_0_t1b_t1b = n395_O_0_0_t1b_t1b; // @[Top.scala 294:12]
  assign n403_valid_up = n381_valid_down & n402_valid_down; // @[Top.scala 299:19]
  assign n403_I0_0_0_t0b = n381_O_0_0_t0b; // @[Top.scala 297:13]
  assign n403_I0_0_0_t1b_t0b = n381_O_0_0_t1b_t0b; // @[Top.scala 297:13]
  assign n403_I0_0_0_t1b_t1b = n381_O_0_0_t1b_t1b; // @[Top.scala 297:13]
  assign n403_I1_0_0_t0b = n402_O_0_0_t0b; // @[Top.scala 298:13]
  assign n403_I1_0_0_t1b_t0b = n402_O_0_0_t1b_t0b; // @[Top.scala 298:13]
  assign n403_I1_0_0_t1b_t1b = n402_O_0_0_t1b_t1b; // @[Top.scala 298:13]
  assign n411_valid_up = n410_valid_down & n403_valid_down; // @[Top.scala 303:19]
  assign n411_I0_0_0 = n410_O_0_0; // @[Top.scala 301:13]
  assign n411_I1_0_0_t0b_t0b = n403_O_0_0_t0b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t0b_t1b_t0b = n403_O_0_0_t0b_t1b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t0b_t1b_t1b = n403_O_0_0_t0b_t1b_t1b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t1b_t0b = n403_O_0_0_t1b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t1b_t1b_t0b = n403_O_0_0_t1b_t1b_t0b; // @[Top.scala 302:13]
  assign n411_I1_0_0_t1b_t1b_t1b = n403_O_0_0_t1b_t1b_t1b; // @[Top.scala 302:13]
  assign n422_valid_up = n411_valid_down; // @[Top.scala 306:19]
  assign n422_I_0_0_t0b = n411_O_0_0_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t0b_t0b = n411_O_0_0_t1b_t0b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t0b_t1b_t0b = n411_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t0b_t1b_t1b = n411_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t1b_t0b = n411_O_0_0_t1b_t1b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t1b_t1b_t0b = n411_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 305:12]
  assign n422_I_0_0_t1b_t1b_t1b_t1b = n411_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 305:12]
  assign n423_valid_up = n372_valid_down & n422_valid_down; // @[Top.scala 310:19]
  assign n423_I0_0_0_t0b = n372_O_0_0_t0b; // @[Top.scala 308:13]
  assign n423_I0_0_0_t1b_t0b = n372_O_0_0_t1b_t0b; // @[Top.scala 308:13]
  assign n423_I0_0_0_t1b_t1b = n372_O_0_0_t1b_t1b; // @[Top.scala 308:13]
  assign n423_I1_0_0_t0b = n422_O_0_0_t0b; // @[Top.scala 309:13]
  assign n423_I1_0_0_t1b_t0b = n422_O_0_0_t1b_t0b; // @[Top.scala 309:13]
  assign n423_I1_0_0_t1b_t1b = n422_O_0_0_t1b_t1b; // @[Top.scala 309:13]
  assign n431_valid_up = n430_valid_down & n423_valid_down; // @[Top.scala 314:19]
  assign n431_I0_0_0 = n430_O_0_0; // @[Top.scala 312:13]
  assign n431_I1_0_0_t0b_t0b = n423_O_0_0_t0b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t0b_t1b_t0b = n423_O_0_0_t0b_t1b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t0b_t1b_t1b = n423_O_0_0_t0b_t1b_t1b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t1b_t0b = n423_O_0_0_t1b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t1b_t1b_t0b = n423_O_0_0_t1b_t1b_t0b; // @[Top.scala 313:13]
  assign n431_I1_0_0_t1b_t1b_t1b = n423_O_0_0_t1b_t1b_t1b; // @[Top.scala 313:13]
  assign n442_valid_up = n431_valid_down; // @[Top.scala 317:19]
  assign n442_I_0_0_t0b = n431_O_0_0_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t0b_t0b = n431_O_0_0_t1b_t0b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t0b_t1b_t0b = n431_O_0_0_t1b_t0b_t1b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t0b_t1b_t1b = n431_O_0_0_t1b_t0b_t1b_t1b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t1b_t0b = n431_O_0_0_t1b_t1b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t1b_t1b_t0b = n431_O_0_0_t1b_t1b_t1b_t0b; // @[Top.scala 316:12]
  assign n442_I_0_0_t1b_t1b_t1b_t1b = n431_O_0_0_t1b_t1b_t1b_t1b; // @[Top.scala 316:12]
endmodule
module Map2S_53(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_0_2_0,
  input  [31:0] I0_0_2_1,
  input  [31:0] I0_0_2_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_1_2_0,
  input  [31:0] I0_1_2_1,
  input  [31:0] I0_1_2_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_2_2_0,
  input  [31:0] I0_2_2_1,
  input  [31:0] I0_2_2_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_3_2_0,
  input  [31:0] I0_3_2_1,
  input  [31:0] I0_3_2_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_4_2_0,
  input  [31:0] I0_4_2_1,
  input  [31:0] I0_4_2_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_5_2_0,
  input  [31:0] I0_5_2_1,
  input  [31:0] I0_5_2_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_6_2_0,
  input  [31:0] I0_6_2_1,
  input  [31:0] I0_6_2_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I0_7_2_0,
  input  [31:0] I0_7_2_1,
  input  [31:0] I0_7_2_2,
  input  [31:0] I0_8_0_0,
  input  [31:0] I0_8_0_1,
  input  [31:0] I0_8_0_2,
  input  [31:0] I0_8_1_0,
  input  [31:0] I0_8_1_1,
  input  [31:0] I0_8_1_2,
  input  [31:0] I0_8_2_0,
  input  [31:0] I0_8_2_1,
  input  [31:0] I0_8_2_2,
  input  [31:0] I0_9_0_0,
  input  [31:0] I0_9_0_1,
  input  [31:0] I0_9_0_2,
  input  [31:0] I0_9_1_0,
  input  [31:0] I0_9_1_1,
  input  [31:0] I0_9_1_2,
  input  [31:0] I0_9_2_0,
  input  [31:0] I0_9_2_1,
  input  [31:0] I0_9_2_2,
  input  [31:0] I0_10_0_0,
  input  [31:0] I0_10_0_1,
  input  [31:0] I0_10_0_2,
  input  [31:0] I0_10_1_0,
  input  [31:0] I0_10_1_1,
  input  [31:0] I0_10_1_2,
  input  [31:0] I0_10_2_0,
  input  [31:0] I0_10_2_1,
  input  [31:0] I0_10_2_2,
  input  [31:0] I0_11_0_0,
  input  [31:0] I0_11_0_1,
  input  [31:0] I0_11_0_2,
  input  [31:0] I0_11_1_0,
  input  [31:0] I0_11_1_1,
  input  [31:0] I0_11_1_2,
  input  [31:0] I0_11_2_0,
  input  [31:0] I0_11_2_1,
  input  [31:0] I0_11_2_2,
  input  [31:0] I0_12_0_0,
  input  [31:0] I0_12_0_1,
  input  [31:0] I0_12_0_2,
  input  [31:0] I0_12_1_0,
  input  [31:0] I0_12_1_1,
  input  [31:0] I0_12_1_2,
  input  [31:0] I0_12_2_0,
  input  [31:0] I0_12_2_1,
  input  [31:0] I0_12_2_2,
  input  [31:0] I0_13_0_0,
  input  [31:0] I0_13_0_1,
  input  [31:0] I0_13_0_2,
  input  [31:0] I0_13_1_0,
  input  [31:0] I0_13_1_1,
  input  [31:0] I0_13_1_2,
  input  [31:0] I0_13_2_0,
  input  [31:0] I0_13_2_1,
  input  [31:0] I0_13_2_2,
  input  [31:0] I0_14_0_0,
  input  [31:0] I0_14_0_1,
  input  [31:0] I0_14_0_2,
  input  [31:0] I0_14_1_0,
  input  [31:0] I0_14_1_1,
  input  [31:0] I0_14_1_2,
  input  [31:0] I0_14_2_0,
  input  [31:0] I0_14_2_1,
  input  [31:0] I0_14_2_2,
  input  [31:0] I0_15_0_0,
  input  [31:0] I0_15_0_1,
  input  [31:0] I0_15_0_2,
  input  [31:0] I0_15_1_0,
  input  [31:0] I0_15_1_1,
  input  [31:0] I0_15_1_2,
  input  [31:0] I0_15_2_0,
  input  [31:0] I0_15_2_1,
  input  [31:0] I0_15_2_2,
  input         I1_0_0_0_t0b,
  input         I1_0_0_0_t1b,
  input         I1_1_0_0_t0b,
  input         I1_1_0_0_t1b,
  input         I1_2_0_0_t0b,
  input         I1_2_0_0_t1b,
  input         I1_3_0_0_t0b,
  input         I1_3_0_0_t1b,
  input         I1_4_0_0_t0b,
  input         I1_4_0_0_t1b,
  input         I1_5_0_0_t0b,
  input         I1_5_0_0_t1b,
  input         I1_6_0_0_t0b,
  input         I1_6_0_0_t1b,
  input         I1_7_0_0_t0b,
  input         I1_7_0_0_t1b,
  input         I1_8_0_0_t0b,
  input         I1_8_0_0_t1b,
  input         I1_9_0_0_t0b,
  input         I1_9_0_0_t1b,
  input         I1_10_0_0_t0b,
  input         I1_10_0_0_t1b,
  input         I1_11_0_0_t0b,
  input         I1_11_0_0_t1b,
  input         I1_12_0_0_t0b,
  input         I1_12_0_0_t1b,
  input         I1_13_0_0_t0b,
  input         I1_13_0_0_t1b,
  input         I1_14_0_0_t0b,
  input         I1_14_0_0_t1b,
  input         I1_15_0_0_t0b,
  input         I1_15_0_0_t1b,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b,
  output [31:0] O_8_0_0_t0b,
  output [31:0] O_8_0_0_t1b_t0b,
  output [31:0] O_8_0_0_t1b_t1b,
  output [31:0] O_9_0_0_t0b,
  output [31:0] O_9_0_0_t1b_t0b,
  output [31:0] O_9_0_0_t1b_t1b,
  output [31:0] O_10_0_0_t0b,
  output [31:0] O_10_0_0_t1b_t0b,
  output [31:0] O_10_0_0_t1b_t1b,
  output [31:0] O_11_0_0_t0b,
  output [31:0] O_11_0_0_t1b_t0b,
  output [31:0] O_11_0_0_t1b_t1b,
  output [31:0] O_12_0_0_t0b,
  output [31:0] O_12_0_0_t1b_t0b,
  output [31:0] O_12_0_0_t1b_t1b,
  output [31:0] O_13_0_0_t0b,
  output [31:0] O_13_0_0_t1b_t0b,
  output [31:0] O_13_0_0_t1b_t1b,
  output [31:0] O_14_0_0_t0b,
  output [31:0] O_14_0_0_t1b_t0b,
  output [31:0] O_14_0_0_t1b_t1b,
  output [31:0] O_15_0_0_t0b,
  output [31:0] O_15_0_0_t1b_t0b,
  output [31:0] O_15_0_0_t1b_t1b
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2_0; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2_1; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_I0_2_2; // @[Map2S.scala 9:22]
  wire  fst_op_I1_0_0_t0b; // @[Map2S.scala 9:22]
  wire  fst_op_I1_0_0_t1b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0_t1b_t0b; // @[Map2S.scala 9:22]
  wire [31:0] fst_op_O_0_0_t1b_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_clock; // @[Map2S.scala 10:86]
  wire  other_ops_0_reset; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_0_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_0_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_0_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_clock; // @[Map2S.scala 10:86]
  wire  other_ops_1_reset; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_1_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_1_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_2_clock; // @[Map2S.scala 10:86]
  wire  other_ops_2_reset; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_2_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_2_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_3_clock; // @[Map2S.scala 10:86]
  wire  other_ops_3_reset; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_3_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_3_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_4_clock; // @[Map2S.scala 10:86]
  wire  other_ops_4_reset; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_4_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_4_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_5_clock; // @[Map2S.scala 10:86]
  wire  other_ops_5_reset; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_5_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_5_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_6_clock; // @[Map2S.scala 10:86]
  wire  other_ops_6_reset; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_6_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_6_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_7_clock; // @[Map2S.scala 10:86]
  wire  other_ops_7_reset; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_7_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_7_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_8_clock; // @[Map2S.scala 10:86]
  wire  other_ops_8_reset; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_8_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_8_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_9_clock; // @[Map2S.scala 10:86]
  wire  other_ops_9_reset; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_9_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_9_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_10_clock; // @[Map2S.scala 10:86]
  wire  other_ops_10_reset; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_10_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_10_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_11_clock; // @[Map2S.scala 10:86]
  wire  other_ops_11_reset; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_11_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_11_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_12_clock; // @[Map2S.scala 10:86]
  wire  other_ops_12_reset; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_12_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_12_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_13_clock; // @[Map2S.scala 10:86]
  wire  other_ops_13_reset; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_13_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_13_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_14_clock; // @[Map2S.scala 10:86]
  wire  other_ops_14_reset; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_0_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_1_2; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_2_0; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_2_1; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_I0_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_I1_0_0_t0b; // @[Map2S.scala 10:86]
  wire  other_ops_14_I1_0_0_t1b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_0_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_0_t1b_t0b; // @[Map2S.scala 10:86]
  wire [31:0] other_ops_14_O_0_0_t1b_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Module_6 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I0_2_0(fst_op_I0_2_0),
    .I0_2_1(fst_op_I0_2_1),
    .I0_2_2(fst_op_I0_2_2),
    .I1_0_0_t0b(fst_op_I1_0_0_t0b),
    .I1_0_0_t1b(fst_op_I1_0_0_t1b),
    .O_0_0_t0b(fst_op_O_0_0_t0b),
    .O_0_0_t1b_t0b(fst_op_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(fst_op_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_0 ( // @[Map2S.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I0_2_0(other_ops_0_I0_2_0),
    .I0_2_1(other_ops_0_I0_2_1),
    .I0_2_2(other_ops_0_I0_2_2),
    .I1_0_0_t0b(other_ops_0_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_0_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_0_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_0_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_0_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_1 ( // @[Map2S.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I0_2_0(other_ops_1_I0_2_0),
    .I0_2_1(other_ops_1_I0_2_1),
    .I0_2_2(other_ops_1_I0_2_2),
    .I1_0_0_t0b(other_ops_1_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_1_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_1_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_1_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_1_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_2 ( // @[Map2S.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I0_2_0(other_ops_2_I0_2_0),
    .I0_2_1(other_ops_2_I0_2_1),
    .I0_2_2(other_ops_2_I0_2_2),
    .I1_0_0_t0b(other_ops_2_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_2_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_2_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_2_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_2_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_3 ( // @[Map2S.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I0_2_0(other_ops_3_I0_2_0),
    .I0_2_1(other_ops_3_I0_2_1),
    .I0_2_2(other_ops_3_I0_2_2),
    .I1_0_0_t0b(other_ops_3_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_3_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_3_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_3_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_3_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_4 ( // @[Map2S.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I0_2_0(other_ops_4_I0_2_0),
    .I0_2_1(other_ops_4_I0_2_1),
    .I0_2_2(other_ops_4_I0_2_2),
    .I1_0_0_t0b(other_ops_4_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_4_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_4_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_4_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_4_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_5 ( // @[Map2S.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I0_2_0(other_ops_5_I0_2_0),
    .I0_2_1(other_ops_5_I0_2_1),
    .I0_2_2(other_ops_5_I0_2_2),
    .I1_0_0_t0b(other_ops_5_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_5_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_5_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_5_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_5_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_6 ( // @[Map2S.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I0_2_0(other_ops_6_I0_2_0),
    .I0_2_1(other_ops_6_I0_2_1),
    .I0_2_2(other_ops_6_I0_2_2),
    .I1_0_0_t0b(other_ops_6_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_6_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_6_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_6_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_6_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_7 ( // @[Map2S.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I0_0_1(other_ops_7_I0_0_1),
    .I0_0_2(other_ops_7_I0_0_2),
    .I0_1_0(other_ops_7_I0_1_0),
    .I0_1_1(other_ops_7_I0_1_1),
    .I0_1_2(other_ops_7_I0_1_2),
    .I0_2_0(other_ops_7_I0_2_0),
    .I0_2_1(other_ops_7_I0_2_1),
    .I0_2_2(other_ops_7_I0_2_2),
    .I1_0_0_t0b(other_ops_7_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_7_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_7_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_7_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_7_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_8 ( // @[Map2S.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I0_0_1(other_ops_8_I0_0_1),
    .I0_0_2(other_ops_8_I0_0_2),
    .I0_1_0(other_ops_8_I0_1_0),
    .I0_1_1(other_ops_8_I0_1_1),
    .I0_1_2(other_ops_8_I0_1_2),
    .I0_2_0(other_ops_8_I0_2_0),
    .I0_2_1(other_ops_8_I0_2_1),
    .I0_2_2(other_ops_8_I0_2_2),
    .I1_0_0_t0b(other_ops_8_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_8_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_8_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_8_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_8_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_9 ( // @[Map2S.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I0_0_1(other_ops_9_I0_0_1),
    .I0_0_2(other_ops_9_I0_0_2),
    .I0_1_0(other_ops_9_I0_1_0),
    .I0_1_1(other_ops_9_I0_1_1),
    .I0_1_2(other_ops_9_I0_1_2),
    .I0_2_0(other_ops_9_I0_2_0),
    .I0_2_1(other_ops_9_I0_2_1),
    .I0_2_2(other_ops_9_I0_2_2),
    .I1_0_0_t0b(other_ops_9_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_9_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_9_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_9_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_9_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_10 ( // @[Map2S.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I0_0_1(other_ops_10_I0_0_1),
    .I0_0_2(other_ops_10_I0_0_2),
    .I0_1_0(other_ops_10_I0_1_0),
    .I0_1_1(other_ops_10_I0_1_1),
    .I0_1_2(other_ops_10_I0_1_2),
    .I0_2_0(other_ops_10_I0_2_0),
    .I0_2_1(other_ops_10_I0_2_1),
    .I0_2_2(other_ops_10_I0_2_2),
    .I1_0_0_t0b(other_ops_10_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_10_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_10_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_10_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_10_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_11 ( // @[Map2S.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I0_0_1(other_ops_11_I0_0_1),
    .I0_0_2(other_ops_11_I0_0_2),
    .I0_1_0(other_ops_11_I0_1_0),
    .I0_1_1(other_ops_11_I0_1_1),
    .I0_1_2(other_ops_11_I0_1_2),
    .I0_2_0(other_ops_11_I0_2_0),
    .I0_2_1(other_ops_11_I0_2_1),
    .I0_2_2(other_ops_11_I0_2_2),
    .I1_0_0_t0b(other_ops_11_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_11_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_11_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_11_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_11_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_12 ( // @[Map2S.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I0_0_1(other_ops_12_I0_0_1),
    .I0_0_2(other_ops_12_I0_0_2),
    .I0_1_0(other_ops_12_I0_1_0),
    .I0_1_1(other_ops_12_I0_1_1),
    .I0_1_2(other_ops_12_I0_1_2),
    .I0_2_0(other_ops_12_I0_2_0),
    .I0_2_1(other_ops_12_I0_2_1),
    .I0_2_2(other_ops_12_I0_2_2),
    .I1_0_0_t0b(other_ops_12_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_12_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_12_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_12_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_12_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_13 ( // @[Map2S.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I0_0_1(other_ops_13_I0_0_1),
    .I0_0_2(other_ops_13_I0_0_2),
    .I0_1_0(other_ops_13_I0_1_0),
    .I0_1_1(other_ops_13_I0_1_1),
    .I0_1_2(other_ops_13_I0_1_2),
    .I0_2_0(other_ops_13_I0_2_0),
    .I0_2_1(other_ops_13_I0_2_1),
    .I0_2_2(other_ops_13_I0_2_2),
    .I1_0_0_t0b(other_ops_13_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_13_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_13_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_13_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_13_O_0_0_t1b_t1b)
  );
  Module_6 other_ops_14 ( // @[Map2S.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I0_0_1(other_ops_14_I0_0_1),
    .I0_0_2(other_ops_14_I0_0_2),
    .I0_1_0(other_ops_14_I0_1_0),
    .I0_1_1(other_ops_14_I0_1_1),
    .I0_1_2(other_ops_14_I0_1_2),
    .I0_2_0(other_ops_14_I0_2_0),
    .I0_2_1(other_ops_14_I0_2_1),
    .I0_2_2(other_ops_14_I0_2_2),
    .I1_0_0_t0b(other_ops_14_I1_0_0_t0b),
    .I1_0_0_t1b(other_ops_14_I1_0_0_t1b),
    .O_0_0_t0b(other_ops_14_O_0_0_t0b),
    .O_0_0_t1b_t0b(other_ops_14_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(other_ops_14_O_0_0_t1b_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0_t0b = fst_op_O_0_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_0_t1b_t0b = fst_op_O_0_0_t1b_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_0_t1b_t1b = fst_op_O_0_0_t1b_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_0_t0b = other_ops_0_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_0_t1b_t0b = other_ops_0_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_0_t1b_t1b = other_ops_0_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_0_t0b = other_ops_1_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_0_t1b_t0b = other_ops_1_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_0_t1b_t1b = other_ops_1_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_3_0_0_t0b = other_ops_2_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_3_0_0_t1b_t0b = other_ops_2_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_3_0_0_t1b_t1b = other_ops_2_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_4_0_0_t0b = other_ops_3_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_4_0_0_t1b_t0b = other_ops_3_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_4_0_0_t1b_t1b = other_ops_3_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_5_0_0_t0b = other_ops_4_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_5_0_0_t1b_t0b = other_ops_4_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_5_0_0_t1b_t1b = other_ops_4_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_6_0_0_t0b = other_ops_5_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_6_0_0_t1b_t0b = other_ops_5_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_6_0_0_t1b_t1b = other_ops_5_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_7_0_0_t0b = other_ops_6_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_7_0_0_t1b_t0b = other_ops_6_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_7_0_0_t1b_t1b = other_ops_6_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_8_0_0_t0b = other_ops_7_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_8_0_0_t1b_t0b = other_ops_7_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_8_0_0_t1b_t1b = other_ops_7_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_9_0_0_t0b = other_ops_8_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_9_0_0_t1b_t0b = other_ops_8_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_9_0_0_t1b_t1b = other_ops_8_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_10_0_0_t0b = other_ops_9_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_10_0_0_t1b_t0b = other_ops_9_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_10_0_0_t1b_t1b = other_ops_9_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_11_0_0_t0b = other_ops_10_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_11_0_0_t1b_t0b = other_ops_10_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_11_0_0_t1b_t1b = other_ops_10_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_12_0_0_t0b = other_ops_11_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_12_0_0_t1b_t0b = other_ops_11_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_12_0_0_t1b_t1b = other_ops_11_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_13_0_0_t0b = other_ops_12_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_13_0_0_t1b_t0b = other_ops_12_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_13_0_0_t1b_t1b = other_ops_12_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_14_0_0_t0b = other_ops_13_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_14_0_0_t1b_t0b = other_ops_13_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_14_0_0_t1b_t1b = other_ops_13_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign O_15_0_0_t0b = other_ops_14_O_0_0_t0b; // @[Map2S.scala 24:12]
  assign O_15_0_0_t1b_t0b = other_ops_14_O_0_0_t1b_t0b; // @[Map2S.scala 24:12]
  assign O_15_0_0_t1b_t1b = other_ops_14_O_0_0_t1b_t1b; // @[Map2S.scala 24:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_2_0 = I0_0_2_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_2_1 = I0_0_2_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2_2 = I0_0_2_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0_0_t0b = I1_0_0_0_t0b; // @[Map2S.scala 18:13]
  assign fst_op_I1_0_0_t1b = I1_0_0_0_t1b; // @[Map2S.scala 18:13]
  assign other_ops_0_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_0_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2_0 = I0_1_2_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2_1 = I0_1_2_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2_2 = I0_1_2_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0_0_t0b = I1_1_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_0_0_t1b = I1_1_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_1_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_1_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2_0 = I0_2_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2_1 = I0_2_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2_2 = I0_2_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0_0_t0b = I1_2_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_0_0_t1b = I1_2_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_2_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_2_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2_0 = I0_3_2_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2_1 = I0_3_2_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2_2 = I0_3_2_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0_0_t0b = I1_3_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_0_0_t1b = I1_3_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_3_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_3_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2_0 = I0_4_2_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2_1 = I0_4_2_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2_2 = I0_4_2_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0_0_t0b = I1_4_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_0_0_t1b = I1_4_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_4_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_4_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2_0 = I0_5_2_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2_1 = I0_5_2_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2_2 = I0_5_2_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0_0_t0b = I1_5_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_0_0_t1b = I1_5_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_5_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_5_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2_0 = I0_6_2_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2_1 = I0_6_2_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2_2 = I0_6_2_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0_0_t0b = I1_6_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_0_0_t1b = I1_6_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_6_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_6_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2_0 = I0_7_2_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2_1 = I0_7_2_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2_2 = I0_7_2_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0_0_t0b = I1_7_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_0_0_t1b = I1_7_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_7_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_7_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1 = I0_8_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_2 = I0_8_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_0 = I0_8_1_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_1 = I0_8_1_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_2 = I0_8_1_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2_0 = I0_8_2_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2_1 = I0_8_2_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2_2 = I0_8_2_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0_0_t0b = I1_8_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_0_0_t1b = I1_8_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_8_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_8_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1 = I0_9_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_2 = I0_9_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_0 = I0_9_1_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_1 = I0_9_1_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_2 = I0_9_1_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2_0 = I0_9_2_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2_1 = I0_9_2_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2_2 = I0_9_2_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0_0_t0b = I1_9_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_0_0_t1b = I1_9_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_9_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_9_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1 = I0_10_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_2 = I0_10_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_0 = I0_10_1_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_1 = I0_10_1_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_2 = I0_10_1_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2_0 = I0_10_2_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2_1 = I0_10_2_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2_2 = I0_10_2_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0_0_t0b = I1_10_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_0_0_t1b = I1_10_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_10_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_10_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1 = I0_11_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_2 = I0_11_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_0 = I0_11_1_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_1 = I0_11_1_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_2 = I0_11_1_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2_0 = I0_11_2_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2_1 = I0_11_2_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2_2 = I0_11_2_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0_0_t0b = I1_11_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_0_0_t1b = I1_11_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_11_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_11_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1 = I0_12_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_2 = I0_12_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_0 = I0_12_1_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_1 = I0_12_1_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_2 = I0_12_1_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2_0 = I0_12_2_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2_1 = I0_12_2_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2_2 = I0_12_2_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0_0_t0b = I1_12_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_0_0_t1b = I1_12_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_12_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_12_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1 = I0_13_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_2 = I0_13_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_0 = I0_13_1_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_1 = I0_13_1_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_2 = I0_13_1_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2_0 = I0_13_2_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2_1 = I0_13_2_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2_2 = I0_13_2_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0_0_t0b = I1_13_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_0_0_t1b = I1_13_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_13_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_13_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1 = I0_14_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_2 = I0_14_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_0 = I0_14_1_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_1 = I0_14_1_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_2 = I0_14_1_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2_0 = I0_14_2_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2_1 = I0_14_2_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2_2 = I0_14_2_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0_0_t0b = I1_14_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_0_0_t1b = I1_14_0_0_t1b; // @[Map2S.scala 23:43]
  assign other_ops_14_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_14_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1 = I0_15_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_2 = I0_15_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_0 = I0_15_1_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_1 = I0_15_1_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_2 = I0_15_1_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2_0 = I0_15_2_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2_1 = I0_15_2_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2_2 = I0_15_2_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0_0_t0b = I1_15_0_0_t0b; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_0_0_t1b = I1_15_0_0_t1b; // @[Map2S.scala 23:43]
endmodule
module Map2T_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I0_0_0_0,
  input  [31:0] I0_0_0_1,
  input  [31:0] I0_0_0_2,
  input  [31:0] I0_0_1_0,
  input  [31:0] I0_0_1_1,
  input  [31:0] I0_0_1_2,
  input  [31:0] I0_0_2_0,
  input  [31:0] I0_0_2_1,
  input  [31:0] I0_0_2_2,
  input  [31:0] I0_1_0_0,
  input  [31:0] I0_1_0_1,
  input  [31:0] I0_1_0_2,
  input  [31:0] I0_1_1_0,
  input  [31:0] I0_1_1_1,
  input  [31:0] I0_1_1_2,
  input  [31:0] I0_1_2_0,
  input  [31:0] I0_1_2_1,
  input  [31:0] I0_1_2_2,
  input  [31:0] I0_2_0_0,
  input  [31:0] I0_2_0_1,
  input  [31:0] I0_2_0_2,
  input  [31:0] I0_2_1_0,
  input  [31:0] I0_2_1_1,
  input  [31:0] I0_2_1_2,
  input  [31:0] I0_2_2_0,
  input  [31:0] I0_2_2_1,
  input  [31:0] I0_2_2_2,
  input  [31:0] I0_3_0_0,
  input  [31:0] I0_3_0_1,
  input  [31:0] I0_3_0_2,
  input  [31:0] I0_3_1_0,
  input  [31:0] I0_3_1_1,
  input  [31:0] I0_3_1_2,
  input  [31:0] I0_3_2_0,
  input  [31:0] I0_3_2_1,
  input  [31:0] I0_3_2_2,
  input  [31:0] I0_4_0_0,
  input  [31:0] I0_4_0_1,
  input  [31:0] I0_4_0_2,
  input  [31:0] I0_4_1_0,
  input  [31:0] I0_4_1_1,
  input  [31:0] I0_4_1_2,
  input  [31:0] I0_4_2_0,
  input  [31:0] I0_4_2_1,
  input  [31:0] I0_4_2_2,
  input  [31:0] I0_5_0_0,
  input  [31:0] I0_5_0_1,
  input  [31:0] I0_5_0_2,
  input  [31:0] I0_5_1_0,
  input  [31:0] I0_5_1_1,
  input  [31:0] I0_5_1_2,
  input  [31:0] I0_5_2_0,
  input  [31:0] I0_5_2_1,
  input  [31:0] I0_5_2_2,
  input  [31:0] I0_6_0_0,
  input  [31:0] I0_6_0_1,
  input  [31:0] I0_6_0_2,
  input  [31:0] I0_6_1_0,
  input  [31:0] I0_6_1_1,
  input  [31:0] I0_6_1_2,
  input  [31:0] I0_6_2_0,
  input  [31:0] I0_6_2_1,
  input  [31:0] I0_6_2_2,
  input  [31:0] I0_7_0_0,
  input  [31:0] I0_7_0_1,
  input  [31:0] I0_7_0_2,
  input  [31:0] I0_7_1_0,
  input  [31:0] I0_7_1_1,
  input  [31:0] I0_7_1_2,
  input  [31:0] I0_7_2_0,
  input  [31:0] I0_7_2_1,
  input  [31:0] I0_7_2_2,
  input  [31:0] I0_8_0_0,
  input  [31:0] I0_8_0_1,
  input  [31:0] I0_8_0_2,
  input  [31:0] I0_8_1_0,
  input  [31:0] I0_8_1_1,
  input  [31:0] I0_8_1_2,
  input  [31:0] I0_8_2_0,
  input  [31:0] I0_8_2_1,
  input  [31:0] I0_8_2_2,
  input  [31:0] I0_9_0_0,
  input  [31:0] I0_9_0_1,
  input  [31:0] I0_9_0_2,
  input  [31:0] I0_9_1_0,
  input  [31:0] I0_9_1_1,
  input  [31:0] I0_9_1_2,
  input  [31:0] I0_9_2_0,
  input  [31:0] I0_9_2_1,
  input  [31:0] I0_9_2_2,
  input  [31:0] I0_10_0_0,
  input  [31:0] I0_10_0_1,
  input  [31:0] I0_10_0_2,
  input  [31:0] I0_10_1_0,
  input  [31:0] I0_10_1_1,
  input  [31:0] I0_10_1_2,
  input  [31:0] I0_10_2_0,
  input  [31:0] I0_10_2_1,
  input  [31:0] I0_10_2_2,
  input  [31:0] I0_11_0_0,
  input  [31:0] I0_11_0_1,
  input  [31:0] I0_11_0_2,
  input  [31:0] I0_11_1_0,
  input  [31:0] I0_11_1_1,
  input  [31:0] I0_11_1_2,
  input  [31:0] I0_11_2_0,
  input  [31:0] I0_11_2_1,
  input  [31:0] I0_11_2_2,
  input  [31:0] I0_12_0_0,
  input  [31:0] I0_12_0_1,
  input  [31:0] I0_12_0_2,
  input  [31:0] I0_12_1_0,
  input  [31:0] I0_12_1_1,
  input  [31:0] I0_12_1_2,
  input  [31:0] I0_12_2_0,
  input  [31:0] I0_12_2_1,
  input  [31:0] I0_12_2_2,
  input  [31:0] I0_13_0_0,
  input  [31:0] I0_13_0_1,
  input  [31:0] I0_13_0_2,
  input  [31:0] I0_13_1_0,
  input  [31:0] I0_13_1_1,
  input  [31:0] I0_13_1_2,
  input  [31:0] I0_13_2_0,
  input  [31:0] I0_13_2_1,
  input  [31:0] I0_13_2_2,
  input  [31:0] I0_14_0_0,
  input  [31:0] I0_14_0_1,
  input  [31:0] I0_14_0_2,
  input  [31:0] I0_14_1_0,
  input  [31:0] I0_14_1_1,
  input  [31:0] I0_14_1_2,
  input  [31:0] I0_14_2_0,
  input  [31:0] I0_14_2_1,
  input  [31:0] I0_14_2_2,
  input  [31:0] I0_15_0_0,
  input  [31:0] I0_15_0_1,
  input  [31:0] I0_15_0_2,
  input  [31:0] I0_15_1_0,
  input  [31:0] I0_15_1_1,
  input  [31:0] I0_15_1_2,
  input  [31:0] I0_15_2_0,
  input  [31:0] I0_15_2_1,
  input  [31:0] I0_15_2_2,
  input         I1_0_0_0_t0b,
  input         I1_0_0_0_t1b,
  input         I1_1_0_0_t0b,
  input         I1_1_0_0_t1b,
  input         I1_2_0_0_t0b,
  input         I1_2_0_0_t1b,
  input         I1_3_0_0_t0b,
  input         I1_3_0_0_t1b,
  input         I1_4_0_0_t0b,
  input         I1_4_0_0_t1b,
  input         I1_5_0_0_t0b,
  input         I1_5_0_0_t1b,
  input         I1_6_0_0_t0b,
  input         I1_6_0_0_t1b,
  input         I1_7_0_0_t0b,
  input         I1_7_0_0_t1b,
  input         I1_8_0_0_t0b,
  input         I1_8_0_0_t1b,
  input         I1_9_0_0_t0b,
  input         I1_9_0_0_t1b,
  input         I1_10_0_0_t0b,
  input         I1_10_0_0_t1b,
  input         I1_11_0_0_t0b,
  input         I1_11_0_0_t1b,
  input         I1_12_0_0_t0b,
  input         I1_12_0_0_t1b,
  input         I1_13_0_0_t0b,
  input         I1_13_0_0_t1b,
  input         I1_14_0_0_t0b,
  input         I1_14_0_0_t1b,
  input         I1_15_0_0_t0b,
  input         I1_15_0_0_t1b,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b,
  output [31:0] O_8_0_0_t0b,
  output [31:0] O_8_0_0_t1b_t0b,
  output [31:0] O_8_0_0_t1b_t1b,
  output [31:0] O_9_0_0_t0b,
  output [31:0] O_9_0_0_t1b_t0b,
  output [31:0] O_9_0_0_t1b_t1b,
  output [31:0] O_10_0_0_t0b,
  output [31:0] O_10_0_0_t1b_t0b,
  output [31:0] O_10_0_0_t1b_t1b,
  output [31:0] O_11_0_0_t0b,
  output [31:0] O_11_0_0_t1b_t0b,
  output [31:0] O_11_0_0_t1b_t1b,
  output [31:0] O_12_0_0_t0b,
  output [31:0] O_12_0_0_t1b_t0b,
  output [31:0] O_12_0_0_t1b_t1b,
  output [31:0] O_13_0_0_t0b,
  output [31:0] O_13_0_0_t1b_t0b,
  output [31:0] O_13_0_0_t1b_t1b,
  output [31:0] O_14_0_0_t0b,
  output [31:0] O_14_0_0_t1b_t0b,
  output [31:0] O_14_0_0_t1b_t1b,
  output [31:0] O_15_0_0_t0b,
  output [31:0] O_15_0_0_t1b_t0b,
  output [31:0] O_15_0_0_t1b_t1b
);
  wire  op_clock; // @[Map2T.scala 8:20]
  wire  op_reset; // @[Map2T.scala 8:20]
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_0_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_1_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_2_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_3_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_4_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_5_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_6_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_7_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_8_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_9_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_10_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_11_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_12_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_13_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_14_2_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_0_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_1_2; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_2_0; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_2_1; // @[Map2T.scala 8:20]
  wire [31:0] op_I0_15_2_2; // @[Map2T.scala 8:20]
  wire  op_I1_0_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_0_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_1_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_1_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_2_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_2_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_3_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_3_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_4_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_4_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_5_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_5_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_6_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_6_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_7_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_7_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_8_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_8_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_9_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_9_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_10_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_10_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_11_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_11_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_12_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_12_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_13_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_13_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_14_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_14_0_0_t1b; // @[Map2T.scala 8:20]
  wire  op_I1_15_0_0_t0b; // @[Map2T.scala 8:20]
  wire  op_I1_15_0_0_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_8_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_9_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_10_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_11_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_12_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_13_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_14_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_0_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_0_t1b_t0b; // @[Map2T.scala 8:20]
  wire [31:0] op_O_15_0_0_t1b_t1b; // @[Map2T.scala 8:20]
  Map2S_53 op ( // @[Map2T.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_0_2_0(op_I0_0_2_0),
    .I0_0_2_1(op_I0_0_2_1),
    .I0_0_2_2(op_I0_0_2_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_1_2_0(op_I0_1_2_0),
    .I0_1_2_1(op_I0_1_2_1),
    .I0_1_2_2(op_I0_1_2_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_2_2_0(op_I0_2_2_0),
    .I0_2_2_1(op_I0_2_2_1),
    .I0_2_2_2(op_I0_2_2_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_3_2_0(op_I0_3_2_0),
    .I0_3_2_1(op_I0_3_2_1),
    .I0_3_2_2(op_I0_3_2_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_4_2_0(op_I0_4_2_0),
    .I0_4_2_1(op_I0_4_2_1),
    .I0_4_2_2(op_I0_4_2_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_5_2_0(op_I0_5_2_0),
    .I0_5_2_1(op_I0_5_2_1),
    .I0_5_2_2(op_I0_5_2_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_6_2_0(op_I0_6_2_0),
    .I0_6_2_1(op_I0_6_2_1),
    .I0_6_2_2(op_I0_6_2_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I0_7_2_0(op_I0_7_2_0),
    .I0_7_2_1(op_I0_7_2_1),
    .I0_7_2_2(op_I0_7_2_2),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_8_0_1(op_I0_8_0_1),
    .I0_8_0_2(op_I0_8_0_2),
    .I0_8_1_0(op_I0_8_1_0),
    .I0_8_1_1(op_I0_8_1_1),
    .I0_8_1_2(op_I0_8_1_2),
    .I0_8_2_0(op_I0_8_2_0),
    .I0_8_2_1(op_I0_8_2_1),
    .I0_8_2_2(op_I0_8_2_2),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_9_0_1(op_I0_9_0_1),
    .I0_9_0_2(op_I0_9_0_2),
    .I0_9_1_0(op_I0_9_1_0),
    .I0_9_1_1(op_I0_9_1_1),
    .I0_9_1_2(op_I0_9_1_2),
    .I0_9_2_0(op_I0_9_2_0),
    .I0_9_2_1(op_I0_9_2_1),
    .I0_9_2_2(op_I0_9_2_2),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_10_0_1(op_I0_10_0_1),
    .I0_10_0_2(op_I0_10_0_2),
    .I0_10_1_0(op_I0_10_1_0),
    .I0_10_1_1(op_I0_10_1_1),
    .I0_10_1_2(op_I0_10_1_2),
    .I0_10_2_0(op_I0_10_2_0),
    .I0_10_2_1(op_I0_10_2_1),
    .I0_10_2_2(op_I0_10_2_2),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_11_0_1(op_I0_11_0_1),
    .I0_11_0_2(op_I0_11_0_2),
    .I0_11_1_0(op_I0_11_1_0),
    .I0_11_1_1(op_I0_11_1_1),
    .I0_11_1_2(op_I0_11_1_2),
    .I0_11_2_0(op_I0_11_2_0),
    .I0_11_2_1(op_I0_11_2_1),
    .I0_11_2_2(op_I0_11_2_2),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_12_0_1(op_I0_12_0_1),
    .I0_12_0_2(op_I0_12_0_2),
    .I0_12_1_0(op_I0_12_1_0),
    .I0_12_1_1(op_I0_12_1_1),
    .I0_12_1_2(op_I0_12_1_2),
    .I0_12_2_0(op_I0_12_2_0),
    .I0_12_2_1(op_I0_12_2_1),
    .I0_12_2_2(op_I0_12_2_2),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_13_0_1(op_I0_13_0_1),
    .I0_13_0_2(op_I0_13_0_2),
    .I0_13_1_0(op_I0_13_1_0),
    .I0_13_1_1(op_I0_13_1_1),
    .I0_13_1_2(op_I0_13_1_2),
    .I0_13_2_0(op_I0_13_2_0),
    .I0_13_2_1(op_I0_13_2_1),
    .I0_13_2_2(op_I0_13_2_2),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_14_0_1(op_I0_14_0_1),
    .I0_14_0_2(op_I0_14_0_2),
    .I0_14_1_0(op_I0_14_1_0),
    .I0_14_1_1(op_I0_14_1_1),
    .I0_14_1_2(op_I0_14_1_2),
    .I0_14_2_0(op_I0_14_2_0),
    .I0_14_2_1(op_I0_14_2_1),
    .I0_14_2_2(op_I0_14_2_2),
    .I0_15_0_0(op_I0_15_0_0),
    .I0_15_0_1(op_I0_15_0_1),
    .I0_15_0_2(op_I0_15_0_2),
    .I0_15_1_0(op_I0_15_1_0),
    .I0_15_1_1(op_I0_15_1_1),
    .I0_15_1_2(op_I0_15_1_2),
    .I0_15_2_0(op_I0_15_2_0),
    .I0_15_2_1(op_I0_15_2_1),
    .I0_15_2_2(op_I0_15_2_2),
    .I1_0_0_0_t0b(op_I1_0_0_0_t0b),
    .I1_0_0_0_t1b(op_I1_0_0_0_t1b),
    .I1_1_0_0_t0b(op_I1_1_0_0_t0b),
    .I1_1_0_0_t1b(op_I1_1_0_0_t1b),
    .I1_2_0_0_t0b(op_I1_2_0_0_t0b),
    .I1_2_0_0_t1b(op_I1_2_0_0_t1b),
    .I1_3_0_0_t0b(op_I1_3_0_0_t0b),
    .I1_3_0_0_t1b(op_I1_3_0_0_t1b),
    .I1_4_0_0_t0b(op_I1_4_0_0_t0b),
    .I1_4_0_0_t1b(op_I1_4_0_0_t1b),
    .I1_5_0_0_t0b(op_I1_5_0_0_t0b),
    .I1_5_0_0_t1b(op_I1_5_0_0_t1b),
    .I1_6_0_0_t0b(op_I1_6_0_0_t0b),
    .I1_6_0_0_t1b(op_I1_6_0_0_t1b),
    .I1_7_0_0_t0b(op_I1_7_0_0_t0b),
    .I1_7_0_0_t1b(op_I1_7_0_0_t1b),
    .I1_8_0_0_t0b(op_I1_8_0_0_t0b),
    .I1_8_0_0_t1b(op_I1_8_0_0_t1b),
    .I1_9_0_0_t0b(op_I1_9_0_0_t0b),
    .I1_9_0_0_t1b(op_I1_9_0_0_t1b),
    .I1_10_0_0_t0b(op_I1_10_0_0_t0b),
    .I1_10_0_0_t1b(op_I1_10_0_0_t1b),
    .I1_11_0_0_t0b(op_I1_11_0_0_t0b),
    .I1_11_0_0_t1b(op_I1_11_0_0_t1b),
    .I1_12_0_0_t0b(op_I1_12_0_0_t0b),
    .I1_12_0_0_t1b(op_I1_12_0_0_t1b),
    .I1_13_0_0_t0b(op_I1_13_0_0_t0b),
    .I1_13_0_0_t1b(op_I1_13_0_0_t1b),
    .I1_14_0_0_t0b(op_I1_14_0_0_t0b),
    .I1_14_0_0_t1b(op_I1_14_0_0_t1b),
    .I1_15_0_0_t0b(op_I1_15_0_0_t0b),
    .I1_15_0_0_t1b(op_I1_15_0_0_t1b),
    .O_0_0_0_t0b(op_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(op_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(op_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(op_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(op_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(op_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(op_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(op_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(op_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(op_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(op_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(op_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(op_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(op_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(op_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(op_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(op_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(op_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(op_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(op_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(op_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(op_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(op_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(op_O_7_0_0_t1b_t1b),
    .O_8_0_0_t0b(op_O_8_0_0_t0b),
    .O_8_0_0_t1b_t0b(op_O_8_0_0_t1b_t0b),
    .O_8_0_0_t1b_t1b(op_O_8_0_0_t1b_t1b),
    .O_9_0_0_t0b(op_O_9_0_0_t0b),
    .O_9_0_0_t1b_t0b(op_O_9_0_0_t1b_t0b),
    .O_9_0_0_t1b_t1b(op_O_9_0_0_t1b_t1b),
    .O_10_0_0_t0b(op_O_10_0_0_t0b),
    .O_10_0_0_t1b_t0b(op_O_10_0_0_t1b_t0b),
    .O_10_0_0_t1b_t1b(op_O_10_0_0_t1b_t1b),
    .O_11_0_0_t0b(op_O_11_0_0_t0b),
    .O_11_0_0_t1b_t0b(op_O_11_0_0_t1b_t0b),
    .O_11_0_0_t1b_t1b(op_O_11_0_0_t1b_t1b),
    .O_12_0_0_t0b(op_O_12_0_0_t0b),
    .O_12_0_0_t1b_t0b(op_O_12_0_0_t1b_t0b),
    .O_12_0_0_t1b_t1b(op_O_12_0_0_t1b_t1b),
    .O_13_0_0_t0b(op_O_13_0_0_t0b),
    .O_13_0_0_t1b_t0b(op_O_13_0_0_t1b_t0b),
    .O_13_0_0_t1b_t1b(op_O_13_0_0_t1b_t1b),
    .O_14_0_0_t0b(op_O_14_0_0_t0b),
    .O_14_0_0_t1b_t0b(op_O_14_0_0_t1b_t0b),
    .O_14_0_0_t1b_t1b(op_O_14_0_0_t1b_t1b),
    .O_15_0_0_t0b(op_O_15_0_0_t0b),
    .O_15_0_0_t1b_t0b(op_O_15_0_0_t1b_t0b),
    .O_15_0_0_t1b_t1b(op_O_15_0_0_t1b_t1b)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0_t0b = op_O_0_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_0_0_0_t1b_t0b = op_O_0_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_0_0_0_t1b_t1b = op_O_0_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_1_0_0_t0b = op_O_1_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_1_0_0_t1b_t0b = op_O_1_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_1_0_0_t1b_t1b = op_O_1_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_2_0_0_t0b = op_O_2_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_2_0_0_t1b_t0b = op_O_2_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_2_0_0_t1b_t1b = op_O_2_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_3_0_0_t0b = op_O_3_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_3_0_0_t1b_t0b = op_O_3_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_3_0_0_t1b_t1b = op_O_3_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_4_0_0_t0b = op_O_4_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_4_0_0_t1b_t0b = op_O_4_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_4_0_0_t1b_t1b = op_O_4_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_5_0_0_t0b = op_O_5_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_5_0_0_t1b_t0b = op_O_5_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_5_0_0_t1b_t1b = op_O_5_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_6_0_0_t0b = op_O_6_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_6_0_0_t1b_t0b = op_O_6_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_6_0_0_t1b_t1b = op_O_6_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_7_0_0_t0b = op_O_7_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_7_0_0_t1b_t0b = op_O_7_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_7_0_0_t1b_t1b = op_O_7_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_8_0_0_t0b = op_O_8_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_8_0_0_t1b_t0b = op_O_8_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_8_0_0_t1b_t1b = op_O_8_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_9_0_0_t0b = op_O_9_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_9_0_0_t1b_t0b = op_O_9_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_9_0_0_t1b_t1b = op_O_9_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_10_0_0_t0b = op_O_10_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_10_0_0_t1b_t0b = op_O_10_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_10_0_0_t1b_t1b = op_O_10_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_11_0_0_t0b = op_O_11_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_11_0_0_t1b_t0b = op_O_11_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_11_0_0_t1b_t1b = op_O_11_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_12_0_0_t0b = op_O_12_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_12_0_0_t1b_t0b = op_O_12_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_12_0_0_t1b_t1b = op_O_12_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_13_0_0_t0b = op_O_13_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_13_0_0_t1b_t0b = op_O_13_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_13_0_0_t1b_t1b = op_O_13_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_14_0_0_t0b = op_O_14_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_14_0_0_t1b_t0b = op_O_14_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_14_0_0_t1b_t1b = op_O_14_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign O_15_0_0_t0b = op_O_15_0_0_t0b; // @[Map2T.scala 17:7]
  assign O_15_0_0_t1b_t0b = op_O_15_0_0_t1b_t0b; // @[Map2T.scala 17:7]
  assign O_15_0_0_t1b_t1b = op_O_15_0_0_t1b_t1b; // @[Map2T.scala 17:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_0_2_0 = I0_0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_0_2_1 = I0_0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2_2 = I0_0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_2_0 = I0_1_2_0; // @[Map2T.scala 15:11]
  assign op_I0_1_2_1 = I0_1_2_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2_2 = I0_1_2_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_2_0 = I0_2_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_2_1 = I0_2_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2_2 = I0_2_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_2_0 = I0_3_2_0; // @[Map2T.scala 15:11]
  assign op_I0_3_2_1 = I0_3_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2_2 = I0_3_2_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_2_0 = I0_4_2_0; // @[Map2T.scala 15:11]
  assign op_I0_4_2_1 = I0_4_2_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2_2 = I0_4_2_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_2_0 = I0_5_2_0; // @[Map2T.scala 15:11]
  assign op_I0_5_2_1 = I0_5_2_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2_2 = I0_5_2_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_2_0 = I0_6_2_0; // @[Map2T.scala 15:11]
  assign op_I0_6_2_1 = I0_6_2_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2_2 = I0_6_2_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_2_0 = I0_7_2_0; // @[Map2T.scala 15:11]
  assign op_I0_7_2_1 = I0_7_2_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2_2 = I0_7_2_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1 = I0_8_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_2 = I0_8_0_2; // @[Map2T.scala 15:11]
  assign op_I0_8_1_0 = I0_8_1_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1_1 = I0_8_1_1; // @[Map2T.scala 15:11]
  assign op_I0_8_1_2 = I0_8_1_2; // @[Map2T.scala 15:11]
  assign op_I0_8_2_0 = I0_8_2_0; // @[Map2T.scala 15:11]
  assign op_I0_8_2_1 = I0_8_2_1; // @[Map2T.scala 15:11]
  assign op_I0_8_2_2 = I0_8_2_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1 = I0_9_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_2 = I0_9_0_2; // @[Map2T.scala 15:11]
  assign op_I0_9_1_0 = I0_9_1_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1_1 = I0_9_1_1; // @[Map2T.scala 15:11]
  assign op_I0_9_1_2 = I0_9_1_2; // @[Map2T.scala 15:11]
  assign op_I0_9_2_0 = I0_9_2_0; // @[Map2T.scala 15:11]
  assign op_I0_9_2_1 = I0_9_2_1; // @[Map2T.scala 15:11]
  assign op_I0_9_2_2 = I0_9_2_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1 = I0_10_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_2 = I0_10_0_2; // @[Map2T.scala 15:11]
  assign op_I0_10_1_0 = I0_10_1_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1_1 = I0_10_1_1; // @[Map2T.scala 15:11]
  assign op_I0_10_1_2 = I0_10_1_2; // @[Map2T.scala 15:11]
  assign op_I0_10_2_0 = I0_10_2_0; // @[Map2T.scala 15:11]
  assign op_I0_10_2_1 = I0_10_2_1; // @[Map2T.scala 15:11]
  assign op_I0_10_2_2 = I0_10_2_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1 = I0_11_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_2 = I0_11_0_2; // @[Map2T.scala 15:11]
  assign op_I0_11_1_0 = I0_11_1_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1_1 = I0_11_1_1; // @[Map2T.scala 15:11]
  assign op_I0_11_1_2 = I0_11_1_2; // @[Map2T.scala 15:11]
  assign op_I0_11_2_0 = I0_11_2_0; // @[Map2T.scala 15:11]
  assign op_I0_11_2_1 = I0_11_2_1; // @[Map2T.scala 15:11]
  assign op_I0_11_2_2 = I0_11_2_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1 = I0_12_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_2 = I0_12_0_2; // @[Map2T.scala 15:11]
  assign op_I0_12_1_0 = I0_12_1_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1_1 = I0_12_1_1; // @[Map2T.scala 15:11]
  assign op_I0_12_1_2 = I0_12_1_2; // @[Map2T.scala 15:11]
  assign op_I0_12_2_0 = I0_12_2_0; // @[Map2T.scala 15:11]
  assign op_I0_12_2_1 = I0_12_2_1; // @[Map2T.scala 15:11]
  assign op_I0_12_2_2 = I0_12_2_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1 = I0_13_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_2 = I0_13_0_2; // @[Map2T.scala 15:11]
  assign op_I0_13_1_0 = I0_13_1_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1_1 = I0_13_1_1; // @[Map2T.scala 15:11]
  assign op_I0_13_1_2 = I0_13_1_2; // @[Map2T.scala 15:11]
  assign op_I0_13_2_0 = I0_13_2_0; // @[Map2T.scala 15:11]
  assign op_I0_13_2_1 = I0_13_2_1; // @[Map2T.scala 15:11]
  assign op_I0_13_2_2 = I0_13_2_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1 = I0_14_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_2 = I0_14_0_2; // @[Map2T.scala 15:11]
  assign op_I0_14_1_0 = I0_14_1_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1_1 = I0_14_1_1; // @[Map2T.scala 15:11]
  assign op_I0_14_1_2 = I0_14_1_2; // @[Map2T.scala 15:11]
  assign op_I0_14_2_0 = I0_14_2_0; // @[Map2T.scala 15:11]
  assign op_I0_14_2_1 = I0_14_2_1; // @[Map2T.scala 15:11]
  assign op_I0_14_2_2 = I0_14_2_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1 = I0_15_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_2 = I0_15_0_2; // @[Map2T.scala 15:11]
  assign op_I0_15_1_0 = I0_15_1_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1_1 = I0_15_1_1; // @[Map2T.scala 15:11]
  assign op_I0_15_1_2 = I0_15_1_2; // @[Map2T.scala 15:11]
  assign op_I0_15_2_0 = I0_15_2_0; // @[Map2T.scala 15:11]
  assign op_I0_15_2_1 = I0_15_2_1; // @[Map2T.scala 15:11]
  assign op_I0_15_2_2 = I0_15_2_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0_0_t0b = I1_0_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_0_0_0_t1b = I1_0_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0_t0b = I1_1_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_1_0_0_t1b = I1_1_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0_t0b = I1_2_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_2_0_0_t1b = I1_2_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0_t0b = I1_3_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_3_0_0_t1b = I1_3_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0_t0b = I1_4_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_4_0_0_t1b = I1_4_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0_t0b = I1_5_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_5_0_0_t1b = I1_5_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0_t0b = I1_6_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_6_0_0_t1b = I1_6_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0_t0b = I1_7_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_7_0_0_t1b = I1_7_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0_t0b = I1_8_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_8_0_0_t1b = I1_8_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0_t0b = I1_9_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_9_0_0_t1b = I1_9_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0_t0b = I1_10_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_10_0_0_t1b = I1_10_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0_t0b = I1_11_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_11_0_0_t1b = I1_11_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0_t0b = I1_12_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_12_0_0_t1b = I1_12_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0_t0b = I1_13_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_13_0_0_t1b = I1_13_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0_t0b = I1_14_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_14_0_0_t1b = I1_14_0_0_t1b; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0_t0b = I1_15_0_0_t0b; // @[Map2T.scala 16:11]
  assign op_I1_15_0_0_t1b = I1_15_0_0_t1b; // @[Map2T.scala 16:11]
endmodule
module Module_7(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_8_1_0,
  input  [31:0] I_8_1_1,
  input  [31:0] I_8_1_2,
  input  [31:0] I_8_2_0,
  input  [31:0] I_8_2_1,
  input  [31:0] I_8_2_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_9_1_0,
  input  [31:0] I_9_1_1,
  input  [31:0] I_9_1_2,
  input  [31:0] I_9_2_0,
  input  [31:0] I_9_2_1,
  input  [31:0] I_9_2_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_10_1_0,
  input  [31:0] I_10_1_1,
  input  [31:0] I_10_1_2,
  input  [31:0] I_10_2_0,
  input  [31:0] I_10_2_1,
  input  [31:0] I_10_2_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_11_1_0,
  input  [31:0] I_11_1_1,
  input  [31:0] I_11_1_2,
  input  [31:0] I_11_2_0,
  input  [31:0] I_11_2_1,
  input  [31:0] I_11_2_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_12_1_0,
  input  [31:0] I_12_1_1,
  input  [31:0] I_12_1_2,
  input  [31:0] I_12_2_0,
  input  [31:0] I_12_2_1,
  input  [31:0] I_12_2_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_13_1_0,
  input  [31:0] I_13_1_1,
  input  [31:0] I_13_1_2,
  input  [31:0] I_13_2_0,
  input  [31:0] I_13_2_1,
  input  [31:0] I_13_2_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_14_1_0,
  input  [31:0] I_14_1_1,
  input  [31:0] I_14_1_2,
  input  [31:0] I_14_2_0,
  input  [31:0] I_14_2_1,
  input  [31:0] I_14_2_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  input  [31:0] I_15_1_0,
  input  [31:0] I_15_1_1,
  input  [31:0] I_15_1_2,
  input  [31:0] I_15_2_0,
  input  [31:0] I_15_2_1,
  input  [31:0] I_15_2_2,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b,
  output [31:0] O_8_0_0_t0b,
  output [31:0] O_8_0_0_t1b_t0b,
  output [31:0] O_8_0_0_t1b_t1b,
  output [31:0] O_9_0_0_t0b,
  output [31:0] O_9_0_0_t1b_t0b,
  output [31:0] O_9_0_0_t1b_t1b,
  output [31:0] O_10_0_0_t0b,
  output [31:0] O_10_0_0_t1b_t0b,
  output [31:0] O_10_0_0_t1b_t1b,
  output [31:0] O_11_0_0_t0b,
  output [31:0] O_11_0_0_t1b_t0b,
  output [31:0] O_11_0_0_t1b_t1b,
  output [31:0] O_12_0_0_t0b,
  output [31:0] O_12_0_0_t1b_t0b,
  output [31:0] O_12_0_0_t1b_t1b,
  output [31:0] O_13_0_0_t0b,
  output [31:0] O_13_0_0_t1b_t0b,
  output [31:0] O_13_0_0_t1b_t1b,
  output [31:0] O_14_0_0_t0b,
  output [31:0] O_14_0_0_t1b_t0b,
  output [31:0] O_14_0_0_t1b_t1b,
  output [31:0] O_15_0_0_t0b,
  output [31:0] O_15_0_0_t1b_t0b,
  output [31:0] O_15_0_0_t1b_t1b
);
  wire  counter108_clock; // @[Top.scala 325:28]
  wire  counter108_reset; // @[Top.scala 325:28]
  wire [31:0] counter108_O_0; // @[Top.scala 325:28]
  wire [31:0] counter108_O_1; // @[Top.scala 325:28]
  wire [31:0] counter108_O_2; // @[Top.scala 325:28]
  wire [31:0] counter108_O_3; // @[Top.scala 325:28]
  wire [31:0] counter108_O_4; // @[Top.scala 325:28]
  wire [31:0] counter108_O_5; // @[Top.scala 325:28]
  wire [31:0] counter108_O_6; // @[Top.scala 325:28]
  wire [31:0] counter108_O_7; // @[Top.scala 325:28]
  wire [31:0] counter108_O_8; // @[Top.scala 325:28]
  wire [31:0] counter108_O_9; // @[Top.scala 325:28]
  wire [31:0] counter108_O_10; // @[Top.scala 325:28]
  wire [31:0] counter108_O_11; // @[Top.scala 325:28]
  wire [31:0] counter108_O_12; // @[Top.scala 325:28]
  wire [31:0] counter108_O_13; // @[Top.scala 325:28]
  wire [31:0] counter108_O_14; // @[Top.scala 325:28]
  wire [31:0] counter108_O_15; // @[Top.scala 325:28]
  wire  n116_valid_down; // @[Top.scala 327:22]
  wire [31:0] n116_I_0; // @[Top.scala 327:22]
  wire [31:0] n116_I_1; // @[Top.scala 327:22]
  wire [31:0] n116_I_2; // @[Top.scala 327:22]
  wire [31:0] n116_I_3; // @[Top.scala 327:22]
  wire [31:0] n116_I_4; // @[Top.scala 327:22]
  wire [31:0] n116_I_5; // @[Top.scala 327:22]
  wire [31:0] n116_I_6; // @[Top.scala 327:22]
  wire [31:0] n116_I_7; // @[Top.scala 327:22]
  wire [31:0] n116_I_8; // @[Top.scala 327:22]
  wire [31:0] n116_I_9; // @[Top.scala 327:22]
  wire [31:0] n116_I_10; // @[Top.scala 327:22]
  wire [31:0] n116_I_11; // @[Top.scala 327:22]
  wire [31:0] n116_I_12; // @[Top.scala 327:22]
  wire [31:0] n116_I_13; // @[Top.scala 327:22]
  wire [31:0] n116_I_14; // @[Top.scala 327:22]
  wire [31:0] n116_I_15; // @[Top.scala 327:22]
  wire  n116_O_0; // @[Top.scala 327:22]
  wire  n116_O_1; // @[Top.scala 327:22]
  wire  n116_O_2; // @[Top.scala 327:22]
  wire  n116_O_3; // @[Top.scala 327:22]
  wire  n116_O_4; // @[Top.scala 327:22]
  wire  n116_O_5; // @[Top.scala 327:22]
  wire  n116_O_6; // @[Top.scala 327:22]
  wire  n116_O_7; // @[Top.scala 327:22]
  wire  n116_O_8; // @[Top.scala 327:22]
  wire  n116_O_9; // @[Top.scala 327:22]
  wire  n116_O_10; // @[Top.scala 327:22]
  wire  n116_O_11; // @[Top.scala 327:22]
  wire  n116_O_12; // @[Top.scala 327:22]
  wire  n116_O_13; // @[Top.scala 327:22]
  wire  n116_O_14; // @[Top.scala 327:22]
  wire  n116_O_15; // @[Top.scala 327:22]
  wire  n128_valid_down; // @[Top.scala 330:22]
  wire [31:0] n128_I_0; // @[Top.scala 330:22]
  wire [31:0] n128_I_1; // @[Top.scala 330:22]
  wire [31:0] n128_I_2; // @[Top.scala 330:22]
  wire [31:0] n128_I_3; // @[Top.scala 330:22]
  wire [31:0] n128_I_4; // @[Top.scala 330:22]
  wire [31:0] n128_I_5; // @[Top.scala 330:22]
  wire [31:0] n128_I_6; // @[Top.scala 330:22]
  wire [31:0] n128_I_7; // @[Top.scala 330:22]
  wire [31:0] n128_I_8; // @[Top.scala 330:22]
  wire [31:0] n128_I_9; // @[Top.scala 330:22]
  wire [31:0] n128_I_10; // @[Top.scala 330:22]
  wire [31:0] n128_I_11; // @[Top.scala 330:22]
  wire [31:0] n128_I_12; // @[Top.scala 330:22]
  wire [31:0] n128_I_13; // @[Top.scala 330:22]
  wire [31:0] n128_I_14; // @[Top.scala 330:22]
  wire [31:0] n128_I_15; // @[Top.scala 330:22]
  wire  n128_O_0; // @[Top.scala 330:22]
  wire  n128_O_1; // @[Top.scala 330:22]
  wire  n128_O_2; // @[Top.scala 330:22]
  wire  n128_O_3; // @[Top.scala 330:22]
  wire  n128_O_4; // @[Top.scala 330:22]
  wire  n128_O_5; // @[Top.scala 330:22]
  wire  n128_O_6; // @[Top.scala 330:22]
  wire  n128_O_7; // @[Top.scala 330:22]
  wire  n128_O_8; // @[Top.scala 330:22]
  wire  n128_O_9; // @[Top.scala 330:22]
  wire  n128_O_10; // @[Top.scala 330:22]
  wire  n128_O_11; // @[Top.scala 330:22]
  wire  n128_O_12; // @[Top.scala 330:22]
  wire  n128_O_13; // @[Top.scala 330:22]
  wire  n128_O_14; // @[Top.scala 330:22]
  wire  n128_O_15; // @[Top.scala 330:22]
  wire  n129_valid_up; // @[Top.scala 333:22]
  wire  n129_valid_down; // @[Top.scala 333:22]
  wire  n129_I0_0; // @[Top.scala 333:22]
  wire  n129_I0_1; // @[Top.scala 333:22]
  wire  n129_I0_2; // @[Top.scala 333:22]
  wire  n129_I0_3; // @[Top.scala 333:22]
  wire  n129_I0_4; // @[Top.scala 333:22]
  wire  n129_I0_5; // @[Top.scala 333:22]
  wire  n129_I0_6; // @[Top.scala 333:22]
  wire  n129_I0_7; // @[Top.scala 333:22]
  wire  n129_I0_8; // @[Top.scala 333:22]
  wire  n129_I0_9; // @[Top.scala 333:22]
  wire  n129_I0_10; // @[Top.scala 333:22]
  wire  n129_I0_11; // @[Top.scala 333:22]
  wire  n129_I0_12; // @[Top.scala 333:22]
  wire  n129_I0_13; // @[Top.scala 333:22]
  wire  n129_I0_14; // @[Top.scala 333:22]
  wire  n129_I0_15; // @[Top.scala 333:22]
  wire  n129_I1_0; // @[Top.scala 333:22]
  wire  n129_I1_1; // @[Top.scala 333:22]
  wire  n129_I1_2; // @[Top.scala 333:22]
  wire  n129_I1_3; // @[Top.scala 333:22]
  wire  n129_I1_4; // @[Top.scala 333:22]
  wire  n129_I1_5; // @[Top.scala 333:22]
  wire  n129_I1_6; // @[Top.scala 333:22]
  wire  n129_I1_7; // @[Top.scala 333:22]
  wire  n129_I1_8; // @[Top.scala 333:22]
  wire  n129_I1_9; // @[Top.scala 333:22]
  wire  n129_I1_10; // @[Top.scala 333:22]
  wire  n129_I1_11; // @[Top.scala 333:22]
  wire  n129_I1_12; // @[Top.scala 333:22]
  wire  n129_I1_13; // @[Top.scala 333:22]
  wire  n129_I1_14; // @[Top.scala 333:22]
  wire  n129_I1_15; // @[Top.scala 333:22]
  wire  n129_O_0_t0b; // @[Top.scala 333:22]
  wire  n129_O_0_t1b; // @[Top.scala 333:22]
  wire  n129_O_1_t0b; // @[Top.scala 333:22]
  wire  n129_O_1_t1b; // @[Top.scala 333:22]
  wire  n129_O_2_t0b; // @[Top.scala 333:22]
  wire  n129_O_2_t1b; // @[Top.scala 333:22]
  wire  n129_O_3_t0b; // @[Top.scala 333:22]
  wire  n129_O_3_t1b; // @[Top.scala 333:22]
  wire  n129_O_4_t0b; // @[Top.scala 333:22]
  wire  n129_O_4_t1b; // @[Top.scala 333:22]
  wire  n129_O_5_t0b; // @[Top.scala 333:22]
  wire  n129_O_5_t1b; // @[Top.scala 333:22]
  wire  n129_O_6_t0b; // @[Top.scala 333:22]
  wire  n129_O_6_t1b; // @[Top.scala 333:22]
  wire  n129_O_7_t0b; // @[Top.scala 333:22]
  wire  n129_O_7_t1b; // @[Top.scala 333:22]
  wire  n129_O_8_t0b; // @[Top.scala 333:22]
  wire  n129_O_8_t1b; // @[Top.scala 333:22]
  wire  n129_O_9_t0b; // @[Top.scala 333:22]
  wire  n129_O_9_t1b; // @[Top.scala 333:22]
  wire  n129_O_10_t0b; // @[Top.scala 333:22]
  wire  n129_O_10_t1b; // @[Top.scala 333:22]
  wire  n129_O_11_t0b; // @[Top.scala 333:22]
  wire  n129_O_11_t1b; // @[Top.scala 333:22]
  wire  n129_O_12_t0b; // @[Top.scala 333:22]
  wire  n129_O_12_t1b; // @[Top.scala 333:22]
  wire  n129_O_13_t0b; // @[Top.scala 333:22]
  wire  n129_O_13_t1b; // @[Top.scala 333:22]
  wire  n129_O_14_t0b; // @[Top.scala 333:22]
  wire  n129_O_14_t1b; // @[Top.scala 333:22]
  wire  n129_O_15_t0b; // @[Top.scala 333:22]
  wire  n129_O_15_t1b; // @[Top.scala 333:22]
  wire  n138_valid_up; // @[Top.scala 337:22]
  wire  n138_valid_down; // @[Top.scala 337:22]
  wire  n138_I_0_t0b; // @[Top.scala 337:22]
  wire  n138_I_0_t1b; // @[Top.scala 337:22]
  wire  n138_I_1_t0b; // @[Top.scala 337:22]
  wire  n138_I_1_t1b; // @[Top.scala 337:22]
  wire  n138_I_2_t0b; // @[Top.scala 337:22]
  wire  n138_I_2_t1b; // @[Top.scala 337:22]
  wire  n138_I_3_t0b; // @[Top.scala 337:22]
  wire  n138_I_3_t1b; // @[Top.scala 337:22]
  wire  n138_I_4_t0b; // @[Top.scala 337:22]
  wire  n138_I_4_t1b; // @[Top.scala 337:22]
  wire  n138_I_5_t0b; // @[Top.scala 337:22]
  wire  n138_I_5_t1b; // @[Top.scala 337:22]
  wire  n138_I_6_t0b; // @[Top.scala 337:22]
  wire  n138_I_6_t1b; // @[Top.scala 337:22]
  wire  n138_I_7_t0b; // @[Top.scala 337:22]
  wire  n138_I_7_t1b; // @[Top.scala 337:22]
  wire  n138_I_8_t0b; // @[Top.scala 337:22]
  wire  n138_I_8_t1b; // @[Top.scala 337:22]
  wire  n138_I_9_t0b; // @[Top.scala 337:22]
  wire  n138_I_9_t1b; // @[Top.scala 337:22]
  wire  n138_I_10_t0b; // @[Top.scala 337:22]
  wire  n138_I_10_t1b; // @[Top.scala 337:22]
  wire  n138_I_11_t0b; // @[Top.scala 337:22]
  wire  n138_I_11_t1b; // @[Top.scala 337:22]
  wire  n138_I_12_t0b; // @[Top.scala 337:22]
  wire  n138_I_12_t1b; // @[Top.scala 337:22]
  wire  n138_I_13_t0b; // @[Top.scala 337:22]
  wire  n138_I_13_t1b; // @[Top.scala 337:22]
  wire  n138_I_14_t0b; // @[Top.scala 337:22]
  wire  n138_I_14_t1b; // @[Top.scala 337:22]
  wire  n138_I_15_t0b; // @[Top.scala 337:22]
  wire  n138_I_15_t1b; // @[Top.scala 337:22]
  wire  n138_O_0_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_0_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_1_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_1_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_2_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_2_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_3_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_3_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_4_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_4_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_5_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_5_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_6_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_6_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_7_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_7_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_8_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_8_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_9_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_9_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_10_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_10_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_11_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_11_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_12_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_12_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_13_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_13_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_14_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_14_0_t1b; // @[Top.scala 337:22]
  wire  n138_O_15_0_t0b; // @[Top.scala 337:22]
  wire  n138_O_15_0_t1b; // @[Top.scala 337:22]
  wire  n141_valid_up; // @[Top.scala 340:22]
  wire  n141_valid_down; // @[Top.scala 340:22]
  wire  n141_I_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_1_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_1_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_2_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_2_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_3_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_3_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_4_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_4_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_5_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_5_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_6_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_6_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_7_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_7_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_8_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_8_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_9_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_9_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_10_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_10_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_11_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_11_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_12_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_12_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_13_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_13_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_14_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_14_0_t1b; // @[Top.scala 340:22]
  wire  n141_I_15_0_t0b; // @[Top.scala 340:22]
  wire  n141_I_15_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_0_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_0_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_1_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_1_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_2_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_2_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_3_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_3_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_4_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_4_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_5_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_5_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_6_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_6_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_7_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_7_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_8_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_8_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_9_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_9_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_10_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_10_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_11_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_11_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_12_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_12_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_13_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_13_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_14_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_14_0_0_t1b; // @[Top.scala 340:22]
  wire  n141_O_15_0_0_t0b; // @[Top.scala 340:22]
  wire  n141_O_15_0_0_t1b; // @[Top.scala 340:22]
  wire  n142_clock; // @[Top.scala 343:22]
  wire  n142_reset; // @[Top.scala 343:22]
  wire  n142_valid_up; // @[Top.scala 343:22]
  wire  n142_valid_down; // @[Top.scala 343:22]
  wire  n142_I_0_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_0_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_1_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_1_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_2_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_2_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_3_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_3_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_4_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_4_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_5_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_5_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_6_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_6_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_7_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_7_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_8_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_8_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_9_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_9_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_10_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_10_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_11_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_11_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_12_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_12_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_13_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_13_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_14_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_14_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_I_15_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_I_15_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_0_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_0_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_1_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_1_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_2_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_2_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_3_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_3_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_4_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_4_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_5_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_5_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_6_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_6_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_7_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_7_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_8_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_8_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_9_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_9_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_10_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_10_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_11_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_11_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_12_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_12_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_13_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_13_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_14_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_14_0_0_t1b; // @[Top.scala 343:22]
  wire  n142_O_15_0_0_t0b; // @[Top.scala 343:22]
  wire  n142_O_15_0_0_t1b; // @[Top.scala 343:22]
  wire  n143_clock; // @[Top.scala 346:22]
  wire  n143_reset; // @[Top.scala 346:22]
  wire  n143_valid_up; // @[Top.scala 346:22]
  wire  n143_valid_down; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_0_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_1_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_2_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_3_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_4_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_5_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_6_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_7_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_8_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_9_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_10_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_11_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_12_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_13_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_14_2_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_0_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_0_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_0_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_1_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_1_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_1_2; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_2_0; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_2_1; // @[Top.scala 346:22]
  wire [31:0] n143_I0_15_2_2; // @[Top.scala 346:22]
  wire  n143_I1_0_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_0_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_1_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_1_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_2_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_2_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_3_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_3_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_4_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_4_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_5_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_5_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_6_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_6_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_7_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_7_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_8_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_8_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_9_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_9_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_10_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_10_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_11_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_11_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_12_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_12_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_13_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_13_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_14_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_14_0_0_t1b; // @[Top.scala 346:22]
  wire  n143_I1_15_0_0_t0b; // @[Top.scala 346:22]
  wire  n143_I1_15_0_0_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_0_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_0_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_0_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_1_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_1_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_1_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_2_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_2_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_2_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_3_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_3_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_3_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_4_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_4_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_4_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_5_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_5_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_5_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_6_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_6_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_6_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_7_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_7_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_7_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_8_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_8_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_8_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_9_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_9_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_9_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_10_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_10_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_10_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_11_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_11_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_11_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_12_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_12_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_12_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_13_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_13_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_13_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_14_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_14_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_14_0_0_t1b_t1b; // @[Top.scala 346:22]
  wire [31:0] n143_O_15_0_0_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_15_0_0_t1b_t0b; // @[Top.scala 346:22]
  wire [31:0] n143_O_15_0_0_t1b_t1b; // @[Top.scala 346:22]
  Counter_TS counter108 ( // @[Top.scala 325:28]
    .clock(counter108_clock),
    .reset(counter108_reset),
    .O_0(counter108_O_0),
    .O_1(counter108_O_1),
    .O_2(counter108_O_2),
    .O_3(counter108_O_3),
    .O_4(counter108_O_4),
    .O_5(counter108_O_5),
    .O_6(counter108_O_6),
    .O_7(counter108_O_7),
    .O_8(counter108_O_8),
    .O_9(counter108_O_9),
    .O_10(counter108_O_10),
    .O_11(counter108_O_11),
    .O_12(counter108_O_12),
    .O_13(counter108_O_13),
    .O_14(counter108_O_14),
    .O_15(counter108_O_15)
  );
  MapT_8 n116 ( // @[Top.scala 327:22]
    .valid_down(n116_valid_down),
    .I_0(n116_I_0),
    .I_1(n116_I_1),
    .I_2(n116_I_2),
    .I_3(n116_I_3),
    .I_4(n116_I_4),
    .I_5(n116_I_5),
    .I_6(n116_I_6),
    .I_7(n116_I_7),
    .I_8(n116_I_8),
    .I_9(n116_I_9),
    .I_10(n116_I_10),
    .I_11(n116_I_11),
    .I_12(n116_I_12),
    .I_13(n116_I_13),
    .I_14(n116_I_14),
    .I_15(n116_I_15),
    .O_0(n116_O_0),
    .O_1(n116_O_1),
    .O_2(n116_O_2),
    .O_3(n116_O_3),
    .O_4(n116_O_4),
    .O_5(n116_O_5),
    .O_6(n116_O_6),
    .O_7(n116_O_7),
    .O_8(n116_O_8),
    .O_9(n116_O_9),
    .O_10(n116_O_10),
    .O_11(n116_O_11),
    .O_12(n116_O_12),
    .O_13(n116_O_13),
    .O_14(n116_O_14),
    .O_15(n116_O_15)
  );
  MapT_9 n128 ( // @[Top.scala 330:22]
    .valid_down(n128_valid_down),
    .I_0(n128_I_0),
    .I_1(n128_I_1),
    .I_2(n128_I_2),
    .I_3(n128_I_3),
    .I_4(n128_I_4),
    .I_5(n128_I_5),
    .I_6(n128_I_6),
    .I_7(n128_I_7),
    .I_8(n128_I_8),
    .I_9(n128_I_9),
    .I_10(n128_I_10),
    .I_11(n128_I_11),
    .I_12(n128_I_12),
    .I_13(n128_I_13),
    .I_14(n128_I_14),
    .I_15(n128_I_15),
    .O_0(n128_O_0),
    .O_1(n128_O_1),
    .O_2(n128_O_2),
    .O_3(n128_O_3),
    .O_4(n128_O_4),
    .O_5(n128_O_5),
    .O_6(n128_O_6),
    .O_7(n128_O_7),
    .O_8(n128_O_8),
    .O_9(n128_O_9),
    .O_10(n128_O_10),
    .O_11(n128_O_11),
    .O_12(n128_O_12),
    .O_13(n128_O_13),
    .O_14(n128_O_14),
    .O_15(n128_O_15)
  );
  Map2T_8 n129 ( // @[Top.scala 333:22]
    .valid_up(n129_valid_up),
    .valid_down(n129_valid_down),
    .I0_0(n129_I0_0),
    .I0_1(n129_I0_1),
    .I0_2(n129_I0_2),
    .I0_3(n129_I0_3),
    .I0_4(n129_I0_4),
    .I0_5(n129_I0_5),
    .I0_6(n129_I0_6),
    .I0_7(n129_I0_7),
    .I0_8(n129_I0_8),
    .I0_9(n129_I0_9),
    .I0_10(n129_I0_10),
    .I0_11(n129_I0_11),
    .I0_12(n129_I0_12),
    .I0_13(n129_I0_13),
    .I0_14(n129_I0_14),
    .I0_15(n129_I0_15),
    .I1_0(n129_I1_0),
    .I1_1(n129_I1_1),
    .I1_2(n129_I1_2),
    .I1_3(n129_I1_3),
    .I1_4(n129_I1_4),
    .I1_5(n129_I1_5),
    .I1_6(n129_I1_6),
    .I1_7(n129_I1_7),
    .I1_8(n129_I1_8),
    .I1_9(n129_I1_9),
    .I1_10(n129_I1_10),
    .I1_11(n129_I1_11),
    .I1_12(n129_I1_12),
    .I1_13(n129_I1_13),
    .I1_14(n129_I1_14),
    .I1_15(n129_I1_15),
    .O_0_t0b(n129_O_0_t0b),
    .O_0_t1b(n129_O_0_t1b),
    .O_1_t0b(n129_O_1_t0b),
    .O_1_t1b(n129_O_1_t1b),
    .O_2_t0b(n129_O_2_t0b),
    .O_2_t1b(n129_O_2_t1b),
    .O_3_t0b(n129_O_3_t0b),
    .O_3_t1b(n129_O_3_t1b),
    .O_4_t0b(n129_O_4_t0b),
    .O_4_t1b(n129_O_4_t1b),
    .O_5_t0b(n129_O_5_t0b),
    .O_5_t1b(n129_O_5_t1b),
    .O_6_t0b(n129_O_6_t0b),
    .O_6_t1b(n129_O_6_t1b),
    .O_7_t0b(n129_O_7_t0b),
    .O_7_t1b(n129_O_7_t1b),
    .O_8_t0b(n129_O_8_t0b),
    .O_8_t1b(n129_O_8_t1b),
    .O_9_t0b(n129_O_9_t0b),
    .O_9_t1b(n129_O_9_t1b),
    .O_10_t0b(n129_O_10_t0b),
    .O_10_t1b(n129_O_10_t1b),
    .O_11_t0b(n129_O_11_t0b),
    .O_11_t1b(n129_O_11_t1b),
    .O_12_t0b(n129_O_12_t0b),
    .O_12_t1b(n129_O_12_t1b),
    .O_13_t0b(n129_O_13_t0b),
    .O_13_t1b(n129_O_13_t1b),
    .O_14_t0b(n129_O_14_t0b),
    .O_14_t1b(n129_O_14_t1b),
    .O_15_t0b(n129_O_15_t0b),
    .O_15_t1b(n129_O_15_t1b)
  );
  MapT_10 n138 ( // @[Top.scala 337:22]
    .valid_up(n138_valid_up),
    .valid_down(n138_valid_down),
    .I_0_t0b(n138_I_0_t0b),
    .I_0_t1b(n138_I_0_t1b),
    .I_1_t0b(n138_I_1_t0b),
    .I_1_t1b(n138_I_1_t1b),
    .I_2_t0b(n138_I_2_t0b),
    .I_2_t1b(n138_I_2_t1b),
    .I_3_t0b(n138_I_3_t0b),
    .I_3_t1b(n138_I_3_t1b),
    .I_4_t0b(n138_I_4_t0b),
    .I_4_t1b(n138_I_4_t1b),
    .I_5_t0b(n138_I_5_t0b),
    .I_5_t1b(n138_I_5_t1b),
    .I_6_t0b(n138_I_6_t0b),
    .I_6_t1b(n138_I_6_t1b),
    .I_7_t0b(n138_I_7_t0b),
    .I_7_t1b(n138_I_7_t1b),
    .I_8_t0b(n138_I_8_t0b),
    .I_8_t1b(n138_I_8_t1b),
    .I_9_t0b(n138_I_9_t0b),
    .I_9_t1b(n138_I_9_t1b),
    .I_10_t0b(n138_I_10_t0b),
    .I_10_t1b(n138_I_10_t1b),
    .I_11_t0b(n138_I_11_t0b),
    .I_11_t1b(n138_I_11_t1b),
    .I_12_t0b(n138_I_12_t0b),
    .I_12_t1b(n138_I_12_t1b),
    .I_13_t0b(n138_I_13_t0b),
    .I_13_t1b(n138_I_13_t1b),
    .I_14_t0b(n138_I_14_t0b),
    .I_14_t1b(n138_I_14_t1b),
    .I_15_t0b(n138_I_15_t0b),
    .I_15_t1b(n138_I_15_t1b),
    .O_0_0_t0b(n138_O_0_0_t0b),
    .O_0_0_t1b(n138_O_0_0_t1b),
    .O_1_0_t0b(n138_O_1_0_t0b),
    .O_1_0_t1b(n138_O_1_0_t1b),
    .O_2_0_t0b(n138_O_2_0_t0b),
    .O_2_0_t1b(n138_O_2_0_t1b),
    .O_3_0_t0b(n138_O_3_0_t0b),
    .O_3_0_t1b(n138_O_3_0_t1b),
    .O_4_0_t0b(n138_O_4_0_t0b),
    .O_4_0_t1b(n138_O_4_0_t1b),
    .O_5_0_t0b(n138_O_5_0_t0b),
    .O_5_0_t1b(n138_O_5_0_t1b),
    .O_6_0_t0b(n138_O_6_0_t0b),
    .O_6_0_t1b(n138_O_6_0_t1b),
    .O_7_0_t0b(n138_O_7_0_t0b),
    .O_7_0_t1b(n138_O_7_0_t1b),
    .O_8_0_t0b(n138_O_8_0_t0b),
    .O_8_0_t1b(n138_O_8_0_t1b),
    .O_9_0_t0b(n138_O_9_0_t0b),
    .O_9_0_t1b(n138_O_9_0_t1b),
    .O_10_0_t0b(n138_O_10_0_t0b),
    .O_10_0_t1b(n138_O_10_0_t1b),
    .O_11_0_t0b(n138_O_11_0_t0b),
    .O_11_0_t1b(n138_O_11_0_t1b),
    .O_12_0_t0b(n138_O_12_0_t0b),
    .O_12_0_t1b(n138_O_12_0_t1b),
    .O_13_0_t0b(n138_O_13_0_t0b),
    .O_13_0_t1b(n138_O_13_0_t1b),
    .O_14_0_t0b(n138_O_14_0_t0b),
    .O_14_0_t1b(n138_O_14_0_t1b),
    .O_15_0_t0b(n138_O_15_0_t0b),
    .O_15_0_t1b(n138_O_15_0_t1b)
  );
  MapT_11 n141 ( // @[Top.scala 340:22]
    .valid_up(n141_valid_up),
    .valid_down(n141_valid_down),
    .I_0_0_t0b(n141_I_0_0_t0b),
    .I_0_0_t1b(n141_I_0_0_t1b),
    .I_1_0_t0b(n141_I_1_0_t0b),
    .I_1_0_t1b(n141_I_1_0_t1b),
    .I_2_0_t0b(n141_I_2_0_t0b),
    .I_2_0_t1b(n141_I_2_0_t1b),
    .I_3_0_t0b(n141_I_3_0_t0b),
    .I_3_0_t1b(n141_I_3_0_t1b),
    .I_4_0_t0b(n141_I_4_0_t0b),
    .I_4_0_t1b(n141_I_4_0_t1b),
    .I_5_0_t0b(n141_I_5_0_t0b),
    .I_5_0_t1b(n141_I_5_0_t1b),
    .I_6_0_t0b(n141_I_6_0_t0b),
    .I_6_0_t1b(n141_I_6_0_t1b),
    .I_7_0_t0b(n141_I_7_0_t0b),
    .I_7_0_t1b(n141_I_7_0_t1b),
    .I_8_0_t0b(n141_I_8_0_t0b),
    .I_8_0_t1b(n141_I_8_0_t1b),
    .I_9_0_t0b(n141_I_9_0_t0b),
    .I_9_0_t1b(n141_I_9_0_t1b),
    .I_10_0_t0b(n141_I_10_0_t0b),
    .I_10_0_t1b(n141_I_10_0_t1b),
    .I_11_0_t0b(n141_I_11_0_t0b),
    .I_11_0_t1b(n141_I_11_0_t1b),
    .I_12_0_t0b(n141_I_12_0_t0b),
    .I_12_0_t1b(n141_I_12_0_t1b),
    .I_13_0_t0b(n141_I_13_0_t0b),
    .I_13_0_t1b(n141_I_13_0_t1b),
    .I_14_0_t0b(n141_I_14_0_t0b),
    .I_14_0_t1b(n141_I_14_0_t1b),
    .I_15_0_t0b(n141_I_15_0_t0b),
    .I_15_0_t1b(n141_I_15_0_t1b),
    .O_0_0_0_t0b(n141_O_0_0_0_t0b),
    .O_0_0_0_t1b(n141_O_0_0_0_t1b),
    .O_1_0_0_t0b(n141_O_1_0_0_t0b),
    .O_1_0_0_t1b(n141_O_1_0_0_t1b),
    .O_2_0_0_t0b(n141_O_2_0_0_t0b),
    .O_2_0_0_t1b(n141_O_2_0_0_t1b),
    .O_3_0_0_t0b(n141_O_3_0_0_t0b),
    .O_3_0_0_t1b(n141_O_3_0_0_t1b),
    .O_4_0_0_t0b(n141_O_4_0_0_t0b),
    .O_4_0_0_t1b(n141_O_4_0_0_t1b),
    .O_5_0_0_t0b(n141_O_5_0_0_t0b),
    .O_5_0_0_t1b(n141_O_5_0_0_t1b),
    .O_6_0_0_t0b(n141_O_6_0_0_t0b),
    .O_6_0_0_t1b(n141_O_6_0_0_t1b),
    .O_7_0_0_t0b(n141_O_7_0_0_t0b),
    .O_7_0_0_t1b(n141_O_7_0_0_t1b),
    .O_8_0_0_t0b(n141_O_8_0_0_t0b),
    .O_8_0_0_t1b(n141_O_8_0_0_t1b),
    .O_9_0_0_t0b(n141_O_9_0_0_t0b),
    .O_9_0_0_t1b(n141_O_9_0_0_t1b),
    .O_10_0_0_t0b(n141_O_10_0_0_t0b),
    .O_10_0_0_t1b(n141_O_10_0_0_t1b),
    .O_11_0_0_t0b(n141_O_11_0_0_t0b),
    .O_11_0_0_t1b(n141_O_11_0_0_t1b),
    .O_12_0_0_t0b(n141_O_12_0_0_t0b),
    .O_12_0_0_t1b(n141_O_12_0_0_t1b),
    .O_13_0_0_t0b(n141_O_13_0_0_t0b),
    .O_13_0_0_t1b(n141_O_13_0_0_t1b),
    .O_14_0_0_t0b(n141_O_14_0_0_t0b),
    .O_14_0_0_t1b(n141_O_14_0_0_t1b),
    .O_15_0_0_t0b(n141_O_15_0_0_t0b),
    .O_15_0_0_t1b(n141_O_15_0_0_t1b)
  );
  FIFO_1 n142 ( // @[Top.scala 343:22]
    .clock(n142_clock),
    .reset(n142_reset),
    .valid_up(n142_valid_up),
    .valid_down(n142_valid_down),
    .I_0_0_0_t0b(n142_I_0_0_0_t0b),
    .I_0_0_0_t1b(n142_I_0_0_0_t1b),
    .I_1_0_0_t0b(n142_I_1_0_0_t0b),
    .I_1_0_0_t1b(n142_I_1_0_0_t1b),
    .I_2_0_0_t0b(n142_I_2_0_0_t0b),
    .I_2_0_0_t1b(n142_I_2_0_0_t1b),
    .I_3_0_0_t0b(n142_I_3_0_0_t0b),
    .I_3_0_0_t1b(n142_I_3_0_0_t1b),
    .I_4_0_0_t0b(n142_I_4_0_0_t0b),
    .I_4_0_0_t1b(n142_I_4_0_0_t1b),
    .I_5_0_0_t0b(n142_I_5_0_0_t0b),
    .I_5_0_0_t1b(n142_I_5_0_0_t1b),
    .I_6_0_0_t0b(n142_I_6_0_0_t0b),
    .I_6_0_0_t1b(n142_I_6_0_0_t1b),
    .I_7_0_0_t0b(n142_I_7_0_0_t0b),
    .I_7_0_0_t1b(n142_I_7_0_0_t1b),
    .I_8_0_0_t0b(n142_I_8_0_0_t0b),
    .I_8_0_0_t1b(n142_I_8_0_0_t1b),
    .I_9_0_0_t0b(n142_I_9_0_0_t0b),
    .I_9_0_0_t1b(n142_I_9_0_0_t1b),
    .I_10_0_0_t0b(n142_I_10_0_0_t0b),
    .I_10_0_0_t1b(n142_I_10_0_0_t1b),
    .I_11_0_0_t0b(n142_I_11_0_0_t0b),
    .I_11_0_0_t1b(n142_I_11_0_0_t1b),
    .I_12_0_0_t0b(n142_I_12_0_0_t0b),
    .I_12_0_0_t1b(n142_I_12_0_0_t1b),
    .I_13_0_0_t0b(n142_I_13_0_0_t0b),
    .I_13_0_0_t1b(n142_I_13_0_0_t1b),
    .I_14_0_0_t0b(n142_I_14_0_0_t0b),
    .I_14_0_0_t1b(n142_I_14_0_0_t1b),
    .I_15_0_0_t0b(n142_I_15_0_0_t0b),
    .I_15_0_0_t1b(n142_I_15_0_0_t1b),
    .O_0_0_0_t0b(n142_O_0_0_0_t0b),
    .O_0_0_0_t1b(n142_O_0_0_0_t1b),
    .O_1_0_0_t0b(n142_O_1_0_0_t0b),
    .O_1_0_0_t1b(n142_O_1_0_0_t1b),
    .O_2_0_0_t0b(n142_O_2_0_0_t0b),
    .O_2_0_0_t1b(n142_O_2_0_0_t1b),
    .O_3_0_0_t0b(n142_O_3_0_0_t0b),
    .O_3_0_0_t1b(n142_O_3_0_0_t1b),
    .O_4_0_0_t0b(n142_O_4_0_0_t0b),
    .O_4_0_0_t1b(n142_O_4_0_0_t1b),
    .O_5_0_0_t0b(n142_O_5_0_0_t0b),
    .O_5_0_0_t1b(n142_O_5_0_0_t1b),
    .O_6_0_0_t0b(n142_O_6_0_0_t0b),
    .O_6_0_0_t1b(n142_O_6_0_0_t1b),
    .O_7_0_0_t0b(n142_O_7_0_0_t0b),
    .O_7_0_0_t1b(n142_O_7_0_0_t1b),
    .O_8_0_0_t0b(n142_O_8_0_0_t0b),
    .O_8_0_0_t1b(n142_O_8_0_0_t1b),
    .O_9_0_0_t0b(n142_O_9_0_0_t0b),
    .O_9_0_0_t1b(n142_O_9_0_0_t1b),
    .O_10_0_0_t0b(n142_O_10_0_0_t0b),
    .O_10_0_0_t1b(n142_O_10_0_0_t1b),
    .O_11_0_0_t0b(n142_O_11_0_0_t0b),
    .O_11_0_0_t1b(n142_O_11_0_0_t1b),
    .O_12_0_0_t0b(n142_O_12_0_0_t0b),
    .O_12_0_0_t1b(n142_O_12_0_0_t1b),
    .O_13_0_0_t0b(n142_O_13_0_0_t0b),
    .O_13_0_0_t1b(n142_O_13_0_0_t1b),
    .O_14_0_0_t0b(n142_O_14_0_0_t0b),
    .O_14_0_0_t1b(n142_O_14_0_0_t1b),
    .O_15_0_0_t0b(n142_O_15_0_0_t0b),
    .O_15_0_0_t1b(n142_O_15_0_0_t1b)
  );
  Map2T_9 n143 ( // @[Top.scala 346:22]
    .clock(n143_clock),
    .reset(n143_reset),
    .valid_up(n143_valid_up),
    .valid_down(n143_valid_down),
    .I0_0_0_0(n143_I0_0_0_0),
    .I0_0_0_1(n143_I0_0_0_1),
    .I0_0_0_2(n143_I0_0_0_2),
    .I0_0_1_0(n143_I0_0_1_0),
    .I0_0_1_1(n143_I0_0_1_1),
    .I0_0_1_2(n143_I0_0_1_2),
    .I0_0_2_0(n143_I0_0_2_0),
    .I0_0_2_1(n143_I0_0_2_1),
    .I0_0_2_2(n143_I0_0_2_2),
    .I0_1_0_0(n143_I0_1_0_0),
    .I0_1_0_1(n143_I0_1_0_1),
    .I0_1_0_2(n143_I0_1_0_2),
    .I0_1_1_0(n143_I0_1_1_0),
    .I0_1_1_1(n143_I0_1_1_1),
    .I0_1_1_2(n143_I0_1_1_2),
    .I0_1_2_0(n143_I0_1_2_0),
    .I0_1_2_1(n143_I0_1_2_1),
    .I0_1_2_2(n143_I0_1_2_2),
    .I0_2_0_0(n143_I0_2_0_0),
    .I0_2_0_1(n143_I0_2_0_1),
    .I0_2_0_2(n143_I0_2_0_2),
    .I0_2_1_0(n143_I0_2_1_0),
    .I0_2_1_1(n143_I0_2_1_1),
    .I0_2_1_2(n143_I0_2_1_2),
    .I0_2_2_0(n143_I0_2_2_0),
    .I0_2_2_1(n143_I0_2_2_1),
    .I0_2_2_2(n143_I0_2_2_2),
    .I0_3_0_0(n143_I0_3_0_0),
    .I0_3_0_1(n143_I0_3_0_1),
    .I0_3_0_2(n143_I0_3_0_2),
    .I0_3_1_0(n143_I0_3_1_0),
    .I0_3_1_1(n143_I0_3_1_1),
    .I0_3_1_2(n143_I0_3_1_2),
    .I0_3_2_0(n143_I0_3_2_0),
    .I0_3_2_1(n143_I0_3_2_1),
    .I0_3_2_2(n143_I0_3_2_2),
    .I0_4_0_0(n143_I0_4_0_0),
    .I0_4_0_1(n143_I0_4_0_1),
    .I0_4_0_2(n143_I0_4_0_2),
    .I0_4_1_0(n143_I0_4_1_0),
    .I0_4_1_1(n143_I0_4_1_1),
    .I0_4_1_2(n143_I0_4_1_2),
    .I0_4_2_0(n143_I0_4_2_0),
    .I0_4_2_1(n143_I0_4_2_1),
    .I0_4_2_2(n143_I0_4_2_2),
    .I0_5_0_0(n143_I0_5_0_0),
    .I0_5_0_1(n143_I0_5_0_1),
    .I0_5_0_2(n143_I0_5_0_2),
    .I0_5_1_0(n143_I0_5_1_0),
    .I0_5_1_1(n143_I0_5_1_1),
    .I0_5_1_2(n143_I0_5_1_2),
    .I0_5_2_0(n143_I0_5_2_0),
    .I0_5_2_1(n143_I0_5_2_1),
    .I0_5_2_2(n143_I0_5_2_2),
    .I0_6_0_0(n143_I0_6_0_0),
    .I0_6_0_1(n143_I0_6_0_1),
    .I0_6_0_2(n143_I0_6_0_2),
    .I0_6_1_0(n143_I0_6_1_0),
    .I0_6_1_1(n143_I0_6_1_1),
    .I0_6_1_2(n143_I0_6_1_2),
    .I0_6_2_0(n143_I0_6_2_0),
    .I0_6_2_1(n143_I0_6_2_1),
    .I0_6_2_2(n143_I0_6_2_2),
    .I0_7_0_0(n143_I0_7_0_0),
    .I0_7_0_1(n143_I0_7_0_1),
    .I0_7_0_2(n143_I0_7_0_2),
    .I0_7_1_0(n143_I0_7_1_0),
    .I0_7_1_1(n143_I0_7_1_1),
    .I0_7_1_2(n143_I0_7_1_2),
    .I0_7_2_0(n143_I0_7_2_0),
    .I0_7_2_1(n143_I0_7_2_1),
    .I0_7_2_2(n143_I0_7_2_2),
    .I0_8_0_0(n143_I0_8_0_0),
    .I0_8_0_1(n143_I0_8_0_1),
    .I0_8_0_2(n143_I0_8_0_2),
    .I0_8_1_0(n143_I0_8_1_0),
    .I0_8_1_1(n143_I0_8_1_1),
    .I0_8_1_2(n143_I0_8_1_2),
    .I0_8_2_0(n143_I0_8_2_0),
    .I0_8_2_1(n143_I0_8_2_1),
    .I0_8_2_2(n143_I0_8_2_2),
    .I0_9_0_0(n143_I0_9_0_0),
    .I0_9_0_1(n143_I0_9_0_1),
    .I0_9_0_2(n143_I0_9_0_2),
    .I0_9_1_0(n143_I0_9_1_0),
    .I0_9_1_1(n143_I0_9_1_1),
    .I0_9_1_2(n143_I0_9_1_2),
    .I0_9_2_0(n143_I0_9_2_0),
    .I0_9_2_1(n143_I0_9_2_1),
    .I0_9_2_2(n143_I0_9_2_2),
    .I0_10_0_0(n143_I0_10_0_0),
    .I0_10_0_1(n143_I0_10_0_1),
    .I0_10_0_2(n143_I0_10_0_2),
    .I0_10_1_0(n143_I0_10_1_0),
    .I0_10_1_1(n143_I0_10_1_1),
    .I0_10_1_2(n143_I0_10_1_2),
    .I0_10_2_0(n143_I0_10_2_0),
    .I0_10_2_1(n143_I0_10_2_1),
    .I0_10_2_2(n143_I0_10_2_2),
    .I0_11_0_0(n143_I0_11_0_0),
    .I0_11_0_1(n143_I0_11_0_1),
    .I0_11_0_2(n143_I0_11_0_2),
    .I0_11_1_0(n143_I0_11_1_0),
    .I0_11_1_1(n143_I0_11_1_1),
    .I0_11_1_2(n143_I0_11_1_2),
    .I0_11_2_0(n143_I0_11_2_0),
    .I0_11_2_1(n143_I0_11_2_1),
    .I0_11_2_2(n143_I0_11_2_2),
    .I0_12_0_0(n143_I0_12_0_0),
    .I0_12_0_1(n143_I0_12_0_1),
    .I0_12_0_2(n143_I0_12_0_2),
    .I0_12_1_0(n143_I0_12_1_0),
    .I0_12_1_1(n143_I0_12_1_1),
    .I0_12_1_2(n143_I0_12_1_2),
    .I0_12_2_0(n143_I0_12_2_0),
    .I0_12_2_1(n143_I0_12_2_1),
    .I0_12_2_2(n143_I0_12_2_2),
    .I0_13_0_0(n143_I0_13_0_0),
    .I0_13_0_1(n143_I0_13_0_1),
    .I0_13_0_2(n143_I0_13_0_2),
    .I0_13_1_0(n143_I0_13_1_0),
    .I0_13_1_1(n143_I0_13_1_1),
    .I0_13_1_2(n143_I0_13_1_2),
    .I0_13_2_0(n143_I0_13_2_0),
    .I0_13_2_1(n143_I0_13_2_1),
    .I0_13_2_2(n143_I0_13_2_2),
    .I0_14_0_0(n143_I0_14_0_0),
    .I0_14_0_1(n143_I0_14_0_1),
    .I0_14_0_2(n143_I0_14_0_2),
    .I0_14_1_0(n143_I0_14_1_0),
    .I0_14_1_1(n143_I0_14_1_1),
    .I0_14_1_2(n143_I0_14_1_2),
    .I0_14_2_0(n143_I0_14_2_0),
    .I0_14_2_1(n143_I0_14_2_1),
    .I0_14_2_2(n143_I0_14_2_2),
    .I0_15_0_0(n143_I0_15_0_0),
    .I0_15_0_1(n143_I0_15_0_1),
    .I0_15_0_2(n143_I0_15_0_2),
    .I0_15_1_0(n143_I0_15_1_0),
    .I0_15_1_1(n143_I0_15_1_1),
    .I0_15_1_2(n143_I0_15_1_2),
    .I0_15_2_0(n143_I0_15_2_0),
    .I0_15_2_1(n143_I0_15_2_1),
    .I0_15_2_2(n143_I0_15_2_2),
    .I1_0_0_0_t0b(n143_I1_0_0_0_t0b),
    .I1_0_0_0_t1b(n143_I1_0_0_0_t1b),
    .I1_1_0_0_t0b(n143_I1_1_0_0_t0b),
    .I1_1_0_0_t1b(n143_I1_1_0_0_t1b),
    .I1_2_0_0_t0b(n143_I1_2_0_0_t0b),
    .I1_2_0_0_t1b(n143_I1_2_0_0_t1b),
    .I1_3_0_0_t0b(n143_I1_3_0_0_t0b),
    .I1_3_0_0_t1b(n143_I1_3_0_0_t1b),
    .I1_4_0_0_t0b(n143_I1_4_0_0_t0b),
    .I1_4_0_0_t1b(n143_I1_4_0_0_t1b),
    .I1_5_0_0_t0b(n143_I1_5_0_0_t0b),
    .I1_5_0_0_t1b(n143_I1_5_0_0_t1b),
    .I1_6_0_0_t0b(n143_I1_6_0_0_t0b),
    .I1_6_0_0_t1b(n143_I1_6_0_0_t1b),
    .I1_7_0_0_t0b(n143_I1_7_0_0_t0b),
    .I1_7_0_0_t1b(n143_I1_7_0_0_t1b),
    .I1_8_0_0_t0b(n143_I1_8_0_0_t0b),
    .I1_8_0_0_t1b(n143_I1_8_0_0_t1b),
    .I1_9_0_0_t0b(n143_I1_9_0_0_t0b),
    .I1_9_0_0_t1b(n143_I1_9_0_0_t1b),
    .I1_10_0_0_t0b(n143_I1_10_0_0_t0b),
    .I1_10_0_0_t1b(n143_I1_10_0_0_t1b),
    .I1_11_0_0_t0b(n143_I1_11_0_0_t0b),
    .I1_11_0_0_t1b(n143_I1_11_0_0_t1b),
    .I1_12_0_0_t0b(n143_I1_12_0_0_t0b),
    .I1_12_0_0_t1b(n143_I1_12_0_0_t1b),
    .I1_13_0_0_t0b(n143_I1_13_0_0_t0b),
    .I1_13_0_0_t1b(n143_I1_13_0_0_t1b),
    .I1_14_0_0_t0b(n143_I1_14_0_0_t0b),
    .I1_14_0_0_t1b(n143_I1_14_0_0_t1b),
    .I1_15_0_0_t0b(n143_I1_15_0_0_t0b),
    .I1_15_0_0_t1b(n143_I1_15_0_0_t1b),
    .O_0_0_0_t0b(n143_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(n143_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(n143_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(n143_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(n143_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(n143_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(n143_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(n143_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(n143_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(n143_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(n143_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(n143_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(n143_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(n143_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(n143_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(n143_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(n143_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(n143_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(n143_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(n143_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(n143_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(n143_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(n143_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(n143_O_7_0_0_t1b_t1b),
    .O_8_0_0_t0b(n143_O_8_0_0_t0b),
    .O_8_0_0_t1b_t0b(n143_O_8_0_0_t1b_t0b),
    .O_8_0_0_t1b_t1b(n143_O_8_0_0_t1b_t1b),
    .O_9_0_0_t0b(n143_O_9_0_0_t0b),
    .O_9_0_0_t1b_t0b(n143_O_9_0_0_t1b_t0b),
    .O_9_0_0_t1b_t1b(n143_O_9_0_0_t1b_t1b),
    .O_10_0_0_t0b(n143_O_10_0_0_t0b),
    .O_10_0_0_t1b_t0b(n143_O_10_0_0_t1b_t0b),
    .O_10_0_0_t1b_t1b(n143_O_10_0_0_t1b_t1b),
    .O_11_0_0_t0b(n143_O_11_0_0_t0b),
    .O_11_0_0_t1b_t0b(n143_O_11_0_0_t1b_t0b),
    .O_11_0_0_t1b_t1b(n143_O_11_0_0_t1b_t1b),
    .O_12_0_0_t0b(n143_O_12_0_0_t0b),
    .O_12_0_0_t1b_t0b(n143_O_12_0_0_t1b_t0b),
    .O_12_0_0_t1b_t1b(n143_O_12_0_0_t1b_t1b),
    .O_13_0_0_t0b(n143_O_13_0_0_t0b),
    .O_13_0_0_t1b_t0b(n143_O_13_0_0_t1b_t0b),
    .O_13_0_0_t1b_t1b(n143_O_13_0_0_t1b_t1b),
    .O_14_0_0_t0b(n143_O_14_0_0_t0b),
    .O_14_0_0_t1b_t0b(n143_O_14_0_0_t1b_t0b),
    .O_14_0_0_t1b_t1b(n143_O_14_0_0_t1b_t1b),
    .O_15_0_0_t0b(n143_O_15_0_0_t0b),
    .O_15_0_0_t1b_t0b(n143_O_15_0_0_t1b_t0b),
    .O_15_0_0_t1b_t1b(n143_O_15_0_0_t1b_t1b)
  );
  assign valid_down = n143_valid_down; // @[Top.scala 351:16]
  assign O_0_0_0_t0b = n143_O_0_0_0_t0b; // @[Top.scala 350:7]
  assign O_0_0_0_t1b_t0b = n143_O_0_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_0_0_0_t1b_t1b = n143_O_0_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_1_0_0_t0b = n143_O_1_0_0_t0b; // @[Top.scala 350:7]
  assign O_1_0_0_t1b_t0b = n143_O_1_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_1_0_0_t1b_t1b = n143_O_1_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_2_0_0_t0b = n143_O_2_0_0_t0b; // @[Top.scala 350:7]
  assign O_2_0_0_t1b_t0b = n143_O_2_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_2_0_0_t1b_t1b = n143_O_2_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_3_0_0_t0b = n143_O_3_0_0_t0b; // @[Top.scala 350:7]
  assign O_3_0_0_t1b_t0b = n143_O_3_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_3_0_0_t1b_t1b = n143_O_3_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_4_0_0_t0b = n143_O_4_0_0_t0b; // @[Top.scala 350:7]
  assign O_4_0_0_t1b_t0b = n143_O_4_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_4_0_0_t1b_t1b = n143_O_4_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_5_0_0_t0b = n143_O_5_0_0_t0b; // @[Top.scala 350:7]
  assign O_5_0_0_t1b_t0b = n143_O_5_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_5_0_0_t1b_t1b = n143_O_5_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_6_0_0_t0b = n143_O_6_0_0_t0b; // @[Top.scala 350:7]
  assign O_6_0_0_t1b_t0b = n143_O_6_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_6_0_0_t1b_t1b = n143_O_6_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_7_0_0_t0b = n143_O_7_0_0_t0b; // @[Top.scala 350:7]
  assign O_7_0_0_t1b_t0b = n143_O_7_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_7_0_0_t1b_t1b = n143_O_7_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_8_0_0_t0b = n143_O_8_0_0_t0b; // @[Top.scala 350:7]
  assign O_8_0_0_t1b_t0b = n143_O_8_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_8_0_0_t1b_t1b = n143_O_8_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_9_0_0_t0b = n143_O_9_0_0_t0b; // @[Top.scala 350:7]
  assign O_9_0_0_t1b_t0b = n143_O_9_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_9_0_0_t1b_t1b = n143_O_9_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_10_0_0_t0b = n143_O_10_0_0_t0b; // @[Top.scala 350:7]
  assign O_10_0_0_t1b_t0b = n143_O_10_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_10_0_0_t1b_t1b = n143_O_10_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_11_0_0_t0b = n143_O_11_0_0_t0b; // @[Top.scala 350:7]
  assign O_11_0_0_t1b_t0b = n143_O_11_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_11_0_0_t1b_t1b = n143_O_11_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_12_0_0_t0b = n143_O_12_0_0_t0b; // @[Top.scala 350:7]
  assign O_12_0_0_t1b_t0b = n143_O_12_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_12_0_0_t1b_t1b = n143_O_12_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_13_0_0_t0b = n143_O_13_0_0_t0b; // @[Top.scala 350:7]
  assign O_13_0_0_t1b_t0b = n143_O_13_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_13_0_0_t1b_t1b = n143_O_13_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_14_0_0_t0b = n143_O_14_0_0_t0b; // @[Top.scala 350:7]
  assign O_14_0_0_t1b_t0b = n143_O_14_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_14_0_0_t1b_t1b = n143_O_14_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign O_15_0_0_t0b = n143_O_15_0_0_t0b; // @[Top.scala 350:7]
  assign O_15_0_0_t1b_t0b = n143_O_15_0_0_t1b_t0b; // @[Top.scala 350:7]
  assign O_15_0_0_t1b_t1b = n143_O_15_0_0_t1b_t1b; // @[Top.scala 350:7]
  assign counter108_clock = clock;
  assign counter108_reset = reset;
  assign n116_I_0 = counter108_O_0; // @[Top.scala 328:12]
  assign n116_I_1 = counter108_O_1; // @[Top.scala 328:12]
  assign n116_I_2 = counter108_O_2; // @[Top.scala 328:12]
  assign n116_I_3 = counter108_O_3; // @[Top.scala 328:12]
  assign n116_I_4 = counter108_O_4; // @[Top.scala 328:12]
  assign n116_I_5 = counter108_O_5; // @[Top.scala 328:12]
  assign n116_I_6 = counter108_O_6; // @[Top.scala 328:12]
  assign n116_I_7 = counter108_O_7; // @[Top.scala 328:12]
  assign n116_I_8 = counter108_O_8; // @[Top.scala 328:12]
  assign n116_I_9 = counter108_O_9; // @[Top.scala 328:12]
  assign n116_I_10 = counter108_O_10; // @[Top.scala 328:12]
  assign n116_I_11 = counter108_O_11; // @[Top.scala 328:12]
  assign n116_I_12 = counter108_O_12; // @[Top.scala 328:12]
  assign n116_I_13 = counter108_O_13; // @[Top.scala 328:12]
  assign n116_I_14 = counter108_O_14; // @[Top.scala 328:12]
  assign n116_I_15 = counter108_O_15; // @[Top.scala 328:12]
  assign n128_I_0 = counter108_O_0; // @[Top.scala 331:12]
  assign n128_I_1 = counter108_O_1; // @[Top.scala 331:12]
  assign n128_I_2 = counter108_O_2; // @[Top.scala 331:12]
  assign n128_I_3 = counter108_O_3; // @[Top.scala 331:12]
  assign n128_I_4 = counter108_O_4; // @[Top.scala 331:12]
  assign n128_I_5 = counter108_O_5; // @[Top.scala 331:12]
  assign n128_I_6 = counter108_O_6; // @[Top.scala 331:12]
  assign n128_I_7 = counter108_O_7; // @[Top.scala 331:12]
  assign n128_I_8 = counter108_O_8; // @[Top.scala 331:12]
  assign n128_I_9 = counter108_O_9; // @[Top.scala 331:12]
  assign n128_I_10 = counter108_O_10; // @[Top.scala 331:12]
  assign n128_I_11 = counter108_O_11; // @[Top.scala 331:12]
  assign n128_I_12 = counter108_O_12; // @[Top.scala 331:12]
  assign n128_I_13 = counter108_O_13; // @[Top.scala 331:12]
  assign n128_I_14 = counter108_O_14; // @[Top.scala 331:12]
  assign n128_I_15 = counter108_O_15; // @[Top.scala 331:12]
  assign n129_valid_up = n116_valid_down & n128_valid_down; // @[Top.scala 336:19]
  assign n129_I0_0 = n116_O_0; // @[Top.scala 334:13]
  assign n129_I0_1 = n116_O_1; // @[Top.scala 334:13]
  assign n129_I0_2 = n116_O_2; // @[Top.scala 334:13]
  assign n129_I0_3 = n116_O_3; // @[Top.scala 334:13]
  assign n129_I0_4 = n116_O_4; // @[Top.scala 334:13]
  assign n129_I0_5 = n116_O_5; // @[Top.scala 334:13]
  assign n129_I0_6 = n116_O_6; // @[Top.scala 334:13]
  assign n129_I0_7 = n116_O_7; // @[Top.scala 334:13]
  assign n129_I0_8 = n116_O_8; // @[Top.scala 334:13]
  assign n129_I0_9 = n116_O_9; // @[Top.scala 334:13]
  assign n129_I0_10 = n116_O_10; // @[Top.scala 334:13]
  assign n129_I0_11 = n116_O_11; // @[Top.scala 334:13]
  assign n129_I0_12 = n116_O_12; // @[Top.scala 334:13]
  assign n129_I0_13 = n116_O_13; // @[Top.scala 334:13]
  assign n129_I0_14 = n116_O_14; // @[Top.scala 334:13]
  assign n129_I0_15 = n116_O_15; // @[Top.scala 334:13]
  assign n129_I1_0 = n128_O_0; // @[Top.scala 335:13]
  assign n129_I1_1 = n128_O_1; // @[Top.scala 335:13]
  assign n129_I1_2 = n128_O_2; // @[Top.scala 335:13]
  assign n129_I1_3 = n128_O_3; // @[Top.scala 335:13]
  assign n129_I1_4 = n128_O_4; // @[Top.scala 335:13]
  assign n129_I1_5 = n128_O_5; // @[Top.scala 335:13]
  assign n129_I1_6 = n128_O_6; // @[Top.scala 335:13]
  assign n129_I1_7 = n128_O_7; // @[Top.scala 335:13]
  assign n129_I1_8 = n128_O_8; // @[Top.scala 335:13]
  assign n129_I1_9 = n128_O_9; // @[Top.scala 335:13]
  assign n129_I1_10 = n128_O_10; // @[Top.scala 335:13]
  assign n129_I1_11 = n128_O_11; // @[Top.scala 335:13]
  assign n129_I1_12 = n128_O_12; // @[Top.scala 335:13]
  assign n129_I1_13 = n128_O_13; // @[Top.scala 335:13]
  assign n129_I1_14 = n128_O_14; // @[Top.scala 335:13]
  assign n129_I1_15 = n128_O_15; // @[Top.scala 335:13]
  assign n138_valid_up = n129_valid_down; // @[Top.scala 339:19]
  assign n138_I_0_t0b = n129_O_0_t0b; // @[Top.scala 338:12]
  assign n138_I_0_t1b = n129_O_0_t1b; // @[Top.scala 338:12]
  assign n138_I_1_t0b = n129_O_1_t0b; // @[Top.scala 338:12]
  assign n138_I_1_t1b = n129_O_1_t1b; // @[Top.scala 338:12]
  assign n138_I_2_t0b = n129_O_2_t0b; // @[Top.scala 338:12]
  assign n138_I_2_t1b = n129_O_2_t1b; // @[Top.scala 338:12]
  assign n138_I_3_t0b = n129_O_3_t0b; // @[Top.scala 338:12]
  assign n138_I_3_t1b = n129_O_3_t1b; // @[Top.scala 338:12]
  assign n138_I_4_t0b = n129_O_4_t0b; // @[Top.scala 338:12]
  assign n138_I_4_t1b = n129_O_4_t1b; // @[Top.scala 338:12]
  assign n138_I_5_t0b = n129_O_5_t0b; // @[Top.scala 338:12]
  assign n138_I_5_t1b = n129_O_5_t1b; // @[Top.scala 338:12]
  assign n138_I_6_t0b = n129_O_6_t0b; // @[Top.scala 338:12]
  assign n138_I_6_t1b = n129_O_6_t1b; // @[Top.scala 338:12]
  assign n138_I_7_t0b = n129_O_7_t0b; // @[Top.scala 338:12]
  assign n138_I_7_t1b = n129_O_7_t1b; // @[Top.scala 338:12]
  assign n138_I_8_t0b = n129_O_8_t0b; // @[Top.scala 338:12]
  assign n138_I_8_t1b = n129_O_8_t1b; // @[Top.scala 338:12]
  assign n138_I_9_t0b = n129_O_9_t0b; // @[Top.scala 338:12]
  assign n138_I_9_t1b = n129_O_9_t1b; // @[Top.scala 338:12]
  assign n138_I_10_t0b = n129_O_10_t0b; // @[Top.scala 338:12]
  assign n138_I_10_t1b = n129_O_10_t1b; // @[Top.scala 338:12]
  assign n138_I_11_t0b = n129_O_11_t0b; // @[Top.scala 338:12]
  assign n138_I_11_t1b = n129_O_11_t1b; // @[Top.scala 338:12]
  assign n138_I_12_t0b = n129_O_12_t0b; // @[Top.scala 338:12]
  assign n138_I_12_t1b = n129_O_12_t1b; // @[Top.scala 338:12]
  assign n138_I_13_t0b = n129_O_13_t0b; // @[Top.scala 338:12]
  assign n138_I_13_t1b = n129_O_13_t1b; // @[Top.scala 338:12]
  assign n138_I_14_t0b = n129_O_14_t0b; // @[Top.scala 338:12]
  assign n138_I_14_t1b = n129_O_14_t1b; // @[Top.scala 338:12]
  assign n138_I_15_t0b = n129_O_15_t0b; // @[Top.scala 338:12]
  assign n138_I_15_t1b = n129_O_15_t1b; // @[Top.scala 338:12]
  assign n141_valid_up = n138_valid_down; // @[Top.scala 342:19]
  assign n141_I_0_0_t0b = n138_O_0_0_t0b; // @[Top.scala 341:12]
  assign n141_I_0_0_t1b = n138_O_0_0_t1b; // @[Top.scala 341:12]
  assign n141_I_1_0_t0b = n138_O_1_0_t0b; // @[Top.scala 341:12]
  assign n141_I_1_0_t1b = n138_O_1_0_t1b; // @[Top.scala 341:12]
  assign n141_I_2_0_t0b = n138_O_2_0_t0b; // @[Top.scala 341:12]
  assign n141_I_2_0_t1b = n138_O_2_0_t1b; // @[Top.scala 341:12]
  assign n141_I_3_0_t0b = n138_O_3_0_t0b; // @[Top.scala 341:12]
  assign n141_I_3_0_t1b = n138_O_3_0_t1b; // @[Top.scala 341:12]
  assign n141_I_4_0_t0b = n138_O_4_0_t0b; // @[Top.scala 341:12]
  assign n141_I_4_0_t1b = n138_O_4_0_t1b; // @[Top.scala 341:12]
  assign n141_I_5_0_t0b = n138_O_5_0_t0b; // @[Top.scala 341:12]
  assign n141_I_5_0_t1b = n138_O_5_0_t1b; // @[Top.scala 341:12]
  assign n141_I_6_0_t0b = n138_O_6_0_t0b; // @[Top.scala 341:12]
  assign n141_I_6_0_t1b = n138_O_6_0_t1b; // @[Top.scala 341:12]
  assign n141_I_7_0_t0b = n138_O_7_0_t0b; // @[Top.scala 341:12]
  assign n141_I_7_0_t1b = n138_O_7_0_t1b; // @[Top.scala 341:12]
  assign n141_I_8_0_t0b = n138_O_8_0_t0b; // @[Top.scala 341:12]
  assign n141_I_8_0_t1b = n138_O_8_0_t1b; // @[Top.scala 341:12]
  assign n141_I_9_0_t0b = n138_O_9_0_t0b; // @[Top.scala 341:12]
  assign n141_I_9_0_t1b = n138_O_9_0_t1b; // @[Top.scala 341:12]
  assign n141_I_10_0_t0b = n138_O_10_0_t0b; // @[Top.scala 341:12]
  assign n141_I_10_0_t1b = n138_O_10_0_t1b; // @[Top.scala 341:12]
  assign n141_I_11_0_t0b = n138_O_11_0_t0b; // @[Top.scala 341:12]
  assign n141_I_11_0_t1b = n138_O_11_0_t1b; // @[Top.scala 341:12]
  assign n141_I_12_0_t0b = n138_O_12_0_t0b; // @[Top.scala 341:12]
  assign n141_I_12_0_t1b = n138_O_12_0_t1b; // @[Top.scala 341:12]
  assign n141_I_13_0_t0b = n138_O_13_0_t0b; // @[Top.scala 341:12]
  assign n141_I_13_0_t1b = n138_O_13_0_t1b; // @[Top.scala 341:12]
  assign n141_I_14_0_t0b = n138_O_14_0_t0b; // @[Top.scala 341:12]
  assign n141_I_14_0_t1b = n138_O_14_0_t1b; // @[Top.scala 341:12]
  assign n141_I_15_0_t0b = n138_O_15_0_t0b; // @[Top.scala 341:12]
  assign n141_I_15_0_t1b = n138_O_15_0_t1b; // @[Top.scala 341:12]
  assign n142_clock = clock;
  assign n142_reset = reset;
  assign n142_valid_up = n141_valid_down; // @[Top.scala 345:19]
  assign n142_I_0_0_0_t0b = n141_O_0_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_0_0_0_t1b = n141_O_0_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_1_0_0_t0b = n141_O_1_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_1_0_0_t1b = n141_O_1_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_2_0_0_t0b = n141_O_2_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_2_0_0_t1b = n141_O_2_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_3_0_0_t0b = n141_O_3_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_3_0_0_t1b = n141_O_3_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_4_0_0_t0b = n141_O_4_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_4_0_0_t1b = n141_O_4_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_5_0_0_t0b = n141_O_5_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_5_0_0_t1b = n141_O_5_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_6_0_0_t0b = n141_O_6_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_6_0_0_t1b = n141_O_6_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_7_0_0_t0b = n141_O_7_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_7_0_0_t1b = n141_O_7_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_8_0_0_t0b = n141_O_8_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_8_0_0_t1b = n141_O_8_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_9_0_0_t0b = n141_O_9_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_9_0_0_t1b = n141_O_9_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_10_0_0_t0b = n141_O_10_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_10_0_0_t1b = n141_O_10_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_11_0_0_t0b = n141_O_11_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_11_0_0_t1b = n141_O_11_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_12_0_0_t0b = n141_O_12_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_12_0_0_t1b = n141_O_12_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_13_0_0_t0b = n141_O_13_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_13_0_0_t1b = n141_O_13_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_14_0_0_t0b = n141_O_14_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_14_0_0_t1b = n141_O_14_0_0_t1b; // @[Top.scala 344:12]
  assign n142_I_15_0_0_t0b = n141_O_15_0_0_t0b; // @[Top.scala 344:12]
  assign n142_I_15_0_0_t1b = n141_O_15_0_0_t1b; // @[Top.scala 344:12]
  assign n143_clock = clock;
  assign n143_reset = reset;
  assign n143_valid_up = valid_up & n142_valid_down; // @[Top.scala 349:19]
  assign n143_I0_0_0_0 = I_0_0_0; // @[Top.scala 347:13]
  assign n143_I0_0_0_1 = I_0_0_1; // @[Top.scala 347:13]
  assign n143_I0_0_0_2 = I_0_0_2; // @[Top.scala 347:13]
  assign n143_I0_0_1_0 = I_0_1_0; // @[Top.scala 347:13]
  assign n143_I0_0_1_1 = I_0_1_1; // @[Top.scala 347:13]
  assign n143_I0_0_1_2 = I_0_1_2; // @[Top.scala 347:13]
  assign n143_I0_0_2_0 = I_0_2_0; // @[Top.scala 347:13]
  assign n143_I0_0_2_1 = I_0_2_1; // @[Top.scala 347:13]
  assign n143_I0_0_2_2 = I_0_2_2; // @[Top.scala 347:13]
  assign n143_I0_1_0_0 = I_1_0_0; // @[Top.scala 347:13]
  assign n143_I0_1_0_1 = I_1_0_1; // @[Top.scala 347:13]
  assign n143_I0_1_0_2 = I_1_0_2; // @[Top.scala 347:13]
  assign n143_I0_1_1_0 = I_1_1_0; // @[Top.scala 347:13]
  assign n143_I0_1_1_1 = I_1_1_1; // @[Top.scala 347:13]
  assign n143_I0_1_1_2 = I_1_1_2; // @[Top.scala 347:13]
  assign n143_I0_1_2_0 = I_1_2_0; // @[Top.scala 347:13]
  assign n143_I0_1_2_1 = I_1_2_1; // @[Top.scala 347:13]
  assign n143_I0_1_2_2 = I_1_2_2; // @[Top.scala 347:13]
  assign n143_I0_2_0_0 = I_2_0_0; // @[Top.scala 347:13]
  assign n143_I0_2_0_1 = I_2_0_1; // @[Top.scala 347:13]
  assign n143_I0_2_0_2 = I_2_0_2; // @[Top.scala 347:13]
  assign n143_I0_2_1_0 = I_2_1_0; // @[Top.scala 347:13]
  assign n143_I0_2_1_1 = I_2_1_1; // @[Top.scala 347:13]
  assign n143_I0_2_1_2 = I_2_1_2; // @[Top.scala 347:13]
  assign n143_I0_2_2_0 = I_2_2_0; // @[Top.scala 347:13]
  assign n143_I0_2_2_1 = I_2_2_1; // @[Top.scala 347:13]
  assign n143_I0_2_2_2 = I_2_2_2; // @[Top.scala 347:13]
  assign n143_I0_3_0_0 = I_3_0_0; // @[Top.scala 347:13]
  assign n143_I0_3_0_1 = I_3_0_1; // @[Top.scala 347:13]
  assign n143_I0_3_0_2 = I_3_0_2; // @[Top.scala 347:13]
  assign n143_I0_3_1_0 = I_3_1_0; // @[Top.scala 347:13]
  assign n143_I0_3_1_1 = I_3_1_1; // @[Top.scala 347:13]
  assign n143_I0_3_1_2 = I_3_1_2; // @[Top.scala 347:13]
  assign n143_I0_3_2_0 = I_3_2_0; // @[Top.scala 347:13]
  assign n143_I0_3_2_1 = I_3_2_1; // @[Top.scala 347:13]
  assign n143_I0_3_2_2 = I_3_2_2; // @[Top.scala 347:13]
  assign n143_I0_4_0_0 = I_4_0_0; // @[Top.scala 347:13]
  assign n143_I0_4_0_1 = I_4_0_1; // @[Top.scala 347:13]
  assign n143_I0_4_0_2 = I_4_0_2; // @[Top.scala 347:13]
  assign n143_I0_4_1_0 = I_4_1_0; // @[Top.scala 347:13]
  assign n143_I0_4_1_1 = I_4_1_1; // @[Top.scala 347:13]
  assign n143_I0_4_1_2 = I_4_1_2; // @[Top.scala 347:13]
  assign n143_I0_4_2_0 = I_4_2_0; // @[Top.scala 347:13]
  assign n143_I0_4_2_1 = I_4_2_1; // @[Top.scala 347:13]
  assign n143_I0_4_2_2 = I_4_2_2; // @[Top.scala 347:13]
  assign n143_I0_5_0_0 = I_5_0_0; // @[Top.scala 347:13]
  assign n143_I0_5_0_1 = I_5_0_1; // @[Top.scala 347:13]
  assign n143_I0_5_0_2 = I_5_0_2; // @[Top.scala 347:13]
  assign n143_I0_5_1_0 = I_5_1_0; // @[Top.scala 347:13]
  assign n143_I0_5_1_1 = I_5_1_1; // @[Top.scala 347:13]
  assign n143_I0_5_1_2 = I_5_1_2; // @[Top.scala 347:13]
  assign n143_I0_5_2_0 = I_5_2_0; // @[Top.scala 347:13]
  assign n143_I0_5_2_1 = I_5_2_1; // @[Top.scala 347:13]
  assign n143_I0_5_2_2 = I_5_2_2; // @[Top.scala 347:13]
  assign n143_I0_6_0_0 = I_6_0_0; // @[Top.scala 347:13]
  assign n143_I0_6_0_1 = I_6_0_1; // @[Top.scala 347:13]
  assign n143_I0_6_0_2 = I_6_0_2; // @[Top.scala 347:13]
  assign n143_I0_6_1_0 = I_6_1_0; // @[Top.scala 347:13]
  assign n143_I0_6_1_1 = I_6_1_1; // @[Top.scala 347:13]
  assign n143_I0_6_1_2 = I_6_1_2; // @[Top.scala 347:13]
  assign n143_I0_6_2_0 = I_6_2_0; // @[Top.scala 347:13]
  assign n143_I0_6_2_1 = I_6_2_1; // @[Top.scala 347:13]
  assign n143_I0_6_2_2 = I_6_2_2; // @[Top.scala 347:13]
  assign n143_I0_7_0_0 = I_7_0_0; // @[Top.scala 347:13]
  assign n143_I0_7_0_1 = I_7_0_1; // @[Top.scala 347:13]
  assign n143_I0_7_0_2 = I_7_0_2; // @[Top.scala 347:13]
  assign n143_I0_7_1_0 = I_7_1_0; // @[Top.scala 347:13]
  assign n143_I0_7_1_1 = I_7_1_1; // @[Top.scala 347:13]
  assign n143_I0_7_1_2 = I_7_1_2; // @[Top.scala 347:13]
  assign n143_I0_7_2_0 = I_7_2_0; // @[Top.scala 347:13]
  assign n143_I0_7_2_1 = I_7_2_1; // @[Top.scala 347:13]
  assign n143_I0_7_2_2 = I_7_2_2; // @[Top.scala 347:13]
  assign n143_I0_8_0_0 = I_8_0_0; // @[Top.scala 347:13]
  assign n143_I0_8_0_1 = I_8_0_1; // @[Top.scala 347:13]
  assign n143_I0_8_0_2 = I_8_0_2; // @[Top.scala 347:13]
  assign n143_I0_8_1_0 = I_8_1_0; // @[Top.scala 347:13]
  assign n143_I0_8_1_1 = I_8_1_1; // @[Top.scala 347:13]
  assign n143_I0_8_1_2 = I_8_1_2; // @[Top.scala 347:13]
  assign n143_I0_8_2_0 = I_8_2_0; // @[Top.scala 347:13]
  assign n143_I0_8_2_1 = I_8_2_1; // @[Top.scala 347:13]
  assign n143_I0_8_2_2 = I_8_2_2; // @[Top.scala 347:13]
  assign n143_I0_9_0_0 = I_9_0_0; // @[Top.scala 347:13]
  assign n143_I0_9_0_1 = I_9_0_1; // @[Top.scala 347:13]
  assign n143_I0_9_0_2 = I_9_0_2; // @[Top.scala 347:13]
  assign n143_I0_9_1_0 = I_9_1_0; // @[Top.scala 347:13]
  assign n143_I0_9_1_1 = I_9_1_1; // @[Top.scala 347:13]
  assign n143_I0_9_1_2 = I_9_1_2; // @[Top.scala 347:13]
  assign n143_I0_9_2_0 = I_9_2_0; // @[Top.scala 347:13]
  assign n143_I0_9_2_1 = I_9_2_1; // @[Top.scala 347:13]
  assign n143_I0_9_2_2 = I_9_2_2; // @[Top.scala 347:13]
  assign n143_I0_10_0_0 = I_10_0_0; // @[Top.scala 347:13]
  assign n143_I0_10_0_1 = I_10_0_1; // @[Top.scala 347:13]
  assign n143_I0_10_0_2 = I_10_0_2; // @[Top.scala 347:13]
  assign n143_I0_10_1_0 = I_10_1_0; // @[Top.scala 347:13]
  assign n143_I0_10_1_1 = I_10_1_1; // @[Top.scala 347:13]
  assign n143_I0_10_1_2 = I_10_1_2; // @[Top.scala 347:13]
  assign n143_I0_10_2_0 = I_10_2_0; // @[Top.scala 347:13]
  assign n143_I0_10_2_1 = I_10_2_1; // @[Top.scala 347:13]
  assign n143_I0_10_2_2 = I_10_2_2; // @[Top.scala 347:13]
  assign n143_I0_11_0_0 = I_11_0_0; // @[Top.scala 347:13]
  assign n143_I0_11_0_1 = I_11_0_1; // @[Top.scala 347:13]
  assign n143_I0_11_0_2 = I_11_0_2; // @[Top.scala 347:13]
  assign n143_I0_11_1_0 = I_11_1_0; // @[Top.scala 347:13]
  assign n143_I0_11_1_1 = I_11_1_1; // @[Top.scala 347:13]
  assign n143_I0_11_1_2 = I_11_1_2; // @[Top.scala 347:13]
  assign n143_I0_11_2_0 = I_11_2_0; // @[Top.scala 347:13]
  assign n143_I0_11_2_1 = I_11_2_1; // @[Top.scala 347:13]
  assign n143_I0_11_2_2 = I_11_2_2; // @[Top.scala 347:13]
  assign n143_I0_12_0_0 = I_12_0_0; // @[Top.scala 347:13]
  assign n143_I0_12_0_1 = I_12_0_1; // @[Top.scala 347:13]
  assign n143_I0_12_0_2 = I_12_0_2; // @[Top.scala 347:13]
  assign n143_I0_12_1_0 = I_12_1_0; // @[Top.scala 347:13]
  assign n143_I0_12_1_1 = I_12_1_1; // @[Top.scala 347:13]
  assign n143_I0_12_1_2 = I_12_1_2; // @[Top.scala 347:13]
  assign n143_I0_12_2_0 = I_12_2_0; // @[Top.scala 347:13]
  assign n143_I0_12_2_1 = I_12_2_1; // @[Top.scala 347:13]
  assign n143_I0_12_2_2 = I_12_2_2; // @[Top.scala 347:13]
  assign n143_I0_13_0_0 = I_13_0_0; // @[Top.scala 347:13]
  assign n143_I0_13_0_1 = I_13_0_1; // @[Top.scala 347:13]
  assign n143_I0_13_0_2 = I_13_0_2; // @[Top.scala 347:13]
  assign n143_I0_13_1_0 = I_13_1_0; // @[Top.scala 347:13]
  assign n143_I0_13_1_1 = I_13_1_1; // @[Top.scala 347:13]
  assign n143_I0_13_1_2 = I_13_1_2; // @[Top.scala 347:13]
  assign n143_I0_13_2_0 = I_13_2_0; // @[Top.scala 347:13]
  assign n143_I0_13_2_1 = I_13_2_1; // @[Top.scala 347:13]
  assign n143_I0_13_2_2 = I_13_2_2; // @[Top.scala 347:13]
  assign n143_I0_14_0_0 = I_14_0_0; // @[Top.scala 347:13]
  assign n143_I0_14_0_1 = I_14_0_1; // @[Top.scala 347:13]
  assign n143_I0_14_0_2 = I_14_0_2; // @[Top.scala 347:13]
  assign n143_I0_14_1_0 = I_14_1_0; // @[Top.scala 347:13]
  assign n143_I0_14_1_1 = I_14_1_1; // @[Top.scala 347:13]
  assign n143_I0_14_1_2 = I_14_1_2; // @[Top.scala 347:13]
  assign n143_I0_14_2_0 = I_14_2_0; // @[Top.scala 347:13]
  assign n143_I0_14_2_1 = I_14_2_1; // @[Top.scala 347:13]
  assign n143_I0_14_2_2 = I_14_2_2; // @[Top.scala 347:13]
  assign n143_I0_15_0_0 = I_15_0_0; // @[Top.scala 347:13]
  assign n143_I0_15_0_1 = I_15_0_1; // @[Top.scala 347:13]
  assign n143_I0_15_0_2 = I_15_0_2; // @[Top.scala 347:13]
  assign n143_I0_15_1_0 = I_15_1_0; // @[Top.scala 347:13]
  assign n143_I0_15_1_1 = I_15_1_1; // @[Top.scala 347:13]
  assign n143_I0_15_1_2 = I_15_1_2; // @[Top.scala 347:13]
  assign n143_I0_15_2_0 = I_15_2_0; // @[Top.scala 347:13]
  assign n143_I0_15_2_1 = I_15_2_1; // @[Top.scala 347:13]
  assign n143_I0_15_2_2 = I_15_2_2; // @[Top.scala 347:13]
  assign n143_I1_0_0_0_t0b = n142_O_0_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_0_0_0_t1b = n142_O_0_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_1_0_0_t0b = n142_O_1_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_1_0_0_t1b = n142_O_1_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_2_0_0_t0b = n142_O_2_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_2_0_0_t1b = n142_O_2_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_3_0_0_t0b = n142_O_3_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_3_0_0_t1b = n142_O_3_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_4_0_0_t0b = n142_O_4_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_4_0_0_t1b = n142_O_4_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_5_0_0_t0b = n142_O_5_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_5_0_0_t1b = n142_O_5_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_6_0_0_t0b = n142_O_6_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_6_0_0_t1b = n142_O_6_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_7_0_0_t0b = n142_O_7_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_7_0_0_t1b = n142_O_7_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_8_0_0_t0b = n142_O_8_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_8_0_0_t1b = n142_O_8_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_9_0_0_t0b = n142_O_9_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_9_0_0_t1b = n142_O_9_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_10_0_0_t0b = n142_O_10_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_10_0_0_t1b = n142_O_10_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_11_0_0_t0b = n142_O_11_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_11_0_0_t1b = n142_O_11_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_12_0_0_t0b = n142_O_12_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_12_0_0_t1b = n142_O_12_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_13_0_0_t0b = n142_O_13_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_13_0_0_t1b = n142_O_13_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_14_0_0_t0b = n142_O_14_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_14_0_0_t1b = n142_O_14_0_0_t1b; // @[Top.scala 348:13]
  assign n143_I1_15_0_0_t0b = n142_O_15_0_0_t0b; // @[Top.scala 348:13]
  assign n143_I1_15_0_0_t1b = n142_O_15_0_0_t1b; // @[Top.scala 348:13]
endmodule
module MapT_12(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0,
  input  [31:0] I_0_0_1,
  input  [31:0] I_0_0_2,
  input  [31:0] I_0_1_0,
  input  [31:0] I_0_1_1,
  input  [31:0] I_0_1_2,
  input  [31:0] I_0_2_0,
  input  [31:0] I_0_2_1,
  input  [31:0] I_0_2_2,
  input  [31:0] I_1_0_0,
  input  [31:0] I_1_0_1,
  input  [31:0] I_1_0_2,
  input  [31:0] I_1_1_0,
  input  [31:0] I_1_1_1,
  input  [31:0] I_1_1_2,
  input  [31:0] I_1_2_0,
  input  [31:0] I_1_2_1,
  input  [31:0] I_1_2_2,
  input  [31:0] I_2_0_0,
  input  [31:0] I_2_0_1,
  input  [31:0] I_2_0_2,
  input  [31:0] I_2_1_0,
  input  [31:0] I_2_1_1,
  input  [31:0] I_2_1_2,
  input  [31:0] I_2_2_0,
  input  [31:0] I_2_2_1,
  input  [31:0] I_2_2_2,
  input  [31:0] I_3_0_0,
  input  [31:0] I_3_0_1,
  input  [31:0] I_3_0_2,
  input  [31:0] I_3_1_0,
  input  [31:0] I_3_1_1,
  input  [31:0] I_3_1_2,
  input  [31:0] I_3_2_0,
  input  [31:0] I_3_2_1,
  input  [31:0] I_3_2_2,
  input  [31:0] I_4_0_0,
  input  [31:0] I_4_0_1,
  input  [31:0] I_4_0_2,
  input  [31:0] I_4_1_0,
  input  [31:0] I_4_1_1,
  input  [31:0] I_4_1_2,
  input  [31:0] I_4_2_0,
  input  [31:0] I_4_2_1,
  input  [31:0] I_4_2_2,
  input  [31:0] I_5_0_0,
  input  [31:0] I_5_0_1,
  input  [31:0] I_5_0_2,
  input  [31:0] I_5_1_0,
  input  [31:0] I_5_1_1,
  input  [31:0] I_5_1_2,
  input  [31:0] I_5_2_0,
  input  [31:0] I_5_2_1,
  input  [31:0] I_5_2_2,
  input  [31:0] I_6_0_0,
  input  [31:0] I_6_0_1,
  input  [31:0] I_6_0_2,
  input  [31:0] I_6_1_0,
  input  [31:0] I_6_1_1,
  input  [31:0] I_6_1_2,
  input  [31:0] I_6_2_0,
  input  [31:0] I_6_2_1,
  input  [31:0] I_6_2_2,
  input  [31:0] I_7_0_0,
  input  [31:0] I_7_0_1,
  input  [31:0] I_7_0_2,
  input  [31:0] I_7_1_0,
  input  [31:0] I_7_1_1,
  input  [31:0] I_7_1_2,
  input  [31:0] I_7_2_0,
  input  [31:0] I_7_2_1,
  input  [31:0] I_7_2_2,
  input  [31:0] I_8_0_0,
  input  [31:0] I_8_0_1,
  input  [31:0] I_8_0_2,
  input  [31:0] I_8_1_0,
  input  [31:0] I_8_1_1,
  input  [31:0] I_8_1_2,
  input  [31:0] I_8_2_0,
  input  [31:0] I_8_2_1,
  input  [31:0] I_8_2_2,
  input  [31:0] I_9_0_0,
  input  [31:0] I_9_0_1,
  input  [31:0] I_9_0_2,
  input  [31:0] I_9_1_0,
  input  [31:0] I_9_1_1,
  input  [31:0] I_9_1_2,
  input  [31:0] I_9_2_0,
  input  [31:0] I_9_2_1,
  input  [31:0] I_9_2_2,
  input  [31:0] I_10_0_0,
  input  [31:0] I_10_0_1,
  input  [31:0] I_10_0_2,
  input  [31:0] I_10_1_0,
  input  [31:0] I_10_1_1,
  input  [31:0] I_10_1_2,
  input  [31:0] I_10_2_0,
  input  [31:0] I_10_2_1,
  input  [31:0] I_10_2_2,
  input  [31:0] I_11_0_0,
  input  [31:0] I_11_0_1,
  input  [31:0] I_11_0_2,
  input  [31:0] I_11_1_0,
  input  [31:0] I_11_1_1,
  input  [31:0] I_11_1_2,
  input  [31:0] I_11_2_0,
  input  [31:0] I_11_2_1,
  input  [31:0] I_11_2_2,
  input  [31:0] I_12_0_0,
  input  [31:0] I_12_0_1,
  input  [31:0] I_12_0_2,
  input  [31:0] I_12_1_0,
  input  [31:0] I_12_1_1,
  input  [31:0] I_12_1_2,
  input  [31:0] I_12_2_0,
  input  [31:0] I_12_2_1,
  input  [31:0] I_12_2_2,
  input  [31:0] I_13_0_0,
  input  [31:0] I_13_0_1,
  input  [31:0] I_13_0_2,
  input  [31:0] I_13_1_0,
  input  [31:0] I_13_1_1,
  input  [31:0] I_13_1_2,
  input  [31:0] I_13_2_0,
  input  [31:0] I_13_2_1,
  input  [31:0] I_13_2_2,
  input  [31:0] I_14_0_0,
  input  [31:0] I_14_0_1,
  input  [31:0] I_14_0_2,
  input  [31:0] I_14_1_0,
  input  [31:0] I_14_1_1,
  input  [31:0] I_14_1_2,
  input  [31:0] I_14_2_0,
  input  [31:0] I_14_2_1,
  input  [31:0] I_14_2_2,
  input  [31:0] I_15_0_0,
  input  [31:0] I_15_0_1,
  input  [31:0] I_15_0_2,
  input  [31:0] I_15_1_0,
  input  [31:0] I_15_1_1,
  input  [31:0] I_15_1_2,
  input  [31:0] I_15_2_0,
  input  [31:0] I_15_2_1,
  input  [31:0] I_15_2_2,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b,
  output [31:0] O_8_0_0_t0b,
  output [31:0] O_8_0_0_t1b_t0b,
  output [31:0] O_8_0_0_t1b_t1b,
  output [31:0] O_9_0_0_t0b,
  output [31:0] O_9_0_0_t1b_t0b,
  output [31:0] O_9_0_0_t1b_t1b,
  output [31:0] O_10_0_0_t0b,
  output [31:0] O_10_0_0_t1b_t0b,
  output [31:0] O_10_0_0_t1b_t1b,
  output [31:0] O_11_0_0_t0b,
  output [31:0] O_11_0_0_t1b_t0b,
  output [31:0] O_11_0_0_t1b_t1b,
  output [31:0] O_12_0_0_t0b,
  output [31:0] O_12_0_0_t1b_t0b,
  output [31:0] O_12_0_0_t1b_t1b,
  output [31:0] O_13_0_0_t0b,
  output [31:0] O_13_0_0_t1b_t0b,
  output [31:0] O_13_0_0_t1b_t1b,
  output [31:0] O_14_0_0_t0b,
  output [31:0] O_14_0_0_t1b_t0b,
  output [31:0] O_14_0_0_t1b_t1b,
  output [31:0] O_15_0_0_t0b,
  output [31:0] O_15_0_0_t1b_t0b,
  output [31:0] O_15_0_0_t1b_t1b
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [31:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_0_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_1_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_2_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_3_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_4_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_5_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_6_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_7_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_8_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_9_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_10_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_11_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_12_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_13_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_14_0_0_t1b_t1b; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0_t1b_t0b; // @[MapT.scala 8:20]
  wire [31:0] op_O_15_0_0_t1b_t1b; // @[MapT.scala 8:20]
  Module_7 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0_t0b(op_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(op_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(op_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(op_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(op_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(op_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(op_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(op_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(op_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(op_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(op_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(op_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(op_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(op_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(op_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(op_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(op_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(op_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(op_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(op_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(op_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(op_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(op_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(op_O_7_0_0_t1b_t1b),
    .O_8_0_0_t0b(op_O_8_0_0_t0b),
    .O_8_0_0_t1b_t0b(op_O_8_0_0_t1b_t0b),
    .O_8_0_0_t1b_t1b(op_O_8_0_0_t1b_t1b),
    .O_9_0_0_t0b(op_O_9_0_0_t0b),
    .O_9_0_0_t1b_t0b(op_O_9_0_0_t1b_t0b),
    .O_9_0_0_t1b_t1b(op_O_9_0_0_t1b_t1b),
    .O_10_0_0_t0b(op_O_10_0_0_t0b),
    .O_10_0_0_t1b_t0b(op_O_10_0_0_t1b_t0b),
    .O_10_0_0_t1b_t1b(op_O_10_0_0_t1b_t1b),
    .O_11_0_0_t0b(op_O_11_0_0_t0b),
    .O_11_0_0_t1b_t0b(op_O_11_0_0_t1b_t0b),
    .O_11_0_0_t1b_t1b(op_O_11_0_0_t1b_t1b),
    .O_12_0_0_t0b(op_O_12_0_0_t0b),
    .O_12_0_0_t1b_t0b(op_O_12_0_0_t1b_t0b),
    .O_12_0_0_t1b_t1b(op_O_12_0_0_t1b_t1b),
    .O_13_0_0_t0b(op_O_13_0_0_t0b),
    .O_13_0_0_t1b_t0b(op_O_13_0_0_t1b_t0b),
    .O_13_0_0_t1b_t1b(op_O_13_0_0_t1b_t1b),
    .O_14_0_0_t0b(op_O_14_0_0_t0b),
    .O_14_0_0_t1b_t0b(op_O_14_0_0_t1b_t0b),
    .O_14_0_0_t1b_t1b(op_O_14_0_0_t1b_t1b),
    .O_15_0_0_t0b(op_O_15_0_0_t0b),
    .O_15_0_0_t1b_t0b(op_O_15_0_0_t1b_t0b),
    .O_15_0_0_t1b_t1b(op_O_15_0_0_t1b_t1b)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_t0b = op_O_0_0_0_t0b; // @[MapT.scala 15:7]
  assign O_0_0_0_t1b_t0b = op_O_0_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_0_0_0_t1b_t1b = op_O_0_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_1_0_0_t0b = op_O_1_0_0_t0b; // @[MapT.scala 15:7]
  assign O_1_0_0_t1b_t0b = op_O_1_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_1_0_0_t1b_t1b = op_O_1_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_2_0_0_t0b = op_O_2_0_0_t0b; // @[MapT.scala 15:7]
  assign O_2_0_0_t1b_t0b = op_O_2_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_2_0_0_t1b_t1b = op_O_2_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_3_0_0_t0b = op_O_3_0_0_t0b; // @[MapT.scala 15:7]
  assign O_3_0_0_t1b_t0b = op_O_3_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_3_0_0_t1b_t1b = op_O_3_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_4_0_0_t0b = op_O_4_0_0_t0b; // @[MapT.scala 15:7]
  assign O_4_0_0_t1b_t0b = op_O_4_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_4_0_0_t1b_t1b = op_O_4_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_5_0_0_t0b = op_O_5_0_0_t0b; // @[MapT.scala 15:7]
  assign O_5_0_0_t1b_t0b = op_O_5_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_5_0_0_t1b_t1b = op_O_5_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_6_0_0_t0b = op_O_6_0_0_t0b; // @[MapT.scala 15:7]
  assign O_6_0_0_t1b_t0b = op_O_6_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_6_0_0_t1b_t1b = op_O_6_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_7_0_0_t0b = op_O_7_0_0_t0b; // @[MapT.scala 15:7]
  assign O_7_0_0_t1b_t0b = op_O_7_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_7_0_0_t1b_t1b = op_O_7_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_8_0_0_t0b = op_O_8_0_0_t0b; // @[MapT.scala 15:7]
  assign O_8_0_0_t1b_t0b = op_O_8_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_8_0_0_t1b_t1b = op_O_8_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_9_0_0_t0b = op_O_9_0_0_t0b; // @[MapT.scala 15:7]
  assign O_9_0_0_t1b_t0b = op_O_9_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_9_0_0_t1b_t1b = op_O_9_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_10_0_0_t0b = op_O_10_0_0_t0b; // @[MapT.scala 15:7]
  assign O_10_0_0_t1b_t0b = op_O_10_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_10_0_0_t1b_t1b = op_O_10_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_11_0_0_t0b = op_O_11_0_0_t0b; // @[MapT.scala 15:7]
  assign O_11_0_0_t1b_t0b = op_O_11_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_11_0_0_t1b_t1b = op_O_11_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_12_0_0_t0b = op_O_12_0_0_t0b; // @[MapT.scala 15:7]
  assign O_12_0_0_t1b_t0b = op_O_12_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_12_0_0_t1b_t1b = op_O_12_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_13_0_0_t0b = op_O_13_0_0_t0b; // @[MapT.scala 15:7]
  assign O_13_0_0_t1b_t0b = op_O_13_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_13_0_0_t1b_t1b = op_O_13_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_14_0_0_t0b = op_O_14_0_0_t0b; // @[MapT.scala 15:7]
  assign O_14_0_0_t1b_t0b = op_O_14_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_14_0_0_t1b_t1b = op_O_14_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign O_15_0_0_t0b = op_O_15_0_0_t0b; // @[MapT.scala 15:7]
  assign O_15_0_0_t1b_t0b = op_O_15_0_0_t1b_t0b; // @[MapT.scala 15:7]
  assign O_15_0_0_t1b_t1b = op_O_15_0_0_t1b_t1b; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough_1(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_t0b,
  input  [31:0] I_0_0_0_t1b_t0b,
  input  [31:0] I_0_0_0_t1b_t1b,
  input  [31:0] I_1_0_0_t0b,
  input  [31:0] I_1_0_0_t1b_t0b,
  input  [31:0] I_1_0_0_t1b_t1b,
  input  [31:0] I_2_0_0_t0b,
  input  [31:0] I_2_0_0_t1b_t0b,
  input  [31:0] I_2_0_0_t1b_t1b,
  input  [31:0] I_3_0_0_t0b,
  input  [31:0] I_3_0_0_t1b_t0b,
  input  [31:0] I_3_0_0_t1b_t1b,
  input  [31:0] I_4_0_0_t0b,
  input  [31:0] I_4_0_0_t1b_t0b,
  input  [31:0] I_4_0_0_t1b_t1b,
  input  [31:0] I_5_0_0_t0b,
  input  [31:0] I_5_0_0_t1b_t0b,
  input  [31:0] I_5_0_0_t1b_t1b,
  input  [31:0] I_6_0_0_t0b,
  input  [31:0] I_6_0_0_t1b_t0b,
  input  [31:0] I_6_0_0_t1b_t1b,
  input  [31:0] I_7_0_0_t0b,
  input  [31:0] I_7_0_0_t1b_t0b,
  input  [31:0] I_7_0_0_t1b_t1b,
  input  [31:0] I_8_0_0_t0b,
  input  [31:0] I_8_0_0_t1b_t0b,
  input  [31:0] I_8_0_0_t1b_t1b,
  input  [31:0] I_9_0_0_t0b,
  input  [31:0] I_9_0_0_t1b_t0b,
  input  [31:0] I_9_0_0_t1b_t1b,
  input  [31:0] I_10_0_0_t0b,
  input  [31:0] I_10_0_0_t1b_t0b,
  input  [31:0] I_10_0_0_t1b_t1b,
  input  [31:0] I_11_0_0_t0b,
  input  [31:0] I_11_0_0_t1b_t0b,
  input  [31:0] I_11_0_0_t1b_t1b,
  input  [31:0] I_12_0_0_t0b,
  input  [31:0] I_12_0_0_t1b_t0b,
  input  [31:0] I_12_0_0_t1b_t1b,
  input  [31:0] I_13_0_0_t0b,
  input  [31:0] I_13_0_0_t1b_t0b,
  input  [31:0] I_13_0_0_t1b_t1b,
  input  [31:0] I_14_0_0_t0b,
  input  [31:0] I_14_0_0_t1b_t0b,
  input  [31:0] I_14_0_0_t1b_t1b,
  input  [31:0] I_15_0_0_t0b,
  input  [31:0] I_15_0_0_t1b_t0b,
  input  [31:0] I_15_0_0_t1b_t1b,
  output [31:0] O_0_0_0_t0b,
  output [31:0] O_0_0_0_t1b_t0b,
  output [31:0] O_0_0_0_t1b_t1b,
  output [31:0] O_1_0_0_t0b,
  output [31:0] O_1_0_0_t1b_t0b,
  output [31:0] O_1_0_0_t1b_t1b,
  output [31:0] O_2_0_0_t0b,
  output [31:0] O_2_0_0_t1b_t0b,
  output [31:0] O_2_0_0_t1b_t1b,
  output [31:0] O_3_0_0_t0b,
  output [31:0] O_3_0_0_t1b_t0b,
  output [31:0] O_3_0_0_t1b_t1b,
  output [31:0] O_4_0_0_t0b,
  output [31:0] O_4_0_0_t1b_t0b,
  output [31:0] O_4_0_0_t1b_t1b,
  output [31:0] O_5_0_0_t0b,
  output [31:0] O_5_0_0_t1b_t0b,
  output [31:0] O_5_0_0_t1b_t1b,
  output [31:0] O_6_0_0_t0b,
  output [31:0] O_6_0_0_t1b_t0b,
  output [31:0] O_6_0_0_t1b_t1b,
  output [31:0] O_7_0_0_t0b,
  output [31:0] O_7_0_0_t1b_t0b,
  output [31:0] O_7_0_0_t1b_t1b,
  output [31:0] O_8_0_0_t0b,
  output [31:0] O_8_0_0_t1b_t0b,
  output [31:0] O_8_0_0_t1b_t1b,
  output [31:0] O_9_0_0_t0b,
  output [31:0] O_9_0_0_t1b_t0b,
  output [31:0] O_9_0_0_t1b_t1b,
  output [31:0] O_10_0_0_t0b,
  output [31:0] O_10_0_0_t1b_t0b,
  output [31:0] O_10_0_0_t1b_t1b,
  output [31:0] O_11_0_0_t0b,
  output [31:0] O_11_0_0_t1b_t0b,
  output [31:0] O_11_0_0_t1b_t1b,
  output [31:0] O_12_0_0_t0b,
  output [31:0] O_12_0_0_t1b_t0b,
  output [31:0] O_12_0_0_t1b_t1b,
  output [31:0] O_13_0_0_t0b,
  output [31:0] O_13_0_0_t1b_t0b,
  output [31:0] O_13_0_0_t1b_t1b,
  output [31:0] O_14_0_0_t0b,
  output [31:0] O_14_0_0_t1b_t0b,
  output [31:0] O_14_0_0_t1b_t1b,
  output [31:0] O_15_0_0_t0b,
  output [31:0] O_15_0_0_t1b_t0b,
  output [31:0] O_15_0_0_t1b_t1b
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0_0_t0b = I_0_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_0_t1b_t0b = I_0_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_0_t1b_t1b = I_0_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_1_0_0_t0b = I_1_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_0_t1b_t0b = I_1_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_0_t1b_t1b = I_1_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_2_0_0_t0b = I_2_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_0_t1b_t0b = I_2_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_0_t1b_t1b = I_2_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_3_0_0_t0b = I_3_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_0_t1b_t0b = I_3_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_0_t1b_t1b = I_3_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_4_0_0_t0b = I_4_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_0_t1b_t0b = I_4_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_0_t1b_t1b = I_4_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_5_0_0_t0b = I_5_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_0_t1b_t0b = I_5_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_0_t1b_t1b = I_5_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_6_0_0_t0b = I_6_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_0_t1b_t0b = I_6_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_0_t1b_t1b = I_6_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_7_0_0_t0b = I_7_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_0_t1b_t0b = I_7_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_0_t1b_t1b = I_7_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_8_0_0_t0b = I_8_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_8_0_0_t1b_t0b = I_8_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_8_0_0_t1b_t1b = I_8_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_9_0_0_t0b = I_9_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_9_0_0_t1b_t0b = I_9_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_9_0_0_t1b_t1b = I_9_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_10_0_0_t0b = I_10_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_10_0_0_t1b_t0b = I_10_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_10_0_0_t1b_t1b = I_10_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_11_0_0_t0b = I_11_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_11_0_0_t1b_t0b = I_11_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_11_0_0_t1b_t1b = I_11_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_12_0_0_t0b = I_12_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_12_0_0_t1b_t0b = I_12_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_12_0_0_t1b_t1b = I_12_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_13_0_0_t0b = I_13_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_13_0_0_t1b_t0b = I_13_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_13_0_0_t1b_t1b = I_13_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_14_0_0_t0b = I_14_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_14_0_0_t1b_t0b = I_14_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_14_0_0_t1b_t1b = I_14_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_15_0_0_t0b = I_15_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_15_0_0_t1b_t0b = I_15_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_15_0_0_t1b_t1b = I_15_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_2(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_0_t0b,
  input  [31:0] I_0_0_0_t1b_t0b,
  input  [31:0] I_0_0_0_t1b_t1b,
  input  [31:0] I_1_0_0_t0b,
  input  [31:0] I_1_0_0_t1b_t0b,
  input  [31:0] I_1_0_0_t1b_t1b,
  input  [31:0] I_2_0_0_t0b,
  input  [31:0] I_2_0_0_t1b_t0b,
  input  [31:0] I_2_0_0_t1b_t1b,
  input  [31:0] I_3_0_0_t0b,
  input  [31:0] I_3_0_0_t1b_t0b,
  input  [31:0] I_3_0_0_t1b_t1b,
  input  [31:0] I_4_0_0_t0b,
  input  [31:0] I_4_0_0_t1b_t0b,
  input  [31:0] I_4_0_0_t1b_t1b,
  input  [31:0] I_5_0_0_t0b,
  input  [31:0] I_5_0_0_t1b_t0b,
  input  [31:0] I_5_0_0_t1b_t1b,
  input  [31:0] I_6_0_0_t0b,
  input  [31:0] I_6_0_0_t1b_t0b,
  input  [31:0] I_6_0_0_t1b_t1b,
  input  [31:0] I_7_0_0_t0b,
  input  [31:0] I_7_0_0_t1b_t0b,
  input  [31:0] I_7_0_0_t1b_t1b,
  input  [31:0] I_8_0_0_t0b,
  input  [31:0] I_8_0_0_t1b_t0b,
  input  [31:0] I_8_0_0_t1b_t1b,
  input  [31:0] I_9_0_0_t0b,
  input  [31:0] I_9_0_0_t1b_t0b,
  input  [31:0] I_9_0_0_t1b_t1b,
  input  [31:0] I_10_0_0_t0b,
  input  [31:0] I_10_0_0_t1b_t0b,
  input  [31:0] I_10_0_0_t1b_t1b,
  input  [31:0] I_11_0_0_t0b,
  input  [31:0] I_11_0_0_t1b_t0b,
  input  [31:0] I_11_0_0_t1b_t1b,
  input  [31:0] I_12_0_0_t0b,
  input  [31:0] I_12_0_0_t1b_t0b,
  input  [31:0] I_12_0_0_t1b_t1b,
  input  [31:0] I_13_0_0_t0b,
  input  [31:0] I_13_0_0_t1b_t0b,
  input  [31:0] I_13_0_0_t1b_t1b,
  input  [31:0] I_14_0_0_t0b,
  input  [31:0] I_14_0_0_t1b_t0b,
  input  [31:0] I_14_0_0_t1b_t1b,
  input  [31:0] I_15_0_0_t0b,
  input  [31:0] I_15_0_0_t1b_t0b,
  input  [31:0] I_15_0_0_t1b_t1b,
  output [31:0] O_0_0_t0b,
  output [31:0] O_0_0_t1b_t0b,
  output [31:0] O_0_0_t1b_t1b,
  output [31:0] O_1_0_t0b,
  output [31:0] O_1_0_t1b_t0b,
  output [31:0] O_1_0_t1b_t1b,
  output [31:0] O_2_0_t0b,
  output [31:0] O_2_0_t1b_t0b,
  output [31:0] O_2_0_t1b_t1b,
  output [31:0] O_3_0_t0b,
  output [31:0] O_3_0_t1b_t0b,
  output [31:0] O_3_0_t1b_t1b,
  output [31:0] O_4_0_t0b,
  output [31:0] O_4_0_t1b_t0b,
  output [31:0] O_4_0_t1b_t1b,
  output [31:0] O_5_0_t0b,
  output [31:0] O_5_0_t1b_t0b,
  output [31:0] O_5_0_t1b_t1b,
  output [31:0] O_6_0_t0b,
  output [31:0] O_6_0_t1b_t0b,
  output [31:0] O_6_0_t1b_t1b,
  output [31:0] O_7_0_t0b,
  output [31:0] O_7_0_t1b_t0b,
  output [31:0] O_7_0_t1b_t1b,
  output [31:0] O_8_0_t0b,
  output [31:0] O_8_0_t1b_t0b,
  output [31:0] O_8_0_t1b_t1b,
  output [31:0] O_9_0_t0b,
  output [31:0] O_9_0_t1b_t0b,
  output [31:0] O_9_0_t1b_t1b,
  output [31:0] O_10_0_t0b,
  output [31:0] O_10_0_t1b_t0b,
  output [31:0] O_10_0_t1b_t1b,
  output [31:0] O_11_0_t0b,
  output [31:0] O_11_0_t1b_t0b,
  output [31:0] O_11_0_t1b_t1b,
  output [31:0] O_12_0_t0b,
  output [31:0] O_12_0_t1b_t0b,
  output [31:0] O_12_0_t1b_t1b,
  output [31:0] O_13_0_t0b,
  output [31:0] O_13_0_t1b_t0b,
  output [31:0] O_13_0_t1b_t1b,
  output [31:0] O_14_0_t0b,
  output [31:0] O_14_0_t1b_t0b,
  output [31:0] O_14_0_t1b_t1b,
  output [31:0] O_15_0_t0b,
  output [31:0] O_15_0_t1b_t0b,
  output [31:0] O_15_0_t1b_t1b
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0_t0b = I_0_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_t1b_t0b = I_0_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_0_0_t1b_t1b = I_0_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_1_0_t0b = I_1_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_t1b_t0b = I_1_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_1_0_t1b_t1b = I_1_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_2_0_t0b = I_2_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_t1b_t0b = I_2_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_2_0_t1b_t1b = I_2_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_3_0_t0b = I_3_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_t1b_t0b = I_3_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_3_0_t1b_t1b = I_3_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_4_0_t0b = I_4_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_t1b_t0b = I_4_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_4_0_t1b_t1b = I_4_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_5_0_t0b = I_5_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_t1b_t0b = I_5_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_5_0_t1b_t1b = I_5_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_6_0_t0b = I_6_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_t1b_t0b = I_6_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_6_0_t1b_t1b = I_6_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_7_0_t0b = I_7_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_t1b_t0b = I_7_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_7_0_t1b_t1b = I_7_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_8_0_t0b = I_8_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_8_0_t1b_t0b = I_8_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_8_0_t1b_t1b = I_8_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_9_0_t0b = I_9_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_9_0_t1b_t0b = I_9_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_9_0_t1b_t1b = I_9_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_10_0_t0b = I_10_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_10_0_t1b_t0b = I_10_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_10_0_t1b_t1b = I_10_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_11_0_t0b = I_11_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_11_0_t1b_t0b = I_11_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_11_0_t1b_t1b = I_11_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_12_0_t0b = I_12_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_12_0_t1b_t0b = I_12_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_12_0_t1b_t1b = I_12_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_13_0_t0b = I_13_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_13_0_t1b_t0b = I_13_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_13_0_t1b_t1b = I_13_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_14_0_t0b = I_14_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_14_0_t1b_t0b = I_14_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_14_0_t1b_t1b = I_14_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_15_0_t0b = I_15_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_15_0_t1b_t0b = I_15_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_15_0_t1b_t1b = I_15_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_3(
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_0_t0b,
  input  [31:0] I_0_0_t1b_t0b,
  input  [31:0] I_0_0_t1b_t1b,
  input  [31:0] I_1_0_t0b,
  input  [31:0] I_1_0_t1b_t0b,
  input  [31:0] I_1_0_t1b_t1b,
  input  [31:0] I_2_0_t0b,
  input  [31:0] I_2_0_t1b_t0b,
  input  [31:0] I_2_0_t1b_t1b,
  input  [31:0] I_3_0_t0b,
  input  [31:0] I_3_0_t1b_t0b,
  input  [31:0] I_3_0_t1b_t1b,
  input  [31:0] I_4_0_t0b,
  input  [31:0] I_4_0_t1b_t0b,
  input  [31:0] I_4_0_t1b_t1b,
  input  [31:0] I_5_0_t0b,
  input  [31:0] I_5_0_t1b_t0b,
  input  [31:0] I_5_0_t1b_t1b,
  input  [31:0] I_6_0_t0b,
  input  [31:0] I_6_0_t1b_t0b,
  input  [31:0] I_6_0_t1b_t1b,
  input  [31:0] I_7_0_t0b,
  input  [31:0] I_7_0_t1b_t0b,
  input  [31:0] I_7_0_t1b_t1b,
  input  [31:0] I_8_0_t0b,
  input  [31:0] I_8_0_t1b_t0b,
  input  [31:0] I_8_0_t1b_t1b,
  input  [31:0] I_9_0_t0b,
  input  [31:0] I_9_0_t1b_t0b,
  input  [31:0] I_9_0_t1b_t1b,
  input  [31:0] I_10_0_t0b,
  input  [31:0] I_10_0_t1b_t0b,
  input  [31:0] I_10_0_t1b_t1b,
  input  [31:0] I_11_0_t0b,
  input  [31:0] I_11_0_t1b_t0b,
  input  [31:0] I_11_0_t1b_t1b,
  input  [31:0] I_12_0_t0b,
  input  [31:0] I_12_0_t1b_t0b,
  input  [31:0] I_12_0_t1b_t1b,
  input  [31:0] I_13_0_t0b,
  input  [31:0] I_13_0_t1b_t0b,
  input  [31:0] I_13_0_t1b_t1b,
  input  [31:0] I_14_0_t0b,
  input  [31:0] I_14_0_t1b_t0b,
  input  [31:0] I_14_0_t1b_t1b,
  input  [31:0] I_15_0_t0b,
  input  [31:0] I_15_0_t1b_t0b,
  input  [31:0] I_15_0_t1b_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b,
  output [31:0] O_8_t0b,
  output [31:0] O_8_t1b_t0b,
  output [31:0] O_8_t1b_t1b,
  output [31:0] O_9_t0b,
  output [31:0] O_9_t1b_t0b,
  output [31:0] O_9_t1b_t1b,
  output [31:0] O_10_t0b,
  output [31:0] O_10_t1b_t0b,
  output [31:0] O_10_t1b_t1b,
  output [31:0] O_11_t0b,
  output [31:0] O_11_t1b_t0b,
  output [31:0] O_11_t1b_t1b,
  output [31:0] O_12_t0b,
  output [31:0] O_12_t1b_t0b,
  output [31:0] O_12_t1b_t1b,
  output [31:0] O_13_t0b,
  output [31:0] O_13_t1b_t0b,
  output [31:0] O_13_t1b_t1b,
  output [31:0] O_14_t0b,
  output [31:0] O_14_t1b_t0b,
  output [31:0] O_14_t1b_t1b,
  output [31:0] O_15_t0b,
  output [31:0] O_15_t1b_t0b,
  output [31:0] O_15_t1b_t1b
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_t0b = I_0_0_t0b; // @[Passthrough.scala 17:68]
  assign O_0_t1b_t0b = I_0_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_0_t1b_t1b = I_0_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_1_t0b = I_1_0_t0b; // @[Passthrough.scala 17:68]
  assign O_1_t1b_t0b = I_1_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_1_t1b_t1b = I_1_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_2_t0b = I_2_0_t0b; // @[Passthrough.scala 17:68]
  assign O_2_t1b_t0b = I_2_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_2_t1b_t1b = I_2_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_3_t0b = I_3_0_t0b; // @[Passthrough.scala 17:68]
  assign O_3_t1b_t0b = I_3_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_3_t1b_t1b = I_3_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_4_t0b = I_4_0_t0b; // @[Passthrough.scala 17:68]
  assign O_4_t1b_t0b = I_4_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_4_t1b_t1b = I_4_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_5_t0b = I_5_0_t0b; // @[Passthrough.scala 17:68]
  assign O_5_t1b_t0b = I_5_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_5_t1b_t1b = I_5_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_6_t0b = I_6_0_t0b; // @[Passthrough.scala 17:68]
  assign O_6_t1b_t0b = I_6_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_6_t1b_t1b = I_6_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_7_t0b = I_7_0_t0b; // @[Passthrough.scala 17:68]
  assign O_7_t1b_t0b = I_7_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_7_t1b_t1b = I_7_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_8_t0b = I_8_0_t0b; // @[Passthrough.scala 17:68]
  assign O_8_t1b_t0b = I_8_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_8_t1b_t1b = I_8_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_9_t0b = I_9_0_t0b; // @[Passthrough.scala 17:68]
  assign O_9_t1b_t0b = I_9_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_9_t1b_t1b = I_9_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_10_t0b = I_10_0_t0b; // @[Passthrough.scala 17:68]
  assign O_10_t1b_t0b = I_10_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_10_t1b_t1b = I_10_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_11_t0b = I_11_0_t0b; // @[Passthrough.scala 17:68]
  assign O_11_t1b_t0b = I_11_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_11_t1b_t1b = I_11_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_12_t0b = I_12_0_t0b; // @[Passthrough.scala 17:68]
  assign O_12_t1b_t0b = I_12_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_12_t1b_t1b = I_12_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_13_t0b = I_13_0_t0b; // @[Passthrough.scala 17:68]
  assign O_13_t1b_t0b = I_13_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_13_t1b_t1b = I_13_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_14_t0b = I_14_0_t0b; // @[Passthrough.scala 17:68]
  assign O_14_t1b_t0b = I_14_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_14_t1b_t1b = I_14_0_t1b_t1b; // @[Passthrough.scala 17:68]
  assign O_15_t0b = I_15_0_t0b; // @[Passthrough.scala 17:68]
  assign O_15_t1b_t0b = I_15_0_t1b_t0b; // @[Passthrough.scala 17:68]
  assign O_15_t1b_t1b = I_15_0_t1b_t1b; // @[Passthrough.scala 17:68]
endmodule
module FIFO_9(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0_t0b,
  input  [31:0] I_0_t1b_t0b,
  input  [31:0] I_0_t1b_t1b,
  input  [31:0] I_1_t0b,
  input  [31:0] I_1_t1b_t0b,
  input  [31:0] I_1_t1b_t1b,
  input  [31:0] I_2_t0b,
  input  [31:0] I_2_t1b_t0b,
  input  [31:0] I_2_t1b_t1b,
  input  [31:0] I_3_t0b,
  input  [31:0] I_3_t1b_t0b,
  input  [31:0] I_3_t1b_t1b,
  input  [31:0] I_4_t0b,
  input  [31:0] I_4_t1b_t0b,
  input  [31:0] I_4_t1b_t1b,
  input  [31:0] I_5_t0b,
  input  [31:0] I_5_t1b_t0b,
  input  [31:0] I_5_t1b_t1b,
  input  [31:0] I_6_t0b,
  input  [31:0] I_6_t1b_t0b,
  input  [31:0] I_6_t1b_t1b,
  input  [31:0] I_7_t0b,
  input  [31:0] I_7_t1b_t0b,
  input  [31:0] I_7_t1b_t1b,
  input  [31:0] I_8_t0b,
  input  [31:0] I_8_t1b_t0b,
  input  [31:0] I_8_t1b_t1b,
  input  [31:0] I_9_t0b,
  input  [31:0] I_9_t1b_t0b,
  input  [31:0] I_9_t1b_t1b,
  input  [31:0] I_10_t0b,
  input  [31:0] I_10_t1b_t0b,
  input  [31:0] I_10_t1b_t1b,
  input  [31:0] I_11_t0b,
  input  [31:0] I_11_t1b_t0b,
  input  [31:0] I_11_t1b_t1b,
  input  [31:0] I_12_t0b,
  input  [31:0] I_12_t1b_t0b,
  input  [31:0] I_12_t1b_t1b,
  input  [31:0] I_13_t0b,
  input  [31:0] I_13_t1b_t0b,
  input  [31:0] I_13_t1b_t1b,
  input  [31:0] I_14_t0b,
  input  [31:0] I_14_t1b_t0b,
  input  [31:0] I_14_t1b_t1b,
  input  [31:0] I_15_t0b,
  input  [31:0] I_15_t1b_t0b,
  input  [31:0] I_15_t1b_t1b,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b,
  output [31:0] O_8_t0b,
  output [31:0] O_8_t1b_t0b,
  output [31:0] O_8_t1b_t1b,
  output [31:0] O_9_t0b,
  output [31:0] O_9_t1b_t0b,
  output [31:0] O_9_t1b_t1b,
  output [31:0] O_10_t0b,
  output [31:0] O_10_t1b_t0b,
  output [31:0] O_10_t1b_t1b,
  output [31:0] O_11_t0b,
  output [31:0] O_11_t1b_t0b,
  output [31:0] O_11_t1b_t1b,
  output [31:0] O_12_t0b,
  output [31:0] O_12_t1b_t0b,
  output [31:0] O_12_t1b_t1b,
  output [31:0] O_13_t0b,
  output [31:0] O_13_t1b_t0b,
  output [31:0] O_13_t1b_t1b,
  output [31:0] O_14_t0b,
  output [31:0] O_14_t1b_t0b,
  output [31:0] O_14_t1b_t1b,
  output [31:0] O_15_t0b,
  output [31:0] O_15_t1b_t0b,
  output [31:0] O_15_t1b_t1b
);
  reg [31:0] _T__0_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [31:0] _T__0_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [31:0] _T__0_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [31:0] _T__1_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [31:0] _T__1_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [31:0] _T__1_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [31:0] _T__2_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [31:0] _T__2_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [31:0] _T__2_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [31:0] _T__3_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [31:0] _T__3_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [31:0] _T__3_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [31:0] _T__4_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [31:0] _T__4_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [31:0] _T__4_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [31:0] _T__5_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg [31:0] _T__5_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_16;
  reg [31:0] _T__5_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_17;
  reg [31:0] _T__6_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_18;
  reg [31:0] _T__6_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_19;
  reg [31:0] _T__6_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_20;
  reg [31:0] _T__7_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_21;
  reg [31:0] _T__7_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_22;
  reg [31:0] _T__7_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_23;
  reg [31:0] _T__8_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_24;
  reg [31:0] _T__8_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_25;
  reg [31:0] _T__8_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_26;
  reg [31:0] _T__9_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_27;
  reg [31:0] _T__9_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_28;
  reg [31:0] _T__9_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_29;
  reg [31:0] _T__10_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_30;
  reg [31:0] _T__10_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_31;
  reg [31:0] _T__10_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_32;
  reg [31:0] _T__11_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_33;
  reg [31:0] _T__11_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_34;
  reg [31:0] _T__11_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_35;
  reg [31:0] _T__12_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_36;
  reg [31:0] _T__12_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_37;
  reg [31:0] _T__12_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_38;
  reg [31:0] _T__13_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_39;
  reg [31:0] _T__13_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_40;
  reg [31:0] _T__13_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_41;
  reg [31:0] _T__14_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_42;
  reg [31:0] _T__14_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_43;
  reg [31:0] _T__14_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_44;
  reg [31:0] _T__15_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_45;
  reg [31:0] _T__15_t1b_t0b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_46;
  reg [31:0] _T__15_t1b_t1b; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_47;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_48;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0_t0b = _T__0_t0b; // @[FIFO.scala 14:7]
  assign O_0_t1b_t0b = _T__0_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_0_t1b_t1b = _T__0_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_1_t0b = _T__1_t0b; // @[FIFO.scala 14:7]
  assign O_1_t1b_t0b = _T__1_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_1_t1b_t1b = _T__1_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_2_t0b = _T__2_t0b; // @[FIFO.scala 14:7]
  assign O_2_t1b_t0b = _T__2_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_2_t1b_t1b = _T__2_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_3_t0b = _T__3_t0b; // @[FIFO.scala 14:7]
  assign O_3_t1b_t0b = _T__3_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_3_t1b_t1b = _T__3_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_4_t0b = _T__4_t0b; // @[FIFO.scala 14:7]
  assign O_4_t1b_t0b = _T__4_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_4_t1b_t1b = _T__4_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_5_t0b = _T__5_t0b; // @[FIFO.scala 14:7]
  assign O_5_t1b_t0b = _T__5_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_5_t1b_t1b = _T__5_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_6_t0b = _T__6_t0b; // @[FIFO.scala 14:7]
  assign O_6_t1b_t0b = _T__6_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_6_t1b_t1b = _T__6_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_7_t0b = _T__7_t0b; // @[FIFO.scala 14:7]
  assign O_7_t1b_t0b = _T__7_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_7_t1b_t1b = _T__7_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_8_t0b = _T__8_t0b; // @[FIFO.scala 14:7]
  assign O_8_t1b_t0b = _T__8_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_8_t1b_t1b = _T__8_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_9_t0b = _T__9_t0b; // @[FIFO.scala 14:7]
  assign O_9_t1b_t0b = _T__9_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_9_t1b_t1b = _T__9_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_10_t0b = _T__10_t0b; // @[FIFO.scala 14:7]
  assign O_10_t1b_t0b = _T__10_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_10_t1b_t1b = _T__10_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_11_t0b = _T__11_t0b; // @[FIFO.scala 14:7]
  assign O_11_t1b_t0b = _T__11_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_11_t1b_t1b = _T__11_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_12_t0b = _T__12_t0b; // @[FIFO.scala 14:7]
  assign O_12_t1b_t0b = _T__12_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_12_t1b_t1b = _T__12_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_13_t0b = _T__13_t0b; // @[FIFO.scala 14:7]
  assign O_13_t1b_t0b = _T__13_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_13_t1b_t1b = _T__13_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_14_t0b = _T__14_t0b; // @[FIFO.scala 14:7]
  assign O_14_t1b_t0b = _T__14_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_14_t1b_t1b = _T__14_t1b_t1b; // @[FIFO.scala 14:7]
  assign O_15_t0b = _T__15_t0b; // @[FIFO.scala 14:7]
  assign O_15_t1b_t0b = _T__15_t1b_t0b; // @[FIFO.scala 14:7]
  assign O_15_t1b_t1b = _T__15_t1b_t1b; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0_t0b = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__0_t1b_t0b = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0_t1b_t1b = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__1_t0b = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__1_t1b_t0b = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__1_t1b_t1b = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__2_t0b = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__2_t1b_t0b = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__2_t1b_t1b = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__3_t0b = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__3_t1b_t0b = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__3_t1b_t1b = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__4_t0b = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__4_t1b_t0b = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__4_t1b_t1b = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__5_t0b = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T__5_t1b_t0b = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T__5_t1b_t1b = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__6_t0b = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__6_t1b_t0b = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T__6_t1b_t1b = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T__7_t0b = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__7_t1b_t0b = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__7_t1b_t1b = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T__8_t0b = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T__8_t1b_t0b = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__8_t1b_t1b = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__9_t0b = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T__9_t1b_t0b = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T__9_t1b_t1b = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__10_t0b = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__10_t1b_t0b = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T__10_t1b_t1b = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T__11_t0b = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__11_t1b_t0b = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__11_t1b_t1b = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T__12_t0b = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T__12_t1b_t0b = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__12_t1b_t1b = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__13_t0b = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T__13_t1b_t0b = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T__13_t1b_t1b = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__14_t0b = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__14_t1b_t0b = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T__14_t1b_t1b = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T__15_t0b = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__15_t1b_t0b = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__15_t1b_t1b = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0_t0b <= I_0_t0b;
    _T__0_t1b_t0b <= I_0_t1b_t0b;
    _T__0_t1b_t1b <= I_0_t1b_t1b;
    _T__1_t0b <= I_1_t0b;
    _T__1_t1b_t0b <= I_1_t1b_t0b;
    _T__1_t1b_t1b <= I_1_t1b_t1b;
    _T__2_t0b <= I_2_t0b;
    _T__2_t1b_t0b <= I_2_t1b_t0b;
    _T__2_t1b_t1b <= I_2_t1b_t1b;
    _T__3_t0b <= I_3_t0b;
    _T__3_t1b_t0b <= I_3_t1b_t0b;
    _T__3_t1b_t1b <= I_3_t1b_t1b;
    _T__4_t0b <= I_4_t0b;
    _T__4_t1b_t0b <= I_4_t1b_t0b;
    _T__4_t1b_t1b <= I_4_t1b_t1b;
    _T__5_t0b <= I_5_t0b;
    _T__5_t1b_t0b <= I_5_t1b_t0b;
    _T__5_t1b_t1b <= I_5_t1b_t1b;
    _T__6_t0b <= I_6_t0b;
    _T__6_t1b_t0b <= I_6_t1b_t0b;
    _T__6_t1b_t1b <= I_6_t1b_t1b;
    _T__7_t0b <= I_7_t0b;
    _T__7_t1b_t0b <= I_7_t1b_t0b;
    _T__7_t1b_t1b <= I_7_t1b_t1b;
    _T__8_t0b <= I_8_t0b;
    _T__8_t1b_t0b <= I_8_t1b_t0b;
    _T__8_t1b_t1b <= I_8_t1b_t1b;
    _T__9_t0b <= I_9_t0b;
    _T__9_t1b_t0b <= I_9_t1b_t0b;
    _T__9_t1b_t1b <= I_9_t1b_t1b;
    _T__10_t0b <= I_10_t0b;
    _T__10_t1b_t0b <= I_10_t1b_t0b;
    _T__10_t1b_t1b <= I_10_t1b_t1b;
    _T__11_t0b <= I_11_t0b;
    _T__11_t1b_t0b <= I_11_t1b_t0b;
    _T__11_t1b_t1b <= I_11_t1b_t1b;
    _T__12_t0b <= I_12_t0b;
    _T__12_t1b_t0b <= I_12_t1b_t0b;
    _T__12_t1b_t1b <= I_12_t1b_t1b;
    _T__13_t0b <= I_13_t0b;
    _T__13_t1b_t0b <= I_13_t1b_t0b;
    _T__13_t1b_t1b <= I_13_t1b_t1b;
    _T__14_t0b <= I_14_t0b;
    _T__14_t1b_t0b <= I_14_t1b_t0b;
    _T__14_t1b_t1b <= I_14_t1b_t1b;
    _T__15_t0b <= I_15_t0b;
    _T__15_t1b_t0b <= I_15_t1b_t0b;
    _T__15_t1b_t1b <= I_15_t1b_t1b;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module Top(
  input         clock,
  input         reset,
  input         valid_up,
  output        valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  input  [31:0] I_4,
  input  [31:0] I_5,
  input  [31:0] I_6,
  input  [31:0] I_7,
  input  [31:0] I_8,
  input  [31:0] I_9,
  input  [31:0] I_10,
  input  [31:0] I_11,
  input  [31:0] I_12,
  input  [31:0] I_13,
  input  [31:0] I_14,
  input  [31:0] I_15,
  output [31:0] O_0_t0b,
  output [31:0] O_0_t1b_t0b,
  output [31:0] O_0_t1b_t1b,
  output [31:0] O_1_t0b,
  output [31:0] O_1_t1b_t0b,
  output [31:0] O_1_t1b_t1b,
  output [31:0] O_2_t0b,
  output [31:0] O_2_t1b_t0b,
  output [31:0] O_2_t1b_t1b,
  output [31:0] O_3_t0b,
  output [31:0] O_3_t1b_t0b,
  output [31:0] O_3_t1b_t1b,
  output [31:0] O_4_t0b,
  output [31:0] O_4_t1b_t0b,
  output [31:0] O_4_t1b_t1b,
  output [31:0] O_5_t0b,
  output [31:0] O_5_t1b_t0b,
  output [31:0] O_5_t1b_t1b,
  output [31:0] O_6_t0b,
  output [31:0] O_6_t1b_t0b,
  output [31:0] O_6_t1b_t1b,
  output [31:0] O_7_t0b,
  output [31:0] O_7_t1b_t0b,
  output [31:0] O_7_t1b_t1b,
  output [31:0] O_8_t0b,
  output [31:0] O_8_t1b_t0b,
  output [31:0] O_8_t1b_t1b,
  output [31:0] O_9_t0b,
  output [31:0] O_9_t1b_t0b,
  output [31:0] O_9_t1b_t1b,
  output [31:0] O_10_t0b,
  output [31:0] O_10_t1b_t0b,
  output [31:0] O_10_t1b_t1b,
  output [31:0] O_11_t0b,
  output [31:0] O_11_t1b_t0b,
  output [31:0] O_11_t1b_t1b,
  output [31:0] O_12_t0b,
  output [31:0] O_12_t1b_t0b,
  output [31:0] O_12_t1b_t1b,
  output [31:0] O_13_t0b,
  output [31:0] O_13_t1b_t0b,
  output [31:0] O_13_t1b_t1b,
  output [31:0] O_14_t0b,
  output [31:0] O_14_t1b_t0b,
  output [31:0] O_14_t1b_t1b,
  output [31:0] O_15_t0b,
  output [31:0] O_15_t1b_t0b,
  output [31:0] O_15_t1b_t1b
);
  wire  n1_clock; // @[Top.scala 357:20]
  wire  n1_reset; // @[Top.scala 357:20]
  wire  n1_valid_up; // @[Top.scala 357:20]
  wire  n1_valid_down; // @[Top.scala 357:20]
  wire [31:0] n1_I_0; // @[Top.scala 357:20]
  wire [31:0] n1_I_1; // @[Top.scala 357:20]
  wire [31:0] n1_I_2; // @[Top.scala 357:20]
  wire [31:0] n1_I_3; // @[Top.scala 357:20]
  wire [31:0] n1_I_4; // @[Top.scala 357:20]
  wire [31:0] n1_I_5; // @[Top.scala 357:20]
  wire [31:0] n1_I_6; // @[Top.scala 357:20]
  wire [31:0] n1_I_7; // @[Top.scala 357:20]
  wire [31:0] n1_I_8; // @[Top.scala 357:20]
  wire [31:0] n1_I_9; // @[Top.scala 357:20]
  wire [31:0] n1_I_10; // @[Top.scala 357:20]
  wire [31:0] n1_I_11; // @[Top.scala 357:20]
  wire [31:0] n1_I_12; // @[Top.scala 357:20]
  wire [31:0] n1_I_13; // @[Top.scala 357:20]
  wire [31:0] n1_I_14; // @[Top.scala 357:20]
  wire [31:0] n1_I_15; // @[Top.scala 357:20]
  wire [31:0] n1_O_0; // @[Top.scala 357:20]
  wire [31:0] n1_O_1; // @[Top.scala 357:20]
  wire [31:0] n1_O_2; // @[Top.scala 357:20]
  wire [31:0] n1_O_3; // @[Top.scala 357:20]
  wire [31:0] n1_O_4; // @[Top.scala 357:20]
  wire [31:0] n1_O_5; // @[Top.scala 357:20]
  wire [31:0] n1_O_6; // @[Top.scala 357:20]
  wire [31:0] n1_O_7; // @[Top.scala 357:20]
  wire [31:0] n1_O_8; // @[Top.scala 357:20]
  wire [31:0] n1_O_9; // @[Top.scala 357:20]
  wire [31:0] n1_O_10; // @[Top.scala 357:20]
  wire [31:0] n1_O_11; // @[Top.scala 357:20]
  wire [31:0] n1_O_12; // @[Top.scala 357:20]
  wire [31:0] n1_O_13; // @[Top.scala 357:20]
  wire [31:0] n1_O_14; // @[Top.scala 357:20]
  wire [31:0] n1_O_15; // @[Top.scala 357:20]
  wire  n2_clock; // @[Top.scala 360:20]
  wire  n2_reset; // @[Top.scala 360:20]
  wire  n2_valid_up; // @[Top.scala 360:20]
  wire  n2_valid_down; // @[Top.scala 360:20]
  wire [31:0] n2_I_0; // @[Top.scala 360:20]
  wire [31:0] n2_I_1; // @[Top.scala 360:20]
  wire [31:0] n2_I_2; // @[Top.scala 360:20]
  wire [31:0] n2_I_3; // @[Top.scala 360:20]
  wire [31:0] n2_I_4; // @[Top.scala 360:20]
  wire [31:0] n2_I_5; // @[Top.scala 360:20]
  wire [31:0] n2_I_6; // @[Top.scala 360:20]
  wire [31:0] n2_I_7; // @[Top.scala 360:20]
  wire [31:0] n2_I_8; // @[Top.scala 360:20]
  wire [31:0] n2_I_9; // @[Top.scala 360:20]
  wire [31:0] n2_I_10; // @[Top.scala 360:20]
  wire [31:0] n2_I_11; // @[Top.scala 360:20]
  wire [31:0] n2_I_12; // @[Top.scala 360:20]
  wire [31:0] n2_I_13; // @[Top.scala 360:20]
  wire [31:0] n2_I_14; // @[Top.scala 360:20]
  wire [31:0] n2_I_15; // @[Top.scala 360:20]
  wire [31:0] n2_O_0; // @[Top.scala 360:20]
  wire [31:0] n2_O_1; // @[Top.scala 360:20]
  wire [31:0] n2_O_2; // @[Top.scala 360:20]
  wire [31:0] n2_O_3; // @[Top.scala 360:20]
  wire [31:0] n2_O_4; // @[Top.scala 360:20]
  wire [31:0] n2_O_5; // @[Top.scala 360:20]
  wire [31:0] n2_O_6; // @[Top.scala 360:20]
  wire [31:0] n2_O_7; // @[Top.scala 360:20]
  wire [31:0] n2_O_8; // @[Top.scala 360:20]
  wire [31:0] n2_O_9; // @[Top.scala 360:20]
  wire [31:0] n2_O_10; // @[Top.scala 360:20]
  wire [31:0] n2_O_11; // @[Top.scala 360:20]
  wire [31:0] n2_O_12; // @[Top.scala 360:20]
  wire [31:0] n2_O_13; // @[Top.scala 360:20]
  wire [31:0] n2_O_14; // @[Top.scala 360:20]
  wire [31:0] n2_O_15; // @[Top.scala 360:20]
  wire  n3_clock; // @[Top.scala 363:20]
  wire  n3_reset; // @[Top.scala 363:20]
  wire  n3_valid_up; // @[Top.scala 363:20]
  wire  n3_valid_down; // @[Top.scala 363:20]
  wire [31:0] n3_I_0; // @[Top.scala 363:20]
  wire [31:0] n3_I_1; // @[Top.scala 363:20]
  wire [31:0] n3_I_2; // @[Top.scala 363:20]
  wire [31:0] n3_I_3; // @[Top.scala 363:20]
  wire [31:0] n3_I_4; // @[Top.scala 363:20]
  wire [31:0] n3_I_5; // @[Top.scala 363:20]
  wire [31:0] n3_I_6; // @[Top.scala 363:20]
  wire [31:0] n3_I_7; // @[Top.scala 363:20]
  wire [31:0] n3_I_8; // @[Top.scala 363:20]
  wire [31:0] n3_I_9; // @[Top.scala 363:20]
  wire [31:0] n3_I_10; // @[Top.scala 363:20]
  wire [31:0] n3_I_11; // @[Top.scala 363:20]
  wire [31:0] n3_I_12; // @[Top.scala 363:20]
  wire [31:0] n3_I_13; // @[Top.scala 363:20]
  wire [31:0] n3_I_14; // @[Top.scala 363:20]
  wire [31:0] n3_I_15; // @[Top.scala 363:20]
  wire [31:0] n3_O_0; // @[Top.scala 363:20]
  wire [31:0] n3_O_1; // @[Top.scala 363:20]
  wire [31:0] n3_O_2; // @[Top.scala 363:20]
  wire [31:0] n3_O_3; // @[Top.scala 363:20]
  wire [31:0] n3_O_4; // @[Top.scala 363:20]
  wire [31:0] n3_O_5; // @[Top.scala 363:20]
  wire [31:0] n3_O_6; // @[Top.scala 363:20]
  wire [31:0] n3_O_7; // @[Top.scala 363:20]
  wire [31:0] n3_O_8; // @[Top.scala 363:20]
  wire [31:0] n3_O_9; // @[Top.scala 363:20]
  wire [31:0] n3_O_10; // @[Top.scala 363:20]
  wire [31:0] n3_O_11; // @[Top.scala 363:20]
  wire [31:0] n3_O_12; // @[Top.scala 363:20]
  wire [31:0] n3_O_13; // @[Top.scala 363:20]
  wire [31:0] n3_O_14; // @[Top.scala 363:20]
  wire [31:0] n3_O_15; // @[Top.scala 363:20]
  wire  n4_clock; // @[Top.scala 366:20]
  wire  n4_valid_up; // @[Top.scala 366:20]
  wire  n4_valid_down; // @[Top.scala 366:20]
  wire [31:0] n4_I_0; // @[Top.scala 366:20]
  wire [31:0] n4_I_1; // @[Top.scala 366:20]
  wire [31:0] n4_I_2; // @[Top.scala 366:20]
  wire [31:0] n4_I_3; // @[Top.scala 366:20]
  wire [31:0] n4_I_4; // @[Top.scala 366:20]
  wire [31:0] n4_I_5; // @[Top.scala 366:20]
  wire [31:0] n4_I_6; // @[Top.scala 366:20]
  wire [31:0] n4_I_7; // @[Top.scala 366:20]
  wire [31:0] n4_I_8; // @[Top.scala 366:20]
  wire [31:0] n4_I_9; // @[Top.scala 366:20]
  wire [31:0] n4_I_10; // @[Top.scala 366:20]
  wire [31:0] n4_I_11; // @[Top.scala 366:20]
  wire [31:0] n4_I_12; // @[Top.scala 366:20]
  wire [31:0] n4_I_13; // @[Top.scala 366:20]
  wire [31:0] n4_I_14; // @[Top.scala 366:20]
  wire [31:0] n4_I_15; // @[Top.scala 366:20]
  wire [31:0] n4_O_0; // @[Top.scala 366:20]
  wire [31:0] n4_O_1; // @[Top.scala 366:20]
  wire [31:0] n4_O_2; // @[Top.scala 366:20]
  wire [31:0] n4_O_3; // @[Top.scala 366:20]
  wire [31:0] n4_O_4; // @[Top.scala 366:20]
  wire [31:0] n4_O_5; // @[Top.scala 366:20]
  wire [31:0] n4_O_6; // @[Top.scala 366:20]
  wire [31:0] n4_O_7; // @[Top.scala 366:20]
  wire [31:0] n4_O_8; // @[Top.scala 366:20]
  wire [31:0] n4_O_9; // @[Top.scala 366:20]
  wire [31:0] n4_O_10; // @[Top.scala 366:20]
  wire [31:0] n4_O_11; // @[Top.scala 366:20]
  wire [31:0] n4_O_12; // @[Top.scala 366:20]
  wire [31:0] n4_O_13; // @[Top.scala 366:20]
  wire [31:0] n4_O_14; // @[Top.scala 366:20]
  wire [31:0] n4_O_15; // @[Top.scala 366:20]
  wire  n5_clock; // @[Top.scala 369:20]
  wire  n5_valid_up; // @[Top.scala 369:20]
  wire  n5_valid_down; // @[Top.scala 369:20]
  wire [31:0] n5_I_0; // @[Top.scala 369:20]
  wire [31:0] n5_I_1; // @[Top.scala 369:20]
  wire [31:0] n5_I_2; // @[Top.scala 369:20]
  wire [31:0] n5_I_3; // @[Top.scala 369:20]
  wire [31:0] n5_I_4; // @[Top.scala 369:20]
  wire [31:0] n5_I_5; // @[Top.scala 369:20]
  wire [31:0] n5_I_6; // @[Top.scala 369:20]
  wire [31:0] n5_I_7; // @[Top.scala 369:20]
  wire [31:0] n5_I_8; // @[Top.scala 369:20]
  wire [31:0] n5_I_9; // @[Top.scala 369:20]
  wire [31:0] n5_I_10; // @[Top.scala 369:20]
  wire [31:0] n5_I_11; // @[Top.scala 369:20]
  wire [31:0] n5_I_12; // @[Top.scala 369:20]
  wire [31:0] n5_I_13; // @[Top.scala 369:20]
  wire [31:0] n5_I_14; // @[Top.scala 369:20]
  wire [31:0] n5_I_15; // @[Top.scala 369:20]
  wire [31:0] n5_O_0; // @[Top.scala 369:20]
  wire [31:0] n5_O_1; // @[Top.scala 369:20]
  wire [31:0] n5_O_2; // @[Top.scala 369:20]
  wire [31:0] n5_O_3; // @[Top.scala 369:20]
  wire [31:0] n5_O_4; // @[Top.scala 369:20]
  wire [31:0] n5_O_5; // @[Top.scala 369:20]
  wire [31:0] n5_O_6; // @[Top.scala 369:20]
  wire [31:0] n5_O_7; // @[Top.scala 369:20]
  wire [31:0] n5_O_8; // @[Top.scala 369:20]
  wire [31:0] n5_O_9; // @[Top.scala 369:20]
  wire [31:0] n5_O_10; // @[Top.scala 369:20]
  wire [31:0] n5_O_11; // @[Top.scala 369:20]
  wire [31:0] n5_O_12; // @[Top.scala 369:20]
  wire [31:0] n5_O_13; // @[Top.scala 369:20]
  wire [31:0] n5_O_14; // @[Top.scala 369:20]
  wire [31:0] n5_O_15; // @[Top.scala 369:20]
  wire  n6_valid_up; // @[Top.scala 372:20]
  wire  n6_valid_down; // @[Top.scala 372:20]
  wire [31:0] n6_I0_0; // @[Top.scala 372:20]
  wire [31:0] n6_I0_1; // @[Top.scala 372:20]
  wire [31:0] n6_I0_2; // @[Top.scala 372:20]
  wire [31:0] n6_I0_3; // @[Top.scala 372:20]
  wire [31:0] n6_I0_4; // @[Top.scala 372:20]
  wire [31:0] n6_I0_5; // @[Top.scala 372:20]
  wire [31:0] n6_I0_6; // @[Top.scala 372:20]
  wire [31:0] n6_I0_7; // @[Top.scala 372:20]
  wire [31:0] n6_I0_8; // @[Top.scala 372:20]
  wire [31:0] n6_I0_9; // @[Top.scala 372:20]
  wire [31:0] n6_I0_10; // @[Top.scala 372:20]
  wire [31:0] n6_I0_11; // @[Top.scala 372:20]
  wire [31:0] n6_I0_12; // @[Top.scala 372:20]
  wire [31:0] n6_I0_13; // @[Top.scala 372:20]
  wire [31:0] n6_I0_14; // @[Top.scala 372:20]
  wire [31:0] n6_I0_15; // @[Top.scala 372:20]
  wire [31:0] n6_I1_0; // @[Top.scala 372:20]
  wire [31:0] n6_I1_1; // @[Top.scala 372:20]
  wire [31:0] n6_I1_2; // @[Top.scala 372:20]
  wire [31:0] n6_I1_3; // @[Top.scala 372:20]
  wire [31:0] n6_I1_4; // @[Top.scala 372:20]
  wire [31:0] n6_I1_5; // @[Top.scala 372:20]
  wire [31:0] n6_I1_6; // @[Top.scala 372:20]
  wire [31:0] n6_I1_7; // @[Top.scala 372:20]
  wire [31:0] n6_I1_8; // @[Top.scala 372:20]
  wire [31:0] n6_I1_9; // @[Top.scala 372:20]
  wire [31:0] n6_I1_10; // @[Top.scala 372:20]
  wire [31:0] n6_I1_11; // @[Top.scala 372:20]
  wire [31:0] n6_I1_12; // @[Top.scala 372:20]
  wire [31:0] n6_I1_13; // @[Top.scala 372:20]
  wire [31:0] n6_I1_14; // @[Top.scala 372:20]
  wire [31:0] n6_I1_15; // @[Top.scala 372:20]
  wire [31:0] n6_O_0_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_0_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_1_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_1_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_2_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_2_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_3_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_3_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_4_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_4_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_5_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_5_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_6_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_6_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_7_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_7_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_8_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_8_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_9_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_9_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_10_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_10_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_11_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_11_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_12_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_12_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_13_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_13_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_14_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_14_1; // @[Top.scala 372:20]
  wire [31:0] n6_O_15_0; // @[Top.scala 372:20]
  wire [31:0] n6_O_15_1; // @[Top.scala 372:20]
  wire  n13_valid_up; // @[Top.scala 376:21]
  wire  n13_valid_down; // @[Top.scala 376:21]
  wire [31:0] n13_I0_0_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_0_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_1_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_1_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_2_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_2_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_3_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_3_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_4_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_4_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_5_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_5_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_6_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_6_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_7_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_7_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_8_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_8_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_9_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_9_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_10_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_10_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_11_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_11_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_12_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_12_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_13_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_13_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_14_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_14_1; // @[Top.scala 376:21]
  wire [31:0] n13_I0_15_0; // @[Top.scala 376:21]
  wire [31:0] n13_I0_15_1; // @[Top.scala 376:21]
  wire [31:0] n13_I1_0; // @[Top.scala 376:21]
  wire [31:0] n13_I1_1; // @[Top.scala 376:21]
  wire [31:0] n13_I1_2; // @[Top.scala 376:21]
  wire [31:0] n13_I1_3; // @[Top.scala 376:21]
  wire [31:0] n13_I1_4; // @[Top.scala 376:21]
  wire [31:0] n13_I1_5; // @[Top.scala 376:21]
  wire [31:0] n13_I1_6; // @[Top.scala 376:21]
  wire [31:0] n13_I1_7; // @[Top.scala 376:21]
  wire [31:0] n13_I1_8; // @[Top.scala 376:21]
  wire [31:0] n13_I1_9; // @[Top.scala 376:21]
  wire [31:0] n13_I1_10; // @[Top.scala 376:21]
  wire [31:0] n13_I1_11; // @[Top.scala 376:21]
  wire [31:0] n13_I1_12; // @[Top.scala 376:21]
  wire [31:0] n13_I1_13; // @[Top.scala 376:21]
  wire [31:0] n13_I1_14; // @[Top.scala 376:21]
  wire [31:0] n13_I1_15; // @[Top.scala 376:21]
  wire [31:0] n13_O_0_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_0_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_0_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_1_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_1_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_1_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_2_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_2_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_2_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_3_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_3_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_3_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_4_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_4_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_4_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_5_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_5_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_5_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_6_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_6_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_6_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_7_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_7_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_7_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_8_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_8_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_8_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_9_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_9_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_9_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_10_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_10_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_10_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_11_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_11_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_11_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_12_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_12_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_12_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_13_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_13_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_13_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_14_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_14_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_14_2; // @[Top.scala 376:21]
  wire [31:0] n13_O_15_0; // @[Top.scala 376:21]
  wire [31:0] n13_O_15_1; // @[Top.scala 376:21]
  wire [31:0] n13_O_15_2; // @[Top.scala 376:21]
  wire  n22_valid_up; // @[Top.scala 380:21]
  wire  n22_valid_down; // @[Top.scala 380:21]
  wire [31:0] n22_I_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_1_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_1_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_1_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_2_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_2_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_2_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_3_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_3_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_3_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_4_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_4_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_4_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_5_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_5_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_5_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_6_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_6_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_6_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_7_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_7_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_7_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_8_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_8_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_8_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_9_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_9_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_9_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_10_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_10_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_10_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_11_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_11_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_11_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_12_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_12_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_12_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_13_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_13_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_13_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_14_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_14_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_14_2; // @[Top.scala 380:21]
  wire [31:0] n22_I_15_0; // @[Top.scala 380:21]
  wire [31:0] n22_I_15_1; // @[Top.scala 380:21]
  wire [31:0] n22_I_15_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_0_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_0_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_0_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_1_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_1_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_1_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_2_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_2_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_2_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_3_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_3_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_3_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_4_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_4_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_4_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_5_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_5_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_5_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_6_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_6_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_6_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_7_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_7_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_7_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_8_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_8_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_8_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_9_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_9_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_9_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_10_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_10_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_10_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_11_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_11_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_11_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_12_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_12_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_12_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_13_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_13_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_13_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_14_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_14_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_14_0_2; // @[Top.scala 380:21]
  wire [31:0] n22_O_15_0_0; // @[Top.scala 380:21]
  wire [31:0] n22_O_15_0_1; // @[Top.scala 380:21]
  wire [31:0] n22_O_15_0_2; // @[Top.scala 380:21]
  wire  n29_valid_up; // @[Top.scala 383:21]
  wire  n29_valid_down; // @[Top.scala 383:21]
  wire [31:0] n29_I_0_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_0_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_0_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_1_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_1_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_1_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_2_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_2_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_2_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_3_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_3_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_3_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_4_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_4_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_4_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_5_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_5_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_5_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_6_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_6_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_6_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_7_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_7_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_7_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_8_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_8_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_8_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_9_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_9_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_9_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_10_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_10_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_10_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_11_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_11_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_11_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_12_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_12_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_12_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_13_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_13_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_13_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_14_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_14_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_14_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_I_15_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_I_15_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_I_15_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_0_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_0_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_0_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_1_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_1_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_1_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_2_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_2_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_2_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_3_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_3_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_3_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_4_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_4_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_4_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_5_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_5_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_5_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_6_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_6_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_6_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_7_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_7_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_7_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_8_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_8_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_8_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_9_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_9_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_9_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_10_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_10_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_10_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_11_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_11_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_11_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_12_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_12_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_12_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_13_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_13_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_13_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_14_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_14_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_14_2; // @[Top.scala 383:21]
  wire [31:0] n29_O_15_0; // @[Top.scala 383:21]
  wire [31:0] n29_O_15_1; // @[Top.scala 383:21]
  wire [31:0] n29_O_15_2; // @[Top.scala 383:21]
  wire  n30_clock; // @[Top.scala 386:21]
  wire  n30_valid_up; // @[Top.scala 386:21]
  wire  n30_valid_down; // @[Top.scala 386:21]
  wire [31:0] n30_I_0; // @[Top.scala 386:21]
  wire [31:0] n30_I_1; // @[Top.scala 386:21]
  wire [31:0] n30_I_2; // @[Top.scala 386:21]
  wire [31:0] n30_I_3; // @[Top.scala 386:21]
  wire [31:0] n30_I_4; // @[Top.scala 386:21]
  wire [31:0] n30_I_5; // @[Top.scala 386:21]
  wire [31:0] n30_I_6; // @[Top.scala 386:21]
  wire [31:0] n30_I_7; // @[Top.scala 386:21]
  wire [31:0] n30_I_8; // @[Top.scala 386:21]
  wire [31:0] n30_I_9; // @[Top.scala 386:21]
  wire [31:0] n30_I_10; // @[Top.scala 386:21]
  wire [31:0] n30_I_11; // @[Top.scala 386:21]
  wire [31:0] n30_I_12; // @[Top.scala 386:21]
  wire [31:0] n30_I_13; // @[Top.scala 386:21]
  wire [31:0] n30_I_14; // @[Top.scala 386:21]
  wire [31:0] n30_I_15; // @[Top.scala 386:21]
  wire [31:0] n30_O_0; // @[Top.scala 386:21]
  wire [31:0] n30_O_1; // @[Top.scala 386:21]
  wire [31:0] n30_O_2; // @[Top.scala 386:21]
  wire [31:0] n30_O_3; // @[Top.scala 386:21]
  wire [31:0] n30_O_4; // @[Top.scala 386:21]
  wire [31:0] n30_O_5; // @[Top.scala 386:21]
  wire [31:0] n30_O_6; // @[Top.scala 386:21]
  wire [31:0] n30_O_7; // @[Top.scala 386:21]
  wire [31:0] n30_O_8; // @[Top.scala 386:21]
  wire [31:0] n30_O_9; // @[Top.scala 386:21]
  wire [31:0] n30_O_10; // @[Top.scala 386:21]
  wire [31:0] n30_O_11; // @[Top.scala 386:21]
  wire [31:0] n30_O_12; // @[Top.scala 386:21]
  wire [31:0] n30_O_13; // @[Top.scala 386:21]
  wire [31:0] n30_O_14; // @[Top.scala 386:21]
  wire [31:0] n30_O_15; // @[Top.scala 386:21]
  wire  n31_clock; // @[Top.scala 389:21]
  wire  n31_valid_up; // @[Top.scala 389:21]
  wire  n31_valid_down; // @[Top.scala 389:21]
  wire [31:0] n31_I_0; // @[Top.scala 389:21]
  wire [31:0] n31_I_1; // @[Top.scala 389:21]
  wire [31:0] n31_I_2; // @[Top.scala 389:21]
  wire [31:0] n31_I_3; // @[Top.scala 389:21]
  wire [31:0] n31_I_4; // @[Top.scala 389:21]
  wire [31:0] n31_I_5; // @[Top.scala 389:21]
  wire [31:0] n31_I_6; // @[Top.scala 389:21]
  wire [31:0] n31_I_7; // @[Top.scala 389:21]
  wire [31:0] n31_I_8; // @[Top.scala 389:21]
  wire [31:0] n31_I_9; // @[Top.scala 389:21]
  wire [31:0] n31_I_10; // @[Top.scala 389:21]
  wire [31:0] n31_I_11; // @[Top.scala 389:21]
  wire [31:0] n31_I_12; // @[Top.scala 389:21]
  wire [31:0] n31_I_13; // @[Top.scala 389:21]
  wire [31:0] n31_I_14; // @[Top.scala 389:21]
  wire [31:0] n31_I_15; // @[Top.scala 389:21]
  wire [31:0] n31_O_0; // @[Top.scala 389:21]
  wire [31:0] n31_O_1; // @[Top.scala 389:21]
  wire [31:0] n31_O_2; // @[Top.scala 389:21]
  wire [31:0] n31_O_3; // @[Top.scala 389:21]
  wire [31:0] n31_O_4; // @[Top.scala 389:21]
  wire [31:0] n31_O_5; // @[Top.scala 389:21]
  wire [31:0] n31_O_6; // @[Top.scala 389:21]
  wire [31:0] n31_O_7; // @[Top.scala 389:21]
  wire [31:0] n31_O_8; // @[Top.scala 389:21]
  wire [31:0] n31_O_9; // @[Top.scala 389:21]
  wire [31:0] n31_O_10; // @[Top.scala 389:21]
  wire [31:0] n31_O_11; // @[Top.scala 389:21]
  wire [31:0] n31_O_12; // @[Top.scala 389:21]
  wire [31:0] n31_O_13; // @[Top.scala 389:21]
  wire [31:0] n31_O_14; // @[Top.scala 389:21]
  wire [31:0] n31_O_15; // @[Top.scala 389:21]
  wire  n32_valid_up; // @[Top.scala 392:21]
  wire  n32_valid_down; // @[Top.scala 392:21]
  wire [31:0] n32_I0_0; // @[Top.scala 392:21]
  wire [31:0] n32_I0_1; // @[Top.scala 392:21]
  wire [31:0] n32_I0_2; // @[Top.scala 392:21]
  wire [31:0] n32_I0_3; // @[Top.scala 392:21]
  wire [31:0] n32_I0_4; // @[Top.scala 392:21]
  wire [31:0] n32_I0_5; // @[Top.scala 392:21]
  wire [31:0] n32_I0_6; // @[Top.scala 392:21]
  wire [31:0] n32_I0_7; // @[Top.scala 392:21]
  wire [31:0] n32_I0_8; // @[Top.scala 392:21]
  wire [31:0] n32_I0_9; // @[Top.scala 392:21]
  wire [31:0] n32_I0_10; // @[Top.scala 392:21]
  wire [31:0] n32_I0_11; // @[Top.scala 392:21]
  wire [31:0] n32_I0_12; // @[Top.scala 392:21]
  wire [31:0] n32_I0_13; // @[Top.scala 392:21]
  wire [31:0] n32_I0_14; // @[Top.scala 392:21]
  wire [31:0] n32_I0_15; // @[Top.scala 392:21]
  wire [31:0] n32_I1_0; // @[Top.scala 392:21]
  wire [31:0] n32_I1_1; // @[Top.scala 392:21]
  wire [31:0] n32_I1_2; // @[Top.scala 392:21]
  wire [31:0] n32_I1_3; // @[Top.scala 392:21]
  wire [31:0] n32_I1_4; // @[Top.scala 392:21]
  wire [31:0] n32_I1_5; // @[Top.scala 392:21]
  wire [31:0] n32_I1_6; // @[Top.scala 392:21]
  wire [31:0] n32_I1_7; // @[Top.scala 392:21]
  wire [31:0] n32_I1_8; // @[Top.scala 392:21]
  wire [31:0] n32_I1_9; // @[Top.scala 392:21]
  wire [31:0] n32_I1_10; // @[Top.scala 392:21]
  wire [31:0] n32_I1_11; // @[Top.scala 392:21]
  wire [31:0] n32_I1_12; // @[Top.scala 392:21]
  wire [31:0] n32_I1_13; // @[Top.scala 392:21]
  wire [31:0] n32_I1_14; // @[Top.scala 392:21]
  wire [31:0] n32_I1_15; // @[Top.scala 392:21]
  wire [31:0] n32_O_0_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_0_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_1_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_1_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_2_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_2_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_3_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_3_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_4_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_4_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_5_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_5_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_6_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_6_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_7_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_7_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_8_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_8_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_9_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_9_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_10_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_10_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_11_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_11_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_12_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_12_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_13_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_13_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_14_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_14_1; // @[Top.scala 392:21]
  wire [31:0] n32_O_15_0; // @[Top.scala 392:21]
  wire [31:0] n32_O_15_1; // @[Top.scala 392:21]
  wire  n39_valid_up; // @[Top.scala 396:21]
  wire  n39_valid_down; // @[Top.scala 396:21]
  wire [31:0] n39_I0_0_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_0_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_1_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_1_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_2_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_2_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_3_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_3_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_4_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_4_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_5_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_5_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_6_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_6_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_7_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_7_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_8_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_8_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_9_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_9_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_10_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_10_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_11_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_11_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_12_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_12_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_13_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_13_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_14_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_14_1; // @[Top.scala 396:21]
  wire [31:0] n39_I0_15_0; // @[Top.scala 396:21]
  wire [31:0] n39_I0_15_1; // @[Top.scala 396:21]
  wire [31:0] n39_I1_0; // @[Top.scala 396:21]
  wire [31:0] n39_I1_1; // @[Top.scala 396:21]
  wire [31:0] n39_I1_2; // @[Top.scala 396:21]
  wire [31:0] n39_I1_3; // @[Top.scala 396:21]
  wire [31:0] n39_I1_4; // @[Top.scala 396:21]
  wire [31:0] n39_I1_5; // @[Top.scala 396:21]
  wire [31:0] n39_I1_6; // @[Top.scala 396:21]
  wire [31:0] n39_I1_7; // @[Top.scala 396:21]
  wire [31:0] n39_I1_8; // @[Top.scala 396:21]
  wire [31:0] n39_I1_9; // @[Top.scala 396:21]
  wire [31:0] n39_I1_10; // @[Top.scala 396:21]
  wire [31:0] n39_I1_11; // @[Top.scala 396:21]
  wire [31:0] n39_I1_12; // @[Top.scala 396:21]
  wire [31:0] n39_I1_13; // @[Top.scala 396:21]
  wire [31:0] n39_I1_14; // @[Top.scala 396:21]
  wire [31:0] n39_I1_15; // @[Top.scala 396:21]
  wire [31:0] n39_O_0_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_0_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_0_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_1_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_1_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_1_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_2_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_2_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_2_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_3_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_3_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_3_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_4_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_4_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_4_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_5_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_5_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_5_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_6_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_6_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_6_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_7_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_7_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_7_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_8_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_8_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_8_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_9_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_9_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_9_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_10_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_10_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_10_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_11_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_11_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_11_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_12_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_12_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_12_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_13_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_13_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_13_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_14_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_14_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_14_2; // @[Top.scala 396:21]
  wire [31:0] n39_O_15_0; // @[Top.scala 396:21]
  wire [31:0] n39_O_15_1; // @[Top.scala 396:21]
  wire [31:0] n39_O_15_2; // @[Top.scala 396:21]
  wire  n48_valid_up; // @[Top.scala 400:21]
  wire  n48_valid_down; // @[Top.scala 400:21]
  wire [31:0] n48_I_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_1_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_1_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_1_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_2_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_2_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_2_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_3_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_3_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_3_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_4_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_4_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_4_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_5_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_5_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_5_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_6_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_6_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_6_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_7_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_7_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_7_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_8_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_8_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_8_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_9_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_9_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_9_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_10_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_10_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_10_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_11_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_11_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_11_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_12_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_12_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_12_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_13_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_13_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_13_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_14_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_14_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_14_2; // @[Top.scala 400:21]
  wire [31:0] n48_I_15_0; // @[Top.scala 400:21]
  wire [31:0] n48_I_15_1; // @[Top.scala 400:21]
  wire [31:0] n48_I_15_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_0_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_0_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_0_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_1_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_1_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_1_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_2_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_2_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_2_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_3_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_3_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_3_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_4_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_4_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_4_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_5_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_5_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_5_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_6_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_6_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_6_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_7_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_7_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_7_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_8_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_8_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_8_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_9_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_9_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_9_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_10_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_10_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_10_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_11_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_11_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_11_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_12_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_12_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_12_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_13_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_13_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_13_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_14_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_14_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_14_0_2; // @[Top.scala 400:21]
  wire [31:0] n48_O_15_0_0; // @[Top.scala 400:21]
  wire [31:0] n48_O_15_0_1; // @[Top.scala 400:21]
  wire [31:0] n48_O_15_0_2; // @[Top.scala 400:21]
  wire  n55_valid_up; // @[Top.scala 403:21]
  wire  n55_valid_down; // @[Top.scala 403:21]
  wire [31:0] n55_I_0_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_0_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_0_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_1_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_1_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_1_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_2_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_2_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_2_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_3_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_3_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_3_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_4_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_4_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_4_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_5_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_5_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_5_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_6_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_6_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_6_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_7_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_7_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_7_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_8_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_8_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_8_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_9_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_9_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_9_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_10_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_10_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_10_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_11_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_11_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_11_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_12_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_12_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_12_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_13_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_13_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_13_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_14_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_14_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_14_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_I_15_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_I_15_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_I_15_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_0_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_0_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_0_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_1_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_1_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_1_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_2_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_2_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_2_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_3_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_3_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_3_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_4_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_4_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_4_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_5_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_5_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_5_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_6_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_6_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_6_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_7_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_7_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_7_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_8_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_8_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_8_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_9_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_9_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_9_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_10_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_10_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_10_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_11_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_11_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_11_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_12_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_12_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_12_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_13_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_13_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_13_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_14_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_14_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_14_2; // @[Top.scala 403:21]
  wire [31:0] n55_O_15_0; // @[Top.scala 403:21]
  wire [31:0] n55_O_15_1; // @[Top.scala 403:21]
  wire [31:0] n55_O_15_2; // @[Top.scala 403:21]
  wire  n56_valid_up; // @[Top.scala 406:21]
  wire  n56_valid_down; // @[Top.scala 406:21]
  wire [31:0] n56_I0_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_2_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_2_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_2_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_3_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_3_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_3_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_4_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_4_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_4_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_5_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_5_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_5_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_6_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_6_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_6_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_7_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_7_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_7_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_8_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_8_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_8_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_9_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_9_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_9_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_10_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_10_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_10_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_11_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_11_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_11_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_12_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_12_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_12_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_13_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_13_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_13_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_14_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_14_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_14_2; // @[Top.scala 406:21]
  wire [31:0] n56_I0_15_0; // @[Top.scala 406:21]
  wire [31:0] n56_I0_15_1; // @[Top.scala 406:21]
  wire [31:0] n56_I0_15_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_2_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_2_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_2_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_3_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_3_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_3_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_4_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_4_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_4_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_5_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_5_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_5_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_6_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_6_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_6_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_7_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_7_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_7_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_8_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_8_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_8_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_9_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_9_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_9_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_10_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_10_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_10_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_11_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_11_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_11_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_12_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_12_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_12_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_13_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_13_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_13_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_14_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_14_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_14_2; // @[Top.scala 406:21]
  wire [31:0] n56_I1_15_0; // @[Top.scala 406:21]
  wire [31:0] n56_I1_15_1; // @[Top.scala 406:21]
  wire [31:0] n56_I1_15_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_0_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_0_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_0_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_0_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_0_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_0_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_1_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_1_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_1_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_1_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_1_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_1_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_2_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_2_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_2_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_2_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_2_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_2_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_3_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_3_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_3_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_3_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_3_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_3_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_4_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_4_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_4_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_4_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_4_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_4_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_5_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_5_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_5_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_5_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_5_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_5_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_6_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_6_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_6_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_6_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_6_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_6_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_7_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_7_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_7_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_7_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_7_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_7_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_8_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_8_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_8_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_8_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_8_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_8_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_9_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_9_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_9_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_9_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_9_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_9_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_10_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_10_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_10_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_10_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_10_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_10_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_11_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_11_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_11_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_11_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_11_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_11_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_12_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_12_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_12_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_12_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_12_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_12_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_13_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_13_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_13_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_13_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_13_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_13_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_14_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_14_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_14_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_14_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_14_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_14_1_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_15_0_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_15_0_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_15_0_2; // @[Top.scala 406:21]
  wire [31:0] n56_O_15_1_0; // @[Top.scala 406:21]
  wire [31:0] n56_O_15_1_1; // @[Top.scala 406:21]
  wire [31:0] n56_O_15_1_2; // @[Top.scala 406:21]
  wire  n63_clock; // @[Top.scala 410:21]
  wire  n63_valid_up; // @[Top.scala 410:21]
  wire  n63_valid_down; // @[Top.scala 410:21]
  wire [31:0] n63_I_0; // @[Top.scala 410:21]
  wire [31:0] n63_I_1; // @[Top.scala 410:21]
  wire [31:0] n63_I_2; // @[Top.scala 410:21]
  wire [31:0] n63_I_3; // @[Top.scala 410:21]
  wire [31:0] n63_I_4; // @[Top.scala 410:21]
  wire [31:0] n63_I_5; // @[Top.scala 410:21]
  wire [31:0] n63_I_6; // @[Top.scala 410:21]
  wire [31:0] n63_I_7; // @[Top.scala 410:21]
  wire [31:0] n63_I_8; // @[Top.scala 410:21]
  wire [31:0] n63_I_9; // @[Top.scala 410:21]
  wire [31:0] n63_I_10; // @[Top.scala 410:21]
  wire [31:0] n63_I_11; // @[Top.scala 410:21]
  wire [31:0] n63_I_12; // @[Top.scala 410:21]
  wire [31:0] n63_I_13; // @[Top.scala 410:21]
  wire [31:0] n63_I_14; // @[Top.scala 410:21]
  wire [31:0] n63_I_15; // @[Top.scala 410:21]
  wire [31:0] n63_O_0; // @[Top.scala 410:21]
  wire [31:0] n63_O_1; // @[Top.scala 410:21]
  wire [31:0] n63_O_2; // @[Top.scala 410:21]
  wire [31:0] n63_O_3; // @[Top.scala 410:21]
  wire [31:0] n63_O_4; // @[Top.scala 410:21]
  wire [31:0] n63_O_5; // @[Top.scala 410:21]
  wire [31:0] n63_O_6; // @[Top.scala 410:21]
  wire [31:0] n63_O_7; // @[Top.scala 410:21]
  wire [31:0] n63_O_8; // @[Top.scala 410:21]
  wire [31:0] n63_O_9; // @[Top.scala 410:21]
  wire [31:0] n63_O_10; // @[Top.scala 410:21]
  wire [31:0] n63_O_11; // @[Top.scala 410:21]
  wire [31:0] n63_O_12; // @[Top.scala 410:21]
  wire [31:0] n63_O_13; // @[Top.scala 410:21]
  wire [31:0] n63_O_14; // @[Top.scala 410:21]
  wire [31:0] n63_O_15; // @[Top.scala 410:21]
  wire  n64_clock; // @[Top.scala 413:21]
  wire  n64_valid_up; // @[Top.scala 413:21]
  wire  n64_valid_down; // @[Top.scala 413:21]
  wire [31:0] n64_I_0; // @[Top.scala 413:21]
  wire [31:0] n64_I_1; // @[Top.scala 413:21]
  wire [31:0] n64_I_2; // @[Top.scala 413:21]
  wire [31:0] n64_I_3; // @[Top.scala 413:21]
  wire [31:0] n64_I_4; // @[Top.scala 413:21]
  wire [31:0] n64_I_5; // @[Top.scala 413:21]
  wire [31:0] n64_I_6; // @[Top.scala 413:21]
  wire [31:0] n64_I_7; // @[Top.scala 413:21]
  wire [31:0] n64_I_8; // @[Top.scala 413:21]
  wire [31:0] n64_I_9; // @[Top.scala 413:21]
  wire [31:0] n64_I_10; // @[Top.scala 413:21]
  wire [31:0] n64_I_11; // @[Top.scala 413:21]
  wire [31:0] n64_I_12; // @[Top.scala 413:21]
  wire [31:0] n64_I_13; // @[Top.scala 413:21]
  wire [31:0] n64_I_14; // @[Top.scala 413:21]
  wire [31:0] n64_I_15; // @[Top.scala 413:21]
  wire [31:0] n64_O_0; // @[Top.scala 413:21]
  wire [31:0] n64_O_1; // @[Top.scala 413:21]
  wire [31:0] n64_O_2; // @[Top.scala 413:21]
  wire [31:0] n64_O_3; // @[Top.scala 413:21]
  wire [31:0] n64_O_4; // @[Top.scala 413:21]
  wire [31:0] n64_O_5; // @[Top.scala 413:21]
  wire [31:0] n64_O_6; // @[Top.scala 413:21]
  wire [31:0] n64_O_7; // @[Top.scala 413:21]
  wire [31:0] n64_O_8; // @[Top.scala 413:21]
  wire [31:0] n64_O_9; // @[Top.scala 413:21]
  wire [31:0] n64_O_10; // @[Top.scala 413:21]
  wire [31:0] n64_O_11; // @[Top.scala 413:21]
  wire [31:0] n64_O_12; // @[Top.scala 413:21]
  wire [31:0] n64_O_13; // @[Top.scala 413:21]
  wire [31:0] n64_O_14; // @[Top.scala 413:21]
  wire [31:0] n64_O_15; // @[Top.scala 413:21]
  wire  n65_valid_up; // @[Top.scala 416:21]
  wire  n65_valid_down; // @[Top.scala 416:21]
  wire [31:0] n65_I0_0; // @[Top.scala 416:21]
  wire [31:0] n65_I0_1; // @[Top.scala 416:21]
  wire [31:0] n65_I0_2; // @[Top.scala 416:21]
  wire [31:0] n65_I0_3; // @[Top.scala 416:21]
  wire [31:0] n65_I0_4; // @[Top.scala 416:21]
  wire [31:0] n65_I0_5; // @[Top.scala 416:21]
  wire [31:0] n65_I0_6; // @[Top.scala 416:21]
  wire [31:0] n65_I0_7; // @[Top.scala 416:21]
  wire [31:0] n65_I0_8; // @[Top.scala 416:21]
  wire [31:0] n65_I0_9; // @[Top.scala 416:21]
  wire [31:0] n65_I0_10; // @[Top.scala 416:21]
  wire [31:0] n65_I0_11; // @[Top.scala 416:21]
  wire [31:0] n65_I0_12; // @[Top.scala 416:21]
  wire [31:0] n65_I0_13; // @[Top.scala 416:21]
  wire [31:0] n65_I0_14; // @[Top.scala 416:21]
  wire [31:0] n65_I0_15; // @[Top.scala 416:21]
  wire [31:0] n65_I1_0; // @[Top.scala 416:21]
  wire [31:0] n65_I1_1; // @[Top.scala 416:21]
  wire [31:0] n65_I1_2; // @[Top.scala 416:21]
  wire [31:0] n65_I1_3; // @[Top.scala 416:21]
  wire [31:0] n65_I1_4; // @[Top.scala 416:21]
  wire [31:0] n65_I1_5; // @[Top.scala 416:21]
  wire [31:0] n65_I1_6; // @[Top.scala 416:21]
  wire [31:0] n65_I1_7; // @[Top.scala 416:21]
  wire [31:0] n65_I1_8; // @[Top.scala 416:21]
  wire [31:0] n65_I1_9; // @[Top.scala 416:21]
  wire [31:0] n65_I1_10; // @[Top.scala 416:21]
  wire [31:0] n65_I1_11; // @[Top.scala 416:21]
  wire [31:0] n65_I1_12; // @[Top.scala 416:21]
  wire [31:0] n65_I1_13; // @[Top.scala 416:21]
  wire [31:0] n65_I1_14; // @[Top.scala 416:21]
  wire [31:0] n65_I1_15; // @[Top.scala 416:21]
  wire [31:0] n65_O_0_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_0_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_1_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_1_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_2_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_2_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_3_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_3_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_4_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_4_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_5_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_5_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_6_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_6_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_7_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_7_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_8_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_8_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_9_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_9_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_10_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_10_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_11_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_11_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_12_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_12_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_13_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_13_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_14_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_14_1; // @[Top.scala 416:21]
  wire [31:0] n65_O_15_0; // @[Top.scala 416:21]
  wire [31:0] n65_O_15_1; // @[Top.scala 416:21]
  wire  n72_valid_up; // @[Top.scala 420:21]
  wire  n72_valid_down; // @[Top.scala 420:21]
  wire [31:0] n72_I0_0_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_0_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_1_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_1_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_2_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_2_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_3_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_3_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_4_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_4_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_5_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_5_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_6_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_6_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_7_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_7_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_8_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_8_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_9_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_9_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_10_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_10_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_11_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_11_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_12_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_12_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_13_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_13_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_14_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_14_1; // @[Top.scala 420:21]
  wire [31:0] n72_I0_15_0; // @[Top.scala 420:21]
  wire [31:0] n72_I0_15_1; // @[Top.scala 420:21]
  wire [31:0] n72_I1_0; // @[Top.scala 420:21]
  wire [31:0] n72_I1_1; // @[Top.scala 420:21]
  wire [31:0] n72_I1_2; // @[Top.scala 420:21]
  wire [31:0] n72_I1_3; // @[Top.scala 420:21]
  wire [31:0] n72_I1_4; // @[Top.scala 420:21]
  wire [31:0] n72_I1_5; // @[Top.scala 420:21]
  wire [31:0] n72_I1_6; // @[Top.scala 420:21]
  wire [31:0] n72_I1_7; // @[Top.scala 420:21]
  wire [31:0] n72_I1_8; // @[Top.scala 420:21]
  wire [31:0] n72_I1_9; // @[Top.scala 420:21]
  wire [31:0] n72_I1_10; // @[Top.scala 420:21]
  wire [31:0] n72_I1_11; // @[Top.scala 420:21]
  wire [31:0] n72_I1_12; // @[Top.scala 420:21]
  wire [31:0] n72_I1_13; // @[Top.scala 420:21]
  wire [31:0] n72_I1_14; // @[Top.scala 420:21]
  wire [31:0] n72_I1_15; // @[Top.scala 420:21]
  wire [31:0] n72_O_0_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_0_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_0_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_1_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_1_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_1_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_2_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_2_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_2_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_3_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_3_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_3_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_4_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_4_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_4_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_5_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_5_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_5_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_6_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_6_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_6_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_7_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_7_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_7_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_8_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_8_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_8_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_9_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_9_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_9_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_10_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_10_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_10_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_11_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_11_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_11_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_12_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_12_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_12_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_13_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_13_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_13_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_14_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_14_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_14_2; // @[Top.scala 420:21]
  wire [31:0] n72_O_15_0; // @[Top.scala 420:21]
  wire [31:0] n72_O_15_1; // @[Top.scala 420:21]
  wire [31:0] n72_O_15_2; // @[Top.scala 420:21]
  wire  n81_valid_up; // @[Top.scala 424:21]
  wire  n81_valid_down; // @[Top.scala 424:21]
  wire [31:0] n81_I_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_1_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_1_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_1_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_2_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_2_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_2_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_3_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_3_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_3_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_4_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_4_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_4_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_5_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_5_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_5_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_6_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_6_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_6_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_7_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_7_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_7_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_8_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_8_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_8_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_9_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_9_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_9_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_10_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_10_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_10_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_11_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_11_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_11_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_12_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_12_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_12_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_13_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_13_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_13_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_14_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_14_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_14_2; // @[Top.scala 424:21]
  wire [31:0] n81_I_15_0; // @[Top.scala 424:21]
  wire [31:0] n81_I_15_1; // @[Top.scala 424:21]
  wire [31:0] n81_I_15_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_0_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_0_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_0_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_1_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_1_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_1_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_2_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_2_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_2_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_3_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_3_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_3_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_4_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_4_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_4_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_5_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_5_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_5_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_6_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_6_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_6_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_7_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_7_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_7_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_8_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_8_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_8_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_9_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_9_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_9_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_10_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_10_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_10_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_11_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_11_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_11_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_12_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_12_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_12_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_13_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_13_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_13_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_14_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_14_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_14_0_2; // @[Top.scala 424:21]
  wire [31:0] n81_O_15_0_0; // @[Top.scala 424:21]
  wire [31:0] n81_O_15_0_1; // @[Top.scala 424:21]
  wire [31:0] n81_O_15_0_2; // @[Top.scala 424:21]
  wire  n88_valid_up; // @[Top.scala 427:21]
  wire  n88_valid_down; // @[Top.scala 427:21]
  wire [31:0] n88_I_0_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_0_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_0_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_1_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_1_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_1_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_2_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_2_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_2_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_3_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_3_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_3_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_4_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_4_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_4_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_5_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_5_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_5_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_6_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_6_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_6_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_7_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_7_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_7_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_8_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_8_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_8_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_9_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_9_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_9_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_10_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_10_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_10_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_11_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_11_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_11_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_12_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_12_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_12_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_13_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_13_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_13_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_14_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_14_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_14_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_I_15_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_I_15_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_I_15_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_0_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_0_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_0_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_1_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_1_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_1_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_2_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_2_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_2_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_3_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_3_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_3_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_4_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_4_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_4_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_5_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_5_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_5_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_6_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_6_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_6_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_7_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_7_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_7_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_8_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_8_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_8_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_9_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_9_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_9_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_10_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_10_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_10_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_11_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_11_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_11_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_12_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_12_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_12_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_13_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_13_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_13_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_14_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_14_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_14_2; // @[Top.scala 427:21]
  wire [31:0] n88_O_15_0; // @[Top.scala 427:21]
  wire [31:0] n88_O_15_1; // @[Top.scala 427:21]
  wire [31:0] n88_O_15_2; // @[Top.scala 427:21]
  wire  n89_valid_up; // @[Top.scala 430:21]
  wire  n89_valid_down; // @[Top.scala 430:21]
  wire [31:0] n89_I0_0_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_0_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_0_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_0_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_0_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_0_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_1_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_1_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_1_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_1_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_1_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_1_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_2_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_2_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_2_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_2_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_2_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_2_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_3_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_3_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_3_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_3_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_3_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_3_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_4_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_4_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_4_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_4_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_4_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_4_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_5_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_5_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_5_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_5_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_5_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_5_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_6_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_6_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_6_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_6_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_6_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_6_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_7_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_7_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_7_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_7_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_7_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_7_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_8_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_8_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_8_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_8_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_8_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_8_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_9_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_9_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_9_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_9_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_9_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_9_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_10_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_10_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_10_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_10_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_10_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_10_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_11_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_11_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_11_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_11_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_11_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_11_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_12_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_12_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_12_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_12_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_12_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_12_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_13_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_13_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_13_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_13_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_13_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_13_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_14_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_14_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_14_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_14_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_14_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_14_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_15_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_15_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_15_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I0_15_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I0_15_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I0_15_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_3_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_3_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_3_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_4_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_4_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_4_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_5_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_5_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_5_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_6_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_6_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_6_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_7_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_7_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_7_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_8_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_8_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_8_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_9_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_9_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_9_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_10_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_10_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_10_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_11_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_11_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_11_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_12_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_12_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_12_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_13_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_13_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_13_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_14_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_14_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_14_2; // @[Top.scala 430:21]
  wire [31:0] n89_I1_15_0; // @[Top.scala 430:21]
  wire [31:0] n89_I1_15_1; // @[Top.scala 430:21]
  wire [31:0] n89_I1_15_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_0_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_1_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_2_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_3_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_4_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_5_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_6_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_7_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_8_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_9_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_10_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_11_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_12_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_13_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_14_2_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_0_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_0_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_0_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_1_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_1_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_1_2; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_2_0; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_2_1; // @[Top.scala 430:21]
  wire [31:0] n89_O_15_2_2; // @[Top.scala 430:21]
  wire  n98_valid_up; // @[Top.scala 434:21]
  wire  n98_valid_down; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_1_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_2_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_3_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_4_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_5_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_6_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_7_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_8_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_9_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_10_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_11_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_12_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_13_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_14_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_I_15_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_0_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_1_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_2_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_3_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_4_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_5_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_6_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_7_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_8_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_9_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_10_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_11_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_12_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_13_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_14_0_2_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_0_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_0_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_0_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_1_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_1_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_1_2; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_2_0; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_2_1; // @[Top.scala 434:21]
  wire [31:0] n98_O_15_0_2_2; // @[Top.scala 434:21]
  wire  n105_valid_up; // @[Top.scala 437:22]
  wire  n105_valid_down; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_0_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_1_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_2_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_3_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_4_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_5_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_6_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_7_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_8_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_9_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_10_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_11_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_12_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_13_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_14_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_I_15_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_0_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_1_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_2_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_3_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_4_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_5_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_6_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_7_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_8_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_9_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_10_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_11_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_12_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_13_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_14_2_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_0_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_0_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_0_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_1_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_1_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_1_2; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_2_0; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_2_1; // @[Top.scala 437:22]
  wire [31:0] n105_O_15_2_2; // @[Top.scala 437:22]
  wire  n106_valid_up; // @[Top.scala 440:22]
  wire  n106_valid_down; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_0_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_1_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_2_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_3_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_4_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_5_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_6_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_7_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_8_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_9_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_10_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_11_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_12_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_13_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_14_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_I_15_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_0_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_1_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_2_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_3_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_4_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_5_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_6_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_7_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_8_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_9_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_10_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_11_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_12_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_13_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_14_2_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_0_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_0_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_0_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_1_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_1_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_1_2; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_2_0; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_2_1; // @[Top.scala 440:22]
  wire [31:0] n106_O_15_2_2; // @[Top.scala 440:22]
  wire  n443_clock; // @[Top.scala 443:22]
  wire  n443_reset; // @[Top.scala 443:22]
  wire  n443_valid_up; // @[Top.scala 443:22]
  wire  n443_valid_down; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_0_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_1_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_2_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_3_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_4_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_5_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_6_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_7_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_8_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_9_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_10_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_11_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_12_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_13_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_14_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_0_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_0_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_0_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_1_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_1_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_1_2; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_2_0; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_2_1; // @[Top.scala 443:22]
  wire [31:0] n443_I_15_2_2; // @[Top.scala 443:22]
  wire [31:0] n443_O_0_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_0_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_0_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_1_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_1_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_1_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_2_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_2_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_2_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_3_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_3_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_3_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_4_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_4_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_4_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_5_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_5_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_5_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_6_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_6_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_6_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_7_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_7_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_7_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_8_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_8_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_8_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_9_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_9_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_9_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_10_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_10_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_10_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_11_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_11_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_11_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_12_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_12_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_12_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_13_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_13_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_13_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_14_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_14_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_14_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire [31:0] n443_O_15_0_0_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_15_0_0_t1b_t0b; // @[Top.scala 443:22]
  wire [31:0] n443_O_15_0_0_t1b_t1b; // @[Top.scala 443:22]
  wire  n444_valid_up; // @[Top.scala 446:22]
  wire  n444_valid_down; // @[Top.scala 446:22]
  wire [31:0] n444_I_0_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_0_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_0_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_1_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_1_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_1_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_2_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_2_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_2_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_3_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_3_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_3_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_4_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_4_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_4_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_5_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_5_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_5_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_6_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_6_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_6_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_7_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_7_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_7_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_8_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_8_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_8_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_9_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_9_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_9_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_10_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_10_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_10_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_11_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_11_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_11_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_12_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_12_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_12_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_13_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_13_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_13_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_14_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_14_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_14_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_I_15_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_15_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_I_15_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_0_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_0_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_0_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_1_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_1_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_1_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_2_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_2_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_2_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_3_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_3_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_3_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_4_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_4_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_4_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_5_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_5_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_5_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_6_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_6_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_6_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_7_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_7_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_7_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_8_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_8_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_8_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_9_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_9_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_9_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_10_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_10_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_10_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_11_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_11_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_11_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_12_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_12_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_12_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_13_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_13_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_13_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_14_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_14_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_14_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire [31:0] n444_O_15_0_0_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_15_0_0_t1b_t0b; // @[Top.scala 446:22]
  wire [31:0] n444_O_15_0_0_t1b_t1b; // @[Top.scala 446:22]
  wire  n445_valid_up; // @[Top.scala 449:22]
  wire  n445_valid_down; // @[Top.scala 449:22]
  wire [31:0] n445_I_0_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_0_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_0_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_1_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_1_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_1_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_2_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_2_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_2_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_3_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_3_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_3_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_4_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_4_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_4_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_5_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_5_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_5_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_6_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_6_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_6_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_7_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_7_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_7_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_8_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_8_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_8_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_9_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_9_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_9_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_10_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_10_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_10_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_11_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_11_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_11_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_12_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_12_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_12_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_13_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_13_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_13_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_14_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_14_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_14_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_I_15_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_15_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_I_15_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_0_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_0_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_0_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_1_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_1_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_1_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_2_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_2_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_2_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_3_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_3_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_3_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_4_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_4_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_4_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_5_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_5_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_5_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_6_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_6_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_6_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_7_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_7_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_7_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_8_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_8_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_8_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_9_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_9_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_9_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_10_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_10_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_10_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_11_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_11_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_11_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_12_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_12_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_12_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_13_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_13_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_13_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_14_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_14_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_14_0_t1b_t1b; // @[Top.scala 449:22]
  wire [31:0] n445_O_15_0_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_15_0_t1b_t0b; // @[Top.scala 449:22]
  wire [31:0] n445_O_15_0_t1b_t1b; // @[Top.scala 449:22]
  wire  n446_valid_up; // @[Top.scala 452:22]
  wire  n446_valid_down; // @[Top.scala 452:22]
  wire [31:0] n446_I_0_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_0_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_0_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_1_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_1_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_1_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_2_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_2_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_2_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_3_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_3_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_3_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_4_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_4_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_4_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_5_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_5_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_5_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_6_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_6_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_6_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_7_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_7_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_7_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_8_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_8_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_8_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_9_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_9_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_9_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_10_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_10_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_10_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_11_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_11_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_11_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_12_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_12_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_12_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_13_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_13_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_13_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_14_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_14_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_14_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_I_15_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_15_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_I_15_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_0_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_0_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_0_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_1_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_1_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_1_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_2_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_2_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_2_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_3_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_3_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_3_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_4_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_4_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_4_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_5_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_5_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_5_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_6_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_6_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_6_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_7_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_7_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_7_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_8_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_8_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_8_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_9_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_9_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_9_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_10_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_10_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_10_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_11_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_11_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_11_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_12_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_12_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_12_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_13_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_13_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_13_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_14_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_14_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_14_t1b_t1b; // @[Top.scala 452:22]
  wire [31:0] n446_O_15_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_15_t1b_t0b; // @[Top.scala 452:22]
  wire [31:0] n446_O_15_t1b_t1b; // @[Top.scala 452:22]
  wire  n447_clock; // @[Top.scala 455:22]
  wire  n447_reset; // @[Top.scala 455:22]
  wire  n447_valid_up; // @[Top.scala 455:22]
  wire  n447_valid_down; // @[Top.scala 455:22]
  wire [31:0] n447_I_0_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_0_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_0_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_1_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_1_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_1_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_2_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_2_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_2_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_3_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_3_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_3_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_4_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_4_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_4_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_5_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_5_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_5_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_6_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_6_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_6_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_7_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_7_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_7_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_8_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_8_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_8_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_9_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_9_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_9_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_10_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_10_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_10_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_11_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_11_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_11_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_12_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_12_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_12_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_13_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_13_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_13_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_14_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_14_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_14_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_I_15_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_15_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_I_15_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_0_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_0_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_0_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_1_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_1_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_1_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_2_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_2_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_2_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_3_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_3_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_3_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_4_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_4_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_4_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_5_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_5_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_5_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_6_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_6_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_6_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_7_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_7_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_7_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_8_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_8_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_8_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_9_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_9_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_9_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_10_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_10_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_10_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_11_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_11_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_11_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_12_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_12_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_12_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_13_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_13_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_13_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_14_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_14_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_14_t1b_t1b; // @[Top.scala 455:22]
  wire [31:0] n447_O_15_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_15_t1b_t0b; // @[Top.scala 455:22]
  wire [31:0] n447_O_15_t1b_t1b; // @[Top.scala 455:22]
  wire  n448_clock; // @[Top.scala 458:22]
  wire  n448_reset; // @[Top.scala 458:22]
  wire  n448_valid_up; // @[Top.scala 458:22]
  wire  n448_valid_down; // @[Top.scala 458:22]
  wire [31:0] n448_I_0_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_0_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_0_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_1_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_1_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_1_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_2_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_2_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_2_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_3_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_3_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_3_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_4_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_4_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_4_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_5_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_5_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_5_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_6_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_6_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_6_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_7_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_7_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_7_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_8_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_8_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_8_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_9_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_9_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_9_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_10_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_10_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_10_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_11_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_11_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_11_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_12_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_12_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_12_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_13_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_13_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_13_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_14_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_14_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_14_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_I_15_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_15_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_I_15_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_0_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_0_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_0_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_1_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_1_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_1_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_2_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_2_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_2_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_3_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_3_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_3_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_4_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_4_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_4_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_5_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_5_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_5_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_6_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_6_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_6_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_7_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_7_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_7_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_8_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_8_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_8_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_9_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_9_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_9_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_10_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_10_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_10_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_11_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_11_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_11_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_12_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_12_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_12_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_13_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_13_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_13_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_14_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_14_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_14_t1b_t1b; // @[Top.scala 458:22]
  wire [31:0] n448_O_15_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_15_t1b_t0b; // @[Top.scala 458:22]
  wire [31:0] n448_O_15_t1b_t1b; // @[Top.scala 458:22]
  wire  n449_clock; // @[Top.scala 461:22]
  wire  n449_reset; // @[Top.scala 461:22]
  wire  n449_valid_up; // @[Top.scala 461:22]
  wire  n449_valid_down; // @[Top.scala 461:22]
  wire [31:0] n449_I_0_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_0_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_0_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_1_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_1_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_1_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_2_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_2_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_2_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_3_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_3_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_3_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_4_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_4_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_4_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_5_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_5_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_5_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_6_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_6_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_6_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_7_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_7_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_7_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_8_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_8_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_8_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_9_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_9_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_9_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_10_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_10_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_10_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_11_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_11_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_11_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_12_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_12_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_12_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_13_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_13_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_13_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_14_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_14_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_14_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_I_15_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_15_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_I_15_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_0_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_0_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_0_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_1_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_1_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_1_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_2_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_2_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_2_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_3_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_3_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_3_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_4_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_4_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_4_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_5_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_5_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_5_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_6_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_6_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_6_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_7_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_7_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_7_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_8_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_8_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_8_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_9_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_9_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_9_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_10_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_10_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_10_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_11_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_11_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_11_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_12_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_12_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_12_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_13_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_13_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_13_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_14_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_14_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_14_t1b_t1b; // @[Top.scala 461:22]
  wire [31:0] n449_O_15_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_15_t1b_t0b; // @[Top.scala 461:22]
  wire [31:0] n449_O_15_t1b_t1b; // @[Top.scala 461:22]
  FIFO n1 ( // @[Top.scala 357:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .I_8(n1_I_8),
    .I_9(n1_I_9),
    .I_10(n1_I_10),
    .I_11(n1_I_11),
    .I_12(n1_I_12),
    .I_13(n1_I_13),
    .I_14(n1_I_14),
    .I_15(n1_I_15),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7),
    .O_8(n1_O_8),
    .O_9(n1_O_9),
    .O_10(n1_O_10),
    .O_11(n1_O_11),
    .O_12(n1_O_12),
    .O_13(n1_O_13),
    .O_14(n1_O_14),
    .O_15(n1_O_15)
  );
  ShiftTS n2 ( // @[Top.scala 360:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .I_4(n2_I_4),
    .I_5(n2_I_5),
    .I_6(n2_I_6),
    .I_7(n2_I_7),
    .I_8(n2_I_8),
    .I_9(n2_I_9),
    .I_10(n2_I_10),
    .I_11(n2_I_11),
    .I_12(n2_I_12),
    .I_13(n2_I_13),
    .I_14(n2_I_14),
    .I_15(n2_I_15),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3),
    .O_4(n2_O_4),
    .O_5(n2_O_5),
    .O_6(n2_O_6),
    .O_7(n2_O_7),
    .O_8(n2_O_8),
    .O_9(n2_O_9),
    .O_10(n2_O_10),
    .O_11(n2_O_11),
    .O_12(n2_O_12),
    .O_13(n2_O_13),
    .O_14(n2_O_14),
    .O_15(n2_O_15)
  );
  ShiftTS n3 ( // @[Top.scala 363:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .I_4(n3_I_4),
    .I_5(n3_I_5),
    .I_6(n3_I_6),
    .I_7(n3_I_7),
    .I_8(n3_I_8),
    .I_9(n3_I_9),
    .I_10(n3_I_10),
    .I_11(n3_I_11),
    .I_12(n3_I_12),
    .I_13(n3_I_13),
    .I_14(n3_I_14),
    .I_15(n3_I_15),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3),
    .O_4(n3_O_4),
    .O_5(n3_O_5),
    .O_6(n3_O_6),
    .O_7(n3_O_7),
    .O_8(n3_O_8),
    .O_9(n3_O_9),
    .O_10(n3_O_10),
    .O_11(n3_O_11),
    .O_12(n3_O_12),
    .O_13(n3_O_13),
    .O_14(n3_O_14),
    .O_15(n3_O_15)
  );
  ShiftTS_2 n4 ( // @[Top.scala 366:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .I_4(n4_I_4),
    .I_5(n4_I_5),
    .I_6(n4_I_6),
    .I_7(n4_I_7),
    .I_8(n4_I_8),
    .I_9(n4_I_9),
    .I_10(n4_I_10),
    .I_11(n4_I_11),
    .I_12(n4_I_12),
    .I_13(n4_I_13),
    .I_14(n4_I_14),
    .I_15(n4_I_15),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3),
    .O_4(n4_O_4),
    .O_5(n4_O_5),
    .O_6(n4_O_6),
    .O_7(n4_O_7),
    .O_8(n4_O_8),
    .O_9(n4_O_9),
    .O_10(n4_O_10),
    .O_11(n4_O_11),
    .O_12(n4_O_12),
    .O_13(n4_O_13),
    .O_14(n4_O_14),
    .O_15(n4_O_15)
  );
  ShiftTS_2 n5 ( // @[Top.scala 369:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .I_4(n5_I_4),
    .I_5(n5_I_5),
    .I_6(n5_I_6),
    .I_7(n5_I_7),
    .I_8(n5_I_8),
    .I_9(n5_I_9),
    .I_10(n5_I_10),
    .I_11(n5_I_11),
    .I_12(n5_I_12),
    .I_13(n5_I_13),
    .I_14(n5_I_14),
    .I_15(n5_I_15),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3),
    .O_4(n5_O_4),
    .O_5(n5_O_5),
    .O_6(n5_O_6),
    .O_7(n5_O_7),
    .O_8(n5_O_8),
    .O_9(n5_O_9),
    .O_10(n5_O_10),
    .O_11(n5_O_11),
    .O_12(n5_O_12),
    .O_13(n5_O_13),
    .O_14(n5_O_14),
    .O_15(n5_O_15)
  );
  Map2T n6 ( // @[Top.scala 372:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I0_2(n6_I0_2),
    .I0_3(n6_I0_3),
    .I0_4(n6_I0_4),
    .I0_5(n6_I0_5),
    .I0_6(n6_I0_6),
    .I0_7(n6_I0_7),
    .I0_8(n6_I0_8),
    .I0_9(n6_I0_9),
    .I0_10(n6_I0_10),
    .I0_11(n6_I0_11),
    .I0_12(n6_I0_12),
    .I0_13(n6_I0_13),
    .I0_14(n6_I0_14),
    .I0_15(n6_I0_15),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .I1_2(n6_I1_2),
    .I1_3(n6_I1_3),
    .I1_4(n6_I1_4),
    .I1_5(n6_I1_5),
    .I1_6(n6_I1_6),
    .I1_7(n6_I1_7),
    .I1_8(n6_I1_8),
    .I1_9(n6_I1_9),
    .I1_10(n6_I1_10),
    .I1_11(n6_I1_11),
    .I1_12(n6_I1_12),
    .I1_13(n6_I1_13),
    .I1_14(n6_I1_14),
    .I1_15(n6_I1_15),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1),
    .O_2_0(n6_O_2_0),
    .O_2_1(n6_O_2_1),
    .O_3_0(n6_O_3_0),
    .O_3_1(n6_O_3_1),
    .O_4_0(n6_O_4_0),
    .O_4_1(n6_O_4_1),
    .O_5_0(n6_O_5_0),
    .O_5_1(n6_O_5_1),
    .O_6_0(n6_O_6_0),
    .O_6_1(n6_O_6_1),
    .O_7_0(n6_O_7_0),
    .O_7_1(n6_O_7_1),
    .O_8_0(n6_O_8_0),
    .O_8_1(n6_O_8_1),
    .O_9_0(n6_O_9_0),
    .O_9_1(n6_O_9_1),
    .O_10_0(n6_O_10_0),
    .O_10_1(n6_O_10_1),
    .O_11_0(n6_O_11_0),
    .O_11_1(n6_O_11_1),
    .O_12_0(n6_O_12_0),
    .O_12_1(n6_O_12_1),
    .O_13_0(n6_O_13_0),
    .O_13_1(n6_O_13_1),
    .O_14_0(n6_O_14_0),
    .O_14_1(n6_O_14_1),
    .O_15_0(n6_O_15_0),
    .O_15_1(n6_O_15_1)
  );
  Map2T_1 n13 ( // @[Top.scala 376:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0_0(n13_I0_0_0),
    .I0_0_1(n13_I0_0_1),
    .I0_1_0(n13_I0_1_0),
    .I0_1_1(n13_I0_1_1),
    .I0_2_0(n13_I0_2_0),
    .I0_2_1(n13_I0_2_1),
    .I0_3_0(n13_I0_3_0),
    .I0_3_1(n13_I0_3_1),
    .I0_4_0(n13_I0_4_0),
    .I0_4_1(n13_I0_4_1),
    .I0_5_0(n13_I0_5_0),
    .I0_5_1(n13_I0_5_1),
    .I0_6_0(n13_I0_6_0),
    .I0_6_1(n13_I0_6_1),
    .I0_7_0(n13_I0_7_0),
    .I0_7_1(n13_I0_7_1),
    .I0_8_0(n13_I0_8_0),
    .I0_8_1(n13_I0_8_1),
    .I0_9_0(n13_I0_9_0),
    .I0_9_1(n13_I0_9_1),
    .I0_10_0(n13_I0_10_0),
    .I0_10_1(n13_I0_10_1),
    .I0_11_0(n13_I0_11_0),
    .I0_11_1(n13_I0_11_1),
    .I0_12_0(n13_I0_12_0),
    .I0_12_1(n13_I0_12_1),
    .I0_13_0(n13_I0_13_0),
    .I0_13_1(n13_I0_13_1),
    .I0_14_0(n13_I0_14_0),
    .I0_14_1(n13_I0_14_1),
    .I0_15_0(n13_I0_15_0),
    .I0_15_1(n13_I0_15_1),
    .I1_0(n13_I1_0),
    .I1_1(n13_I1_1),
    .I1_2(n13_I1_2),
    .I1_3(n13_I1_3),
    .I1_4(n13_I1_4),
    .I1_5(n13_I1_5),
    .I1_6(n13_I1_6),
    .I1_7(n13_I1_7),
    .I1_8(n13_I1_8),
    .I1_9(n13_I1_9),
    .I1_10(n13_I1_10),
    .I1_11(n13_I1_11),
    .I1_12(n13_I1_12),
    .I1_13(n13_I1_13),
    .I1_14(n13_I1_14),
    .I1_15(n13_I1_15),
    .O_0_0(n13_O_0_0),
    .O_0_1(n13_O_0_1),
    .O_0_2(n13_O_0_2),
    .O_1_0(n13_O_1_0),
    .O_1_1(n13_O_1_1),
    .O_1_2(n13_O_1_2),
    .O_2_0(n13_O_2_0),
    .O_2_1(n13_O_2_1),
    .O_2_2(n13_O_2_2),
    .O_3_0(n13_O_3_0),
    .O_3_1(n13_O_3_1),
    .O_3_2(n13_O_3_2),
    .O_4_0(n13_O_4_0),
    .O_4_1(n13_O_4_1),
    .O_4_2(n13_O_4_2),
    .O_5_0(n13_O_5_0),
    .O_5_1(n13_O_5_1),
    .O_5_2(n13_O_5_2),
    .O_6_0(n13_O_6_0),
    .O_6_1(n13_O_6_1),
    .O_6_2(n13_O_6_2),
    .O_7_0(n13_O_7_0),
    .O_7_1(n13_O_7_1),
    .O_7_2(n13_O_7_2),
    .O_8_0(n13_O_8_0),
    .O_8_1(n13_O_8_1),
    .O_8_2(n13_O_8_2),
    .O_9_0(n13_O_9_0),
    .O_9_1(n13_O_9_1),
    .O_9_2(n13_O_9_2),
    .O_10_0(n13_O_10_0),
    .O_10_1(n13_O_10_1),
    .O_10_2(n13_O_10_2),
    .O_11_0(n13_O_11_0),
    .O_11_1(n13_O_11_1),
    .O_11_2(n13_O_11_2),
    .O_12_0(n13_O_12_0),
    .O_12_1(n13_O_12_1),
    .O_12_2(n13_O_12_2),
    .O_13_0(n13_O_13_0),
    .O_13_1(n13_O_13_1),
    .O_13_2(n13_O_13_2),
    .O_14_0(n13_O_14_0),
    .O_14_1(n13_O_14_1),
    .O_14_2(n13_O_14_2),
    .O_15_0(n13_O_15_0),
    .O_15_1(n13_O_15_1),
    .O_15_2(n13_O_15_2)
  );
  MapT n22 ( // @[Top.scala 380:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I_0_0(n22_I_0_0),
    .I_0_1(n22_I_0_1),
    .I_0_2(n22_I_0_2),
    .I_1_0(n22_I_1_0),
    .I_1_1(n22_I_1_1),
    .I_1_2(n22_I_1_2),
    .I_2_0(n22_I_2_0),
    .I_2_1(n22_I_2_1),
    .I_2_2(n22_I_2_2),
    .I_3_0(n22_I_3_0),
    .I_3_1(n22_I_3_1),
    .I_3_2(n22_I_3_2),
    .I_4_0(n22_I_4_0),
    .I_4_1(n22_I_4_1),
    .I_4_2(n22_I_4_2),
    .I_5_0(n22_I_5_0),
    .I_5_1(n22_I_5_1),
    .I_5_2(n22_I_5_2),
    .I_6_0(n22_I_6_0),
    .I_6_1(n22_I_6_1),
    .I_6_2(n22_I_6_2),
    .I_7_0(n22_I_7_0),
    .I_7_1(n22_I_7_1),
    .I_7_2(n22_I_7_2),
    .I_8_0(n22_I_8_0),
    .I_8_1(n22_I_8_1),
    .I_8_2(n22_I_8_2),
    .I_9_0(n22_I_9_0),
    .I_9_1(n22_I_9_1),
    .I_9_2(n22_I_9_2),
    .I_10_0(n22_I_10_0),
    .I_10_1(n22_I_10_1),
    .I_10_2(n22_I_10_2),
    .I_11_0(n22_I_11_0),
    .I_11_1(n22_I_11_1),
    .I_11_2(n22_I_11_2),
    .I_12_0(n22_I_12_0),
    .I_12_1(n22_I_12_1),
    .I_12_2(n22_I_12_2),
    .I_13_0(n22_I_13_0),
    .I_13_1(n22_I_13_1),
    .I_13_2(n22_I_13_2),
    .I_14_0(n22_I_14_0),
    .I_14_1(n22_I_14_1),
    .I_14_2(n22_I_14_2),
    .I_15_0(n22_I_15_0),
    .I_15_1(n22_I_15_1),
    .I_15_2(n22_I_15_2),
    .O_0_0_0(n22_O_0_0_0),
    .O_0_0_1(n22_O_0_0_1),
    .O_0_0_2(n22_O_0_0_2),
    .O_1_0_0(n22_O_1_0_0),
    .O_1_0_1(n22_O_1_0_1),
    .O_1_0_2(n22_O_1_0_2),
    .O_2_0_0(n22_O_2_0_0),
    .O_2_0_1(n22_O_2_0_1),
    .O_2_0_2(n22_O_2_0_2),
    .O_3_0_0(n22_O_3_0_0),
    .O_3_0_1(n22_O_3_0_1),
    .O_3_0_2(n22_O_3_0_2),
    .O_4_0_0(n22_O_4_0_0),
    .O_4_0_1(n22_O_4_0_1),
    .O_4_0_2(n22_O_4_0_2),
    .O_5_0_0(n22_O_5_0_0),
    .O_5_0_1(n22_O_5_0_1),
    .O_5_0_2(n22_O_5_0_2),
    .O_6_0_0(n22_O_6_0_0),
    .O_6_0_1(n22_O_6_0_1),
    .O_6_0_2(n22_O_6_0_2),
    .O_7_0_0(n22_O_7_0_0),
    .O_7_0_1(n22_O_7_0_1),
    .O_7_0_2(n22_O_7_0_2),
    .O_8_0_0(n22_O_8_0_0),
    .O_8_0_1(n22_O_8_0_1),
    .O_8_0_2(n22_O_8_0_2),
    .O_9_0_0(n22_O_9_0_0),
    .O_9_0_1(n22_O_9_0_1),
    .O_9_0_2(n22_O_9_0_2),
    .O_10_0_0(n22_O_10_0_0),
    .O_10_0_1(n22_O_10_0_1),
    .O_10_0_2(n22_O_10_0_2),
    .O_11_0_0(n22_O_11_0_0),
    .O_11_0_1(n22_O_11_0_1),
    .O_11_0_2(n22_O_11_0_2),
    .O_12_0_0(n22_O_12_0_0),
    .O_12_0_1(n22_O_12_0_1),
    .O_12_0_2(n22_O_12_0_2),
    .O_13_0_0(n22_O_13_0_0),
    .O_13_0_1(n22_O_13_0_1),
    .O_13_0_2(n22_O_13_0_2),
    .O_14_0_0(n22_O_14_0_0),
    .O_14_0_1(n22_O_14_0_1),
    .O_14_0_2(n22_O_14_0_2),
    .O_15_0_0(n22_O_15_0_0),
    .O_15_0_1(n22_O_15_0_1),
    .O_15_0_2(n22_O_15_0_2)
  );
  MapT_1 n29 ( // @[Top.scala 383:21]
    .valid_up(n29_valid_up),
    .valid_down(n29_valid_down),
    .I_0_0_0(n29_I_0_0_0),
    .I_0_0_1(n29_I_0_0_1),
    .I_0_0_2(n29_I_0_0_2),
    .I_1_0_0(n29_I_1_0_0),
    .I_1_0_1(n29_I_1_0_1),
    .I_1_0_2(n29_I_1_0_2),
    .I_2_0_0(n29_I_2_0_0),
    .I_2_0_1(n29_I_2_0_1),
    .I_2_0_2(n29_I_2_0_2),
    .I_3_0_0(n29_I_3_0_0),
    .I_3_0_1(n29_I_3_0_1),
    .I_3_0_2(n29_I_3_0_2),
    .I_4_0_0(n29_I_4_0_0),
    .I_4_0_1(n29_I_4_0_1),
    .I_4_0_2(n29_I_4_0_2),
    .I_5_0_0(n29_I_5_0_0),
    .I_5_0_1(n29_I_5_0_1),
    .I_5_0_2(n29_I_5_0_2),
    .I_6_0_0(n29_I_6_0_0),
    .I_6_0_1(n29_I_6_0_1),
    .I_6_0_2(n29_I_6_0_2),
    .I_7_0_0(n29_I_7_0_0),
    .I_7_0_1(n29_I_7_0_1),
    .I_7_0_2(n29_I_7_0_2),
    .I_8_0_0(n29_I_8_0_0),
    .I_8_0_1(n29_I_8_0_1),
    .I_8_0_2(n29_I_8_0_2),
    .I_9_0_0(n29_I_9_0_0),
    .I_9_0_1(n29_I_9_0_1),
    .I_9_0_2(n29_I_9_0_2),
    .I_10_0_0(n29_I_10_0_0),
    .I_10_0_1(n29_I_10_0_1),
    .I_10_0_2(n29_I_10_0_2),
    .I_11_0_0(n29_I_11_0_0),
    .I_11_0_1(n29_I_11_0_1),
    .I_11_0_2(n29_I_11_0_2),
    .I_12_0_0(n29_I_12_0_0),
    .I_12_0_1(n29_I_12_0_1),
    .I_12_0_2(n29_I_12_0_2),
    .I_13_0_0(n29_I_13_0_0),
    .I_13_0_1(n29_I_13_0_1),
    .I_13_0_2(n29_I_13_0_2),
    .I_14_0_0(n29_I_14_0_0),
    .I_14_0_1(n29_I_14_0_1),
    .I_14_0_2(n29_I_14_0_2),
    .I_15_0_0(n29_I_15_0_0),
    .I_15_0_1(n29_I_15_0_1),
    .I_15_0_2(n29_I_15_0_2),
    .O_0_0(n29_O_0_0),
    .O_0_1(n29_O_0_1),
    .O_0_2(n29_O_0_2),
    .O_1_0(n29_O_1_0),
    .O_1_1(n29_O_1_1),
    .O_1_2(n29_O_1_2),
    .O_2_0(n29_O_2_0),
    .O_2_1(n29_O_2_1),
    .O_2_2(n29_O_2_2),
    .O_3_0(n29_O_3_0),
    .O_3_1(n29_O_3_1),
    .O_3_2(n29_O_3_2),
    .O_4_0(n29_O_4_0),
    .O_4_1(n29_O_4_1),
    .O_4_2(n29_O_4_2),
    .O_5_0(n29_O_5_0),
    .O_5_1(n29_O_5_1),
    .O_5_2(n29_O_5_2),
    .O_6_0(n29_O_6_0),
    .O_6_1(n29_O_6_1),
    .O_6_2(n29_O_6_2),
    .O_7_0(n29_O_7_0),
    .O_7_1(n29_O_7_1),
    .O_7_2(n29_O_7_2),
    .O_8_0(n29_O_8_0),
    .O_8_1(n29_O_8_1),
    .O_8_2(n29_O_8_2),
    .O_9_0(n29_O_9_0),
    .O_9_1(n29_O_9_1),
    .O_9_2(n29_O_9_2),
    .O_10_0(n29_O_10_0),
    .O_10_1(n29_O_10_1),
    .O_10_2(n29_O_10_2),
    .O_11_0(n29_O_11_0),
    .O_11_1(n29_O_11_1),
    .O_11_2(n29_O_11_2),
    .O_12_0(n29_O_12_0),
    .O_12_1(n29_O_12_1),
    .O_12_2(n29_O_12_2),
    .O_13_0(n29_O_13_0),
    .O_13_1(n29_O_13_1),
    .O_13_2(n29_O_13_2),
    .O_14_0(n29_O_14_0),
    .O_14_1(n29_O_14_1),
    .O_14_2(n29_O_14_2),
    .O_15_0(n29_O_15_0),
    .O_15_1(n29_O_15_1),
    .O_15_2(n29_O_15_2)
  );
  ShiftTS_2 n30 ( // @[Top.scala 386:21]
    .clock(n30_clock),
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0(n30_I_0),
    .I_1(n30_I_1),
    .I_2(n30_I_2),
    .I_3(n30_I_3),
    .I_4(n30_I_4),
    .I_5(n30_I_5),
    .I_6(n30_I_6),
    .I_7(n30_I_7),
    .I_8(n30_I_8),
    .I_9(n30_I_9),
    .I_10(n30_I_10),
    .I_11(n30_I_11),
    .I_12(n30_I_12),
    .I_13(n30_I_13),
    .I_14(n30_I_14),
    .I_15(n30_I_15),
    .O_0(n30_O_0),
    .O_1(n30_O_1),
    .O_2(n30_O_2),
    .O_3(n30_O_3),
    .O_4(n30_O_4),
    .O_5(n30_O_5),
    .O_6(n30_O_6),
    .O_7(n30_O_7),
    .O_8(n30_O_8),
    .O_9(n30_O_9),
    .O_10(n30_O_10),
    .O_11(n30_O_11),
    .O_12(n30_O_12),
    .O_13(n30_O_13),
    .O_14(n30_O_14),
    .O_15(n30_O_15)
  );
  ShiftTS_2 n31 ( // @[Top.scala 389:21]
    .clock(n31_clock),
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0(n31_I_0),
    .I_1(n31_I_1),
    .I_2(n31_I_2),
    .I_3(n31_I_3),
    .I_4(n31_I_4),
    .I_5(n31_I_5),
    .I_6(n31_I_6),
    .I_7(n31_I_7),
    .I_8(n31_I_8),
    .I_9(n31_I_9),
    .I_10(n31_I_10),
    .I_11(n31_I_11),
    .I_12(n31_I_12),
    .I_13(n31_I_13),
    .I_14(n31_I_14),
    .I_15(n31_I_15),
    .O_0(n31_O_0),
    .O_1(n31_O_1),
    .O_2(n31_O_2),
    .O_3(n31_O_3),
    .O_4(n31_O_4),
    .O_5(n31_O_5),
    .O_6(n31_O_6),
    .O_7(n31_O_7),
    .O_8(n31_O_8),
    .O_9(n31_O_9),
    .O_10(n31_O_10),
    .O_11(n31_O_11),
    .O_12(n31_O_12),
    .O_13(n31_O_13),
    .O_14(n31_O_14),
    .O_15(n31_O_15)
  );
  Map2T n32 ( // @[Top.scala 392:21]
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I0_0(n32_I0_0),
    .I0_1(n32_I0_1),
    .I0_2(n32_I0_2),
    .I0_3(n32_I0_3),
    .I0_4(n32_I0_4),
    .I0_5(n32_I0_5),
    .I0_6(n32_I0_6),
    .I0_7(n32_I0_7),
    .I0_8(n32_I0_8),
    .I0_9(n32_I0_9),
    .I0_10(n32_I0_10),
    .I0_11(n32_I0_11),
    .I0_12(n32_I0_12),
    .I0_13(n32_I0_13),
    .I0_14(n32_I0_14),
    .I0_15(n32_I0_15),
    .I1_0(n32_I1_0),
    .I1_1(n32_I1_1),
    .I1_2(n32_I1_2),
    .I1_3(n32_I1_3),
    .I1_4(n32_I1_4),
    .I1_5(n32_I1_5),
    .I1_6(n32_I1_6),
    .I1_7(n32_I1_7),
    .I1_8(n32_I1_8),
    .I1_9(n32_I1_9),
    .I1_10(n32_I1_10),
    .I1_11(n32_I1_11),
    .I1_12(n32_I1_12),
    .I1_13(n32_I1_13),
    .I1_14(n32_I1_14),
    .I1_15(n32_I1_15),
    .O_0_0(n32_O_0_0),
    .O_0_1(n32_O_0_1),
    .O_1_0(n32_O_1_0),
    .O_1_1(n32_O_1_1),
    .O_2_0(n32_O_2_0),
    .O_2_1(n32_O_2_1),
    .O_3_0(n32_O_3_0),
    .O_3_1(n32_O_3_1),
    .O_4_0(n32_O_4_0),
    .O_4_1(n32_O_4_1),
    .O_5_0(n32_O_5_0),
    .O_5_1(n32_O_5_1),
    .O_6_0(n32_O_6_0),
    .O_6_1(n32_O_6_1),
    .O_7_0(n32_O_7_0),
    .O_7_1(n32_O_7_1),
    .O_8_0(n32_O_8_0),
    .O_8_1(n32_O_8_1),
    .O_9_0(n32_O_9_0),
    .O_9_1(n32_O_9_1),
    .O_10_0(n32_O_10_0),
    .O_10_1(n32_O_10_1),
    .O_11_0(n32_O_11_0),
    .O_11_1(n32_O_11_1),
    .O_12_0(n32_O_12_0),
    .O_12_1(n32_O_12_1),
    .O_13_0(n32_O_13_0),
    .O_13_1(n32_O_13_1),
    .O_14_0(n32_O_14_0),
    .O_14_1(n32_O_14_1),
    .O_15_0(n32_O_15_0),
    .O_15_1(n32_O_15_1)
  );
  Map2T_1 n39 ( // @[Top.scala 396:21]
    .valid_up(n39_valid_up),
    .valid_down(n39_valid_down),
    .I0_0_0(n39_I0_0_0),
    .I0_0_1(n39_I0_0_1),
    .I0_1_0(n39_I0_1_0),
    .I0_1_1(n39_I0_1_1),
    .I0_2_0(n39_I0_2_0),
    .I0_2_1(n39_I0_2_1),
    .I0_3_0(n39_I0_3_0),
    .I0_3_1(n39_I0_3_1),
    .I0_4_0(n39_I0_4_0),
    .I0_4_1(n39_I0_4_1),
    .I0_5_0(n39_I0_5_0),
    .I0_5_1(n39_I0_5_1),
    .I0_6_0(n39_I0_6_0),
    .I0_6_1(n39_I0_6_1),
    .I0_7_0(n39_I0_7_0),
    .I0_7_1(n39_I0_7_1),
    .I0_8_0(n39_I0_8_0),
    .I0_8_1(n39_I0_8_1),
    .I0_9_0(n39_I0_9_0),
    .I0_9_1(n39_I0_9_1),
    .I0_10_0(n39_I0_10_0),
    .I0_10_1(n39_I0_10_1),
    .I0_11_0(n39_I0_11_0),
    .I0_11_1(n39_I0_11_1),
    .I0_12_0(n39_I0_12_0),
    .I0_12_1(n39_I0_12_1),
    .I0_13_0(n39_I0_13_0),
    .I0_13_1(n39_I0_13_1),
    .I0_14_0(n39_I0_14_0),
    .I0_14_1(n39_I0_14_1),
    .I0_15_0(n39_I0_15_0),
    .I0_15_1(n39_I0_15_1),
    .I1_0(n39_I1_0),
    .I1_1(n39_I1_1),
    .I1_2(n39_I1_2),
    .I1_3(n39_I1_3),
    .I1_4(n39_I1_4),
    .I1_5(n39_I1_5),
    .I1_6(n39_I1_6),
    .I1_7(n39_I1_7),
    .I1_8(n39_I1_8),
    .I1_9(n39_I1_9),
    .I1_10(n39_I1_10),
    .I1_11(n39_I1_11),
    .I1_12(n39_I1_12),
    .I1_13(n39_I1_13),
    .I1_14(n39_I1_14),
    .I1_15(n39_I1_15),
    .O_0_0(n39_O_0_0),
    .O_0_1(n39_O_0_1),
    .O_0_2(n39_O_0_2),
    .O_1_0(n39_O_1_0),
    .O_1_1(n39_O_1_1),
    .O_1_2(n39_O_1_2),
    .O_2_0(n39_O_2_0),
    .O_2_1(n39_O_2_1),
    .O_2_2(n39_O_2_2),
    .O_3_0(n39_O_3_0),
    .O_3_1(n39_O_3_1),
    .O_3_2(n39_O_3_2),
    .O_4_0(n39_O_4_0),
    .O_4_1(n39_O_4_1),
    .O_4_2(n39_O_4_2),
    .O_5_0(n39_O_5_0),
    .O_5_1(n39_O_5_1),
    .O_5_2(n39_O_5_2),
    .O_6_0(n39_O_6_0),
    .O_6_1(n39_O_6_1),
    .O_6_2(n39_O_6_2),
    .O_7_0(n39_O_7_0),
    .O_7_1(n39_O_7_1),
    .O_7_2(n39_O_7_2),
    .O_8_0(n39_O_8_0),
    .O_8_1(n39_O_8_1),
    .O_8_2(n39_O_8_2),
    .O_9_0(n39_O_9_0),
    .O_9_1(n39_O_9_1),
    .O_9_2(n39_O_9_2),
    .O_10_0(n39_O_10_0),
    .O_10_1(n39_O_10_1),
    .O_10_2(n39_O_10_2),
    .O_11_0(n39_O_11_0),
    .O_11_1(n39_O_11_1),
    .O_11_2(n39_O_11_2),
    .O_12_0(n39_O_12_0),
    .O_12_1(n39_O_12_1),
    .O_12_2(n39_O_12_2),
    .O_13_0(n39_O_13_0),
    .O_13_1(n39_O_13_1),
    .O_13_2(n39_O_13_2),
    .O_14_0(n39_O_14_0),
    .O_14_1(n39_O_14_1),
    .O_14_2(n39_O_14_2),
    .O_15_0(n39_O_15_0),
    .O_15_1(n39_O_15_1),
    .O_15_2(n39_O_15_2)
  );
  MapT n48 ( // @[Top.scala 400:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I_0_0(n48_I_0_0),
    .I_0_1(n48_I_0_1),
    .I_0_2(n48_I_0_2),
    .I_1_0(n48_I_1_0),
    .I_1_1(n48_I_1_1),
    .I_1_2(n48_I_1_2),
    .I_2_0(n48_I_2_0),
    .I_2_1(n48_I_2_1),
    .I_2_2(n48_I_2_2),
    .I_3_0(n48_I_3_0),
    .I_3_1(n48_I_3_1),
    .I_3_2(n48_I_3_2),
    .I_4_0(n48_I_4_0),
    .I_4_1(n48_I_4_1),
    .I_4_2(n48_I_4_2),
    .I_5_0(n48_I_5_0),
    .I_5_1(n48_I_5_1),
    .I_5_2(n48_I_5_2),
    .I_6_0(n48_I_6_0),
    .I_6_1(n48_I_6_1),
    .I_6_2(n48_I_6_2),
    .I_7_0(n48_I_7_0),
    .I_7_1(n48_I_7_1),
    .I_7_2(n48_I_7_2),
    .I_8_0(n48_I_8_0),
    .I_8_1(n48_I_8_1),
    .I_8_2(n48_I_8_2),
    .I_9_0(n48_I_9_0),
    .I_9_1(n48_I_9_1),
    .I_9_2(n48_I_9_2),
    .I_10_0(n48_I_10_0),
    .I_10_1(n48_I_10_1),
    .I_10_2(n48_I_10_2),
    .I_11_0(n48_I_11_0),
    .I_11_1(n48_I_11_1),
    .I_11_2(n48_I_11_2),
    .I_12_0(n48_I_12_0),
    .I_12_1(n48_I_12_1),
    .I_12_2(n48_I_12_2),
    .I_13_0(n48_I_13_0),
    .I_13_1(n48_I_13_1),
    .I_13_2(n48_I_13_2),
    .I_14_0(n48_I_14_0),
    .I_14_1(n48_I_14_1),
    .I_14_2(n48_I_14_2),
    .I_15_0(n48_I_15_0),
    .I_15_1(n48_I_15_1),
    .I_15_2(n48_I_15_2),
    .O_0_0_0(n48_O_0_0_0),
    .O_0_0_1(n48_O_0_0_1),
    .O_0_0_2(n48_O_0_0_2),
    .O_1_0_0(n48_O_1_0_0),
    .O_1_0_1(n48_O_1_0_1),
    .O_1_0_2(n48_O_1_0_2),
    .O_2_0_0(n48_O_2_0_0),
    .O_2_0_1(n48_O_2_0_1),
    .O_2_0_2(n48_O_2_0_2),
    .O_3_0_0(n48_O_3_0_0),
    .O_3_0_1(n48_O_3_0_1),
    .O_3_0_2(n48_O_3_0_2),
    .O_4_0_0(n48_O_4_0_0),
    .O_4_0_1(n48_O_4_0_1),
    .O_4_0_2(n48_O_4_0_2),
    .O_5_0_0(n48_O_5_0_0),
    .O_5_0_1(n48_O_5_0_1),
    .O_5_0_2(n48_O_5_0_2),
    .O_6_0_0(n48_O_6_0_0),
    .O_6_0_1(n48_O_6_0_1),
    .O_6_0_2(n48_O_6_0_2),
    .O_7_0_0(n48_O_7_0_0),
    .O_7_0_1(n48_O_7_0_1),
    .O_7_0_2(n48_O_7_0_2),
    .O_8_0_0(n48_O_8_0_0),
    .O_8_0_1(n48_O_8_0_1),
    .O_8_0_2(n48_O_8_0_2),
    .O_9_0_0(n48_O_9_0_0),
    .O_9_0_1(n48_O_9_0_1),
    .O_9_0_2(n48_O_9_0_2),
    .O_10_0_0(n48_O_10_0_0),
    .O_10_0_1(n48_O_10_0_1),
    .O_10_0_2(n48_O_10_0_2),
    .O_11_0_0(n48_O_11_0_0),
    .O_11_0_1(n48_O_11_0_1),
    .O_11_0_2(n48_O_11_0_2),
    .O_12_0_0(n48_O_12_0_0),
    .O_12_0_1(n48_O_12_0_1),
    .O_12_0_2(n48_O_12_0_2),
    .O_13_0_0(n48_O_13_0_0),
    .O_13_0_1(n48_O_13_0_1),
    .O_13_0_2(n48_O_13_0_2),
    .O_14_0_0(n48_O_14_0_0),
    .O_14_0_1(n48_O_14_0_1),
    .O_14_0_2(n48_O_14_0_2),
    .O_15_0_0(n48_O_15_0_0),
    .O_15_0_1(n48_O_15_0_1),
    .O_15_0_2(n48_O_15_0_2)
  );
  MapT_1 n55 ( // @[Top.scala 403:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .I_2_0_0(n55_I_2_0_0),
    .I_2_0_1(n55_I_2_0_1),
    .I_2_0_2(n55_I_2_0_2),
    .I_3_0_0(n55_I_3_0_0),
    .I_3_0_1(n55_I_3_0_1),
    .I_3_0_2(n55_I_3_0_2),
    .I_4_0_0(n55_I_4_0_0),
    .I_4_0_1(n55_I_4_0_1),
    .I_4_0_2(n55_I_4_0_2),
    .I_5_0_0(n55_I_5_0_0),
    .I_5_0_1(n55_I_5_0_1),
    .I_5_0_2(n55_I_5_0_2),
    .I_6_0_0(n55_I_6_0_0),
    .I_6_0_1(n55_I_6_0_1),
    .I_6_0_2(n55_I_6_0_2),
    .I_7_0_0(n55_I_7_0_0),
    .I_7_0_1(n55_I_7_0_1),
    .I_7_0_2(n55_I_7_0_2),
    .I_8_0_0(n55_I_8_0_0),
    .I_8_0_1(n55_I_8_0_1),
    .I_8_0_2(n55_I_8_0_2),
    .I_9_0_0(n55_I_9_0_0),
    .I_9_0_1(n55_I_9_0_1),
    .I_9_0_2(n55_I_9_0_2),
    .I_10_0_0(n55_I_10_0_0),
    .I_10_0_1(n55_I_10_0_1),
    .I_10_0_2(n55_I_10_0_2),
    .I_11_0_0(n55_I_11_0_0),
    .I_11_0_1(n55_I_11_0_1),
    .I_11_0_2(n55_I_11_0_2),
    .I_12_0_0(n55_I_12_0_0),
    .I_12_0_1(n55_I_12_0_1),
    .I_12_0_2(n55_I_12_0_2),
    .I_13_0_0(n55_I_13_0_0),
    .I_13_0_1(n55_I_13_0_1),
    .I_13_0_2(n55_I_13_0_2),
    .I_14_0_0(n55_I_14_0_0),
    .I_14_0_1(n55_I_14_0_1),
    .I_14_0_2(n55_I_14_0_2),
    .I_15_0_0(n55_I_15_0_0),
    .I_15_0_1(n55_I_15_0_1),
    .I_15_0_2(n55_I_15_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2),
    .O_2_0(n55_O_2_0),
    .O_2_1(n55_O_2_1),
    .O_2_2(n55_O_2_2),
    .O_3_0(n55_O_3_0),
    .O_3_1(n55_O_3_1),
    .O_3_2(n55_O_3_2),
    .O_4_0(n55_O_4_0),
    .O_4_1(n55_O_4_1),
    .O_4_2(n55_O_4_2),
    .O_5_0(n55_O_5_0),
    .O_5_1(n55_O_5_1),
    .O_5_2(n55_O_5_2),
    .O_6_0(n55_O_6_0),
    .O_6_1(n55_O_6_1),
    .O_6_2(n55_O_6_2),
    .O_7_0(n55_O_7_0),
    .O_7_1(n55_O_7_1),
    .O_7_2(n55_O_7_2),
    .O_8_0(n55_O_8_0),
    .O_8_1(n55_O_8_1),
    .O_8_2(n55_O_8_2),
    .O_9_0(n55_O_9_0),
    .O_9_1(n55_O_9_1),
    .O_9_2(n55_O_9_2),
    .O_10_0(n55_O_10_0),
    .O_10_1(n55_O_10_1),
    .O_10_2(n55_O_10_2),
    .O_11_0(n55_O_11_0),
    .O_11_1(n55_O_11_1),
    .O_11_2(n55_O_11_2),
    .O_12_0(n55_O_12_0),
    .O_12_1(n55_O_12_1),
    .O_12_2(n55_O_12_2),
    .O_13_0(n55_O_13_0),
    .O_13_1(n55_O_13_1),
    .O_13_2(n55_O_13_2),
    .O_14_0(n55_O_14_0),
    .O_14_1(n55_O_14_1),
    .O_14_2(n55_O_14_2),
    .O_15_0(n55_O_15_0),
    .O_15_1(n55_O_15_1),
    .O_15_2(n55_O_15_2)
  );
  Map2T_4 n56 ( // @[Top.scala 406:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0(n56_I0_0_0),
    .I0_0_1(n56_I0_0_1),
    .I0_0_2(n56_I0_0_2),
    .I0_1_0(n56_I0_1_0),
    .I0_1_1(n56_I0_1_1),
    .I0_1_2(n56_I0_1_2),
    .I0_2_0(n56_I0_2_0),
    .I0_2_1(n56_I0_2_1),
    .I0_2_2(n56_I0_2_2),
    .I0_3_0(n56_I0_3_0),
    .I0_3_1(n56_I0_3_1),
    .I0_3_2(n56_I0_3_2),
    .I0_4_0(n56_I0_4_0),
    .I0_4_1(n56_I0_4_1),
    .I0_4_2(n56_I0_4_2),
    .I0_5_0(n56_I0_5_0),
    .I0_5_1(n56_I0_5_1),
    .I0_5_2(n56_I0_5_2),
    .I0_6_0(n56_I0_6_0),
    .I0_6_1(n56_I0_6_1),
    .I0_6_2(n56_I0_6_2),
    .I0_7_0(n56_I0_7_0),
    .I0_7_1(n56_I0_7_1),
    .I0_7_2(n56_I0_7_2),
    .I0_8_0(n56_I0_8_0),
    .I0_8_1(n56_I0_8_1),
    .I0_8_2(n56_I0_8_2),
    .I0_9_0(n56_I0_9_0),
    .I0_9_1(n56_I0_9_1),
    .I0_9_2(n56_I0_9_2),
    .I0_10_0(n56_I0_10_0),
    .I0_10_1(n56_I0_10_1),
    .I0_10_2(n56_I0_10_2),
    .I0_11_0(n56_I0_11_0),
    .I0_11_1(n56_I0_11_1),
    .I0_11_2(n56_I0_11_2),
    .I0_12_0(n56_I0_12_0),
    .I0_12_1(n56_I0_12_1),
    .I0_12_2(n56_I0_12_2),
    .I0_13_0(n56_I0_13_0),
    .I0_13_1(n56_I0_13_1),
    .I0_13_2(n56_I0_13_2),
    .I0_14_0(n56_I0_14_0),
    .I0_14_1(n56_I0_14_1),
    .I0_14_2(n56_I0_14_2),
    .I0_15_0(n56_I0_15_0),
    .I0_15_1(n56_I0_15_1),
    .I0_15_2(n56_I0_15_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .I1_2_0(n56_I1_2_0),
    .I1_2_1(n56_I1_2_1),
    .I1_2_2(n56_I1_2_2),
    .I1_3_0(n56_I1_3_0),
    .I1_3_1(n56_I1_3_1),
    .I1_3_2(n56_I1_3_2),
    .I1_4_0(n56_I1_4_0),
    .I1_4_1(n56_I1_4_1),
    .I1_4_2(n56_I1_4_2),
    .I1_5_0(n56_I1_5_0),
    .I1_5_1(n56_I1_5_1),
    .I1_5_2(n56_I1_5_2),
    .I1_6_0(n56_I1_6_0),
    .I1_6_1(n56_I1_6_1),
    .I1_6_2(n56_I1_6_2),
    .I1_7_0(n56_I1_7_0),
    .I1_7_1(n56_I1_7_1),
    .I1_7_2(n56_I1_7_2),
    .I1_8_0(n56_I1_8_0),
    .I1_8_1(n56_I1_8_1),
    .I1_8_2(n56_I1_8_2),
    .I1_9_0(n56_I1_9_0),
    .I1_9_1(n56_I1_9_1),
    .I1_9_2(n56_I1_9_2),
    .I1_10_0(n56_I1_10_0),
    .I1_10_1(n56_I1_10_1),
    .I1_10_2(n56_I1_10_2),
    .I1_11_0(n56_I1_11_0),
    .I1_11_1(n56_I1_11_1),
    .I1_11_2(n56_I1_11_2),
    .I1_12_0(n56_I1_12_0),
    .I1_12_1(n56_I1_12_1),
    .I1_12_2(n56_I1_12_2),
    .I1_13_0(n56_I1_13_0),
    .I1_13_1(n56_I1_13_1),
    .I1_13_2(n56_I1_13_2),
    .I1_14_0(n56_I1_14_0),
    .I1_14_1(n56_I1_14_1),
    .I1_14_2(n56_I1_14_2),
    .I1_15_0(n56_I1_15_0),
    .I1_15_1(n56_I1_15_1),
    .I1_15_2(n56_I1_15_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2),
    .O_2_0_0(n56_O_2_0_0),
    .O_2_0_1(n56_O_2_0_1),
    .O_2_0_2(n56_O_2_0_2),
    .O_2_1_0(n56_O_2_1_0),
    .O_2_1_1(n56_O_2_1_1),
    .O_2_1_2(n56_O_2_1_2),
    .O_3_0_0(n56_O_3_0_0),
    .O_3_0_1(n56_O_3_0_1),
    .O_3_0_2(n56_O_3_0_2),
    .O_3_1_0(n56_O_3_1_0),
    .O_3_1_1(n56_O_3_1_1),
    .O_3_1_2(n56_O_3_1_2),
    .O_4_0_0(n56_O_4_0_0),
    .O_4_0_1(n56_O_4_0_1),
    .O_4_0_2(n56_O_4_0_2),
    .O_4_1_0(n56_O_4_1_0),
    .O_4_1_1(n56_O_4_1_1),
    .O_4_1_2(n56_O_4_1_2),
    .O_5_0_0(n56_O_5_0_0),
    .O_5_0_1(n56_O_5_0_1),
    .O_5_0_2(n56_O_5_0_2),
    .O_5_1_0(n56_O_5_1_0),
    .O_5_1_1(n56_O_5_1_1),
    .O_5_1_2(n56_O_5_1_2),
    .O_6_0_0(n56_O_6_0_0),
    .O_6_0_1(n56_O_6_0_1),
    .O_6_0_2(n56_O_6_0_2),
    .O_6_1_0(n56_O_6_1_0),
    .O_6_1_1(n56_O_6_1_1),
    .O_6_1_2(n56_O_6_1_2),
    .O_7_0_0(n56_O_7_0_0),
    .O_7_0_1(n56_O_7_0_1),
    .O_7_0_2(n56_O_7_0_2),
    .O_7_1_0(n56_O_7_1_0),
    .O_7_1_1(n56_O_7_1_1),
    .O_7_1_2(n56_O_7_1_2),
    .O_8_0_0(n56_O_8_0_0),
    .O_8_0_1(n56_O_8_0_1),
    .O_8_0_2(n56_O_8_0_2),
    .O_8_1_0(n56_O_8_1_0),
    .O_8_1_1(n56_O_8_1_1),
    .O_8_1_2(n56_O_8_1_2),
    .O_9_0_0(n56_O_9_0_0),
    .O_9_0_1(n56_O_9_0_1),
    .O_9_0_2(n56_O_9_0_2),
    .O_9_1_0(n56_O_9_1_0),
    .O_9_1_1(n56_O_9_1_1),
    .O_9_1_2(n56_O_9_1_2),
    .O_10_0_0(n56_O_10_0_0),
    .O_10_0_1(n56_O_10_0_1),
    .O_10_0_2(n56_O_10_0_2),
    .O_10_1_0(n56_O_10_1_0),
    .O_10_1_1(n56_O_10_1_1),
    .O_10_1_2(n56_O_10_1_2),
    .O_11_0_0(n56_O_11_0_0),
    .O_11_0_1(n56_O_11_0_1),
    .O_11_0_2(n56_O_11_0_2),
    .O_11_1_0(n56_O_11_1_0),
    .O_11_1_1(n56_O_11_1_1),
    .O_11_1_2(n56_O_11_1_2),
    .O_12_0_0(n56_O_12_0_0),
    .O_12_0_1(n56_O_12_0_1),
    .O_12_0_2(n56_O_12_0_2),
    .O_12_1_0(n56_O_12_1_0),
    .O_12_1_1(n56_O_12_1_1),
    .O_12_1_2(n56_O_12_1_2),
    .O_13_0_0(n56_O_13_0_0),
    .O_13_0_1(n56_O_13_0_1),
    .O_13_0_2(n56_O_13_0_2),
    .O_13_1_0(n56_O_13_1_0),
    .O_13_1_1(n56_O_13_1_1),
    .O_13_1_2(n56_O_13_1_2),
    .O_14_0_0(n56_O_14_0_0),
    .O_14_0_1(n56_O_14_0_1),
    .O_14_0_2(n56_O_14_0_2),
    .O_14_1_0(n56_O_14_1_0),
    .O_14_1_1(n56_O_14_1_1),
    .O_14_1_2(n56_O_14_1_2),
    .O_15_0_0(n56_O_15_0_0),
    .O_15_0_1(n56_O_15_0_1),
    .O_15_0_2(n56_O_15_0_2),
    .O_15_1_0(n56_O_15_1_0),
    .O_15_1_1(n56_O_15_1_1),
    .O_15_1_2(n56_O_15_1_2)
  );
  ShiftTS_2 n63 ( // @[Top.scala 410:21]
    .clock(n63_clock),
    .valid_up(n63_valid_up),
    .valid_down(n63_valid_down),
    .I_0(n63_I_0),
    .I_1(n63_I_1),
    .I_2(n63_I_2),
    .I_3(n63_I_3),
    .I_4(n63_I_4),
    .I_5(n63_I_5),
    .I_6(n63_I_6),
    .I_7(n63_I_7),
    .I_8(n63_I_8),
    .I_9(n63_I_9),
    .I_10(n63_I_10),
    .I_11(n63_I_11),
    .I_12(n63_I_12),
    .I_13(n63_I_13),
    .I_14(n63_I_14),
    .I_15(n63_I_15),
    .O_0(n63_O_0),
    .O_1(n63_O_1),
    .O_2(n63_O_2),
    .O_3(n63_O_3),
    .O_4(n63_O_4),
    .O_5(n63_O_5),
    .O_6(n63_O_6),
    .O_7(n63_O_7),
    .O_8(n63_O_8),
    .O_9(n63_O_9),
    .O_10(n63_O_10),
    .O_11(n63_O_11),
    .O_12(n63_O_12),
    .O_13(n63_O_13),
    .O_14(n63_O_14),
    .O_15(n63_O_15)
  );
  ShiftTS_2 n64 ( // @[Top.scala 413:21]
    .clock(n64_clock),
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I_0(n64_I_0),
    .I_1(n64_I_1),
    .I_2(n64_I_2),
    .I_3(n64_I_3),
    .I_4(n64_I_4),
    .I_5(n64_I_5),
    .I_6(n64_I_6),
    .I_7(n64_I_7),
    .I_8(n64_I_8),
    .I_9(n64_I_9),
    .I_10(n64_I_10),
    .I_11(n64_I_11),
    .I_12(n64_I_12),
    .I_13(n64_I_13),
    .I_14(n64_I_14),
    .I_15(n64_I_15),
    .O_0(n64_O_0),
    .O_1(n64_O_1),
    .O_2(n64_O_2),
    .O_3(n64_O_3),
    .O_4(n64_O_4),
    .O_5(n64_O_5),
    .O_6(n64_O_6),
    .O_7(n64_O_7),
    .O_8(n64_O_8),
    .O_9(n64_O_9),
    .O_10(n64_O_10),
    .O_11(n64_O_11),
    .O_12(n64_O_12),
    .O_13(n64_O_13),
    .O_14(n64_O_14),
    .O_15(n64_O_15)
  );
  Map2T n65 ( // @[Top.scala 416:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I0_0(n65_I0_0),
    .I0_1(n65_I0_1),
    .I0_2(n65_I0_2),
    .I0_3(n65_I0_3),
    .I0_4(n65_I0_4),
    .I0_5(n65_I0_5),
    .I0_6(n65_I0_6),
    .I0_7(n65_I0_7),
    .I0_8(n65_I0_8),
    .I0_9(n65_I0_9),
    .I0_10(n65_I0_10),
    .I0_11(n65_I0_11),
    .I0_12(n65_I0_12),
    .I0_13(n65_I0_13),
    .I0_14(n65_I0_14),
    .I0_15(n65_I0_15),
    .I1_0(n65_I1_0),
    .I1_1(n65_I1_1),
    .I1_2(n65_I1_2),
    .I1_3(n65_I1_3),
    .I1_4(n65_I1_4),
    .I1_5(n65_I1_5),
    .I1_6(n65_I1_6),
    .I1_7(n65_I1_7),
    .I1_8(n65_I1_8),
    .I1_9(n65_I1_9),
    .I1_10(n65_I1_10),
    .I1_11(n65_I1_11),
    .I1_12(n65_I1_12),
    .I1_13(n65_I1_13),
    .I1_14(n65_I1_14),
    .I1_15(n65_I1_15),
    .O_0_0(n65_O_0_0),
    .O_0_1(n65_O_0_1),
    .O_1_0(n65_O_1_0),
    .O_1_1(n65_O_1_1),
    .O_2_0(n65_O_2_0),
    .O_2_1(n65_O_2_1),
    .O_3_0(n65_O_3_0),
    .O_3_1(n65_O_3_1),
    .O_4_0(n65_O_4_0),
    .O_4_1(n65_O_4_1),
    .O_5_0(n65_O_5_0),
    .O_5_1(n65_O_5_1),
    .O_6_0(n65_O_6_0),
    .O_6_1(n65_O_6_1),
    .O_7_0(n65_O_7_0),
    .O_7_1(n65_O_7_1),
    .O_8_0(n65_O_8_0),
    .O_8_1(n65_O_8_1),
    .O_9_0(n65_O_9_0),
    .O_9_1(n65_O_9_1),
    .O_10_0(n65_O_10_0),
    .O_10_1(n65_O_10_1),
    .O_11_0(n65_O_11_0),
    .O_11_1(n65_O_11_1),
    .O_12_0(n65_O_12_0),
    .O_12_1(n65_O_12_1),
    .O_13_0(n65_O_13_0),
    .O_13_1(n65_O_13_1),
    .O_14_0(n65_O_14_0),
    .O_14_1(n65_O_14_1),
    .O_15_0(n65_O_15_0),
    .O_15_1(n65_O_15_1)
  );
  Map2T_1 n72 ( // @[Top.scala 420:21]
    .valid_up(n72_valid_up),
    .valid_down(n72_valid_down),
    .I0_0_0(n72_I0_0_0),
    .I0_0_1(n72_I0_0_1),
    .I0_1_0(n72_I0_1_0),
    .I0_1_1(n72_I0_1_1),
    .I0_2_0(n72_I0_2_0),
    .I0_2_1(n72_I0_2_1),
    .I0_3_0(n72_I0_3_0),
    .I0_3_1(n72_I0_3_1),
    .I0_4_0(n72_I0_4_0),
    .I0_4_1(n72_I0_4_1),
    .I0_5_0(n72_I0_5_0),
    .I0_5_1(n72_I0_5_1),
    .I0_6_0(n72_I0_6_0),
    .I0_6_1(n72_I0_6_1),
    .I0_7_0(n72_I0_7_0),
    .I0_7_1(n72_I0_7_1),
    .I0_8_0(n72_I0_8_0),
    .I0_8_1(n72_I0_8_1),
    .I0_9_0(n72_I0_9_0),
    .I0_9_1(n72_I0_9_1),
    .I0_10_0(n72_I0_10_0),
    .I0_10_1(n72_I0_10_1),
    .I0_11_0(n72_I0_11_0),
    .I0_11_1(n72_I0_11_1),
    .I0_12_0(n72_I0_12_0),
    .I0_12_1(n72_I0_12_1),
    .I0_13_0(n72_I0_13_0),
    .I0_13_1(n72_I0_13_1),
    .I0_14_0(n72_I0_14_0),
    .I0_14_1(n72_I0_14_1),
    .I0_15_0(n72_I0_15_0),
    .I0_15_1(n72_I0_15_1),
    .I1_0(n72_I1_0),
    .I1_1(n72_I1_1),
    .I1_2(n72_I1_2),
    .I1_3(n72_I1_3),
    .I1_4(n72_I1_4),
    .I1_5(n72_I1_5),
    .I1_6(n72_I1_6),
    .I1_7(n72_I1_7),
    .I1_8(n72_I1_8),
    .I1_9(n72_I1_9),
    .I1_10(n72_I1_10),
    .I1_11(n72_I1_11),
    .I1_12(n72_I1_12),
    .I1_13(n72_I1_13),
    .I1_14(n72_I1_14),
    .I1_15(n72_I1_15),
    .O_0_0(n72_O_0_0),
    .O_0_1(n72_O_0_1),
    .O_0_2(n72_O_0_2),
    .O_1_0(n72_O_1_0),
    .O_1_1(n72_O_1_1),
    .O_1_2(n72_O_1_2),
    .O_2_0(n72_O_2_0),
    .O_2_1(n72_O_2_1),
    .O_2_2(n72_O_2_2),
    .O_3_0(n72_O_3_0),
    .O_3_1(n72_O_3_1),
    .O_3_2(n72_O_3_2),
    .O_4_0(n72_O_4_0),
    .O_4_1(n72_O_4_1),
    .O_4_2(n72_O_4_2),
    .O_5_0(n72_O_5_0),
    .O_5_1(n72_O_5_1),
    .O_5_2(n72_O_5_2),
    .O_6_0(n72_O_6_0),
    .O_6_1(n72_O_6_1),
    .O_6_2(n72_O_6_2),
    .O_7_0(n72_O_7_0),
    .O_7_1(n72_O_7_1),
    .O_7_2(n72_O_7_2),
    .O_8_0(n72_O_8_0),
    .O_8_1(n72_O_8_1),
    .O_8_2(n72_O_8_2),
    .O_9_0(n72_O_9_0),
    .O_9_1(n72_O_9_1),
    .O_9_2(n72_O_9_2),
    .O_10_0(n72_O_10_0),
    .O_10_1(n72_O_10_1),
    .O_10_2(n72_O_10_2),
    .O_11_0(n72_O_11_0),
    .O_11_1(n72_O_11_1),
    .O_11_2(n72_O_11_2),
    .O_12_0(n72_O_12_0),
    .O_12_1(n72_O_12_1),
    .O_12_2(n72_O_12_2),
    .O_13_0(n72_O_13_0),
    .O_13_1(n72_O_13_1),
    .O_13_2(n72_O_13_2),
    .O_14_0(n72_O_14_0),
    .O_14_1(n72_O_14_1),
    .O_14_2(n72_O_14_2),
    .O_15_0(n72_O_15_0),
    .O_15_1(n72_O_15_1),
    .O_15_2(n72_O_15_2)
  );
  MapT n81 ( // @[Top.scala 424:21]
    .valid_up(n81_valid_up),
    .valid_down(n81_valid_down),
    .I_0_0(n81_I_0_0),
    .I_0_1(n81_I_0_1),
    .I_0_2(n81_I_0_2),
    .I_1_0(n81_I_1_0),
    .I_1_1(n81_I_1_1),
    .I_1_2(n81_I_1_2),
    .I_2_0(n81_I_2_0),
    .I_2_1(n81_I_2_1),
    .I_2_2(n81_I_2_2),
    .I_3_0(n81_I_3_0),
    .I_3_1(n81_I_3_1),
    .I_3_2(n81_I_3_2),
    .I_4_0(n81_I_4_0),
    .I_4_1(n81_I_4_1),
    .I_4_2(n81_I_4_2),
    .I_5_0(n81_I_5_0),
    .I_5_1(n81_I_5_1),
    .I_5_2(n81_I_5_2),
    .I_6_0(n81_I_6_0),
    .I_6_1(n81_I_6_1),
    .I_6_2(n81_I_6_2),
    .I_7_0(n81_I_7_0),
    .I_7_1(n81_I_7_1),
    .I_7_2(n81_I_7_2),
    .I_8_0(n81_I_8_0),
    .I_8_1(n81_I_8_1),
    .I_8_2(n81_I_8_2),
    .I_9_0(n81_I_9_0),
    .I_9_1(n81_I_9_1),
    .I_9_2(n81_I_9_2),
    .I_10_0(n81_I_10_0),
    .I_10_1(n81_I_10_1),
    .I_10_2(n81_I_10_2),
    .I_11_0(n81_I_11_0),
    .I_11_1(n81_I_11_1),
    .I_11_2(n81_I_11_2),
    .I_12_0(n81_I_12_0),
    .I_12_1(n81_I_12_1),
    .I_12_2(n81_I_12_2),
    .I_13_0(n81_I_13_0),
    .I_13_1(n81_I_13_1),
    .I_13_2(n81_I_13_2),
    .I_14_0(n81_I_14_0),
    .I_14_1(n81_I_14_1),
    .I_14_2(n81_I_14_2),
    .I_15_0(n81_I_15_0),
    .I_15_1(n81_I_15_1),
    .I_15_2(n81_I_15_2),
    .O_0_0_0(n81_O_0_0_0),
    .O_0_0_1(n81_O_0_0_1),
    .O_0_0_2(n81_O_0_0_2),
    .O_1_0_0(n81_O_1_0_0),
    .O_1_0_1(n81_O_1_0_1),
    .O_1_0_2(n81_O_1_0_2),
    .O_2_0_0(n81_O_2_0_0),
    .O_2_0_1(n81_O_2_0_1),
    .O_2_0_2(n81_O_2_0_2),
    .O_3_0_0(n81_O_3_0_0),
    .O_3_0_1(n81_O_3_0_1),
    .O_3_0_2(n81_O_3_0_2),
    .O_4_0_0(n81_O_4_0_0),
    .O_4_0_1(n81_O_4_0_1),
    .O_4_0_2(n81_O_4_0_2),
    .O_5_0_0(n81_O_5_0_0),
    .O_5_0_1(n81_O_5_0_1),
    .O_5_0_2(n81_O_5_0_2),
    .O_6_0_0(n81_O_6_0_0),
    .O_6_0_1(n81_O_6_0_1),
    .O_6_0_2(n81_O_6_0_2),
    .O_7_0_0(n81_O_7_0_0),
    .O_7_0_1(n81_O_7_0_1),
    .O_7_0_2(n81_O_7_0_2),
    .O_8_0_0(n81_O_8_0_0),
    .O_8_0_1(n81_O_8_0_1),
    .O_8_0_2(n81_O_8_0_2),
    .O_9_0_0(n81_O_9_0_0),
    .O_9_0_1(n81_O_9_0_1),
    .O_9_0_2(n81_O_9_0_2),
    .O_10_0_0(n81_O_10_0_0),
    .O_10_0_1(n81_O_10_0_1),
    .O_10_0_2(n81_O_10_0_2),
    .O_11_0_0(n81_O_11_0_0),
    .O_11_0_1(n81_O_11_0_1),
    .O_11_0_2(n81_O_11_0_2),
    .O_12_0_0(n81_O_12_0_0),
    .O_12_0_1(n81_O_12_0_1),
    .O_12_0_2(n81_O_12_0_2),
    .O_13_0_0(n81_O_13_0_0),
    .O_13_0_1(n81_O_13_0_1),
    .O_13_0_2(n81_O_13_0_2),
    .O_14_0_0(n81_O_14_0_0),
    .O_14_0_1(n81_O_14_0_1),
    .O_14_0_2(n81_O_14_0_2),
    .O_15_0_0(n81_O_15_0_0),
    .O_15_0_1(n81_O_15_0_1),
    .O_15_0_2(n81_O_15_0_2)
  );
  MapT_1 n88 ( // @[Top.scala 427:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_0_0_1(n88_I_0_0_1),
    .I_0_0_2(n88_I_0_0_2),
    .I_1_0_0(n88_I_1_0_0),
    .I_1_0_1(n88_I_1_0_1),
    .I_1_0_2(n88_I_1_0_2),
    .I_2_0_0(n88_I_2_0_0),
    .I_2_0_1(n88_I_2_0_1),
    .I_2_0_2(n88_I_2_0_2),
    .I_3_0_0(n88_I_3_0_0),
    .I_3_0_1(n88_I_3_0_1),
    .I_3_0_2(n88_I_3_0_2),
    .I_4_0_0(n88_I_4_0_0),
    .I_4_0_1(n88_I_4_0_1),
    .I_4_0_2(n88_I_4_0_2),
    .I_5_0_0(n88_I_5_0_0),
    .I_5_0_1(n88_I_5_0_1),
    .I_5_0_2(n88_I_5_0_2),
    .I_6_0_0(n88_I_6_0_0),
    .I_6_0_1(n88_I_6_0_1),
    .I_6_0_2(n88_I_6_0_2),
    .I_7_0_0(n88_I_7_0_0),
    .I_7_0_1(n88_I_7_0_1),
    .I_7_0_2(n88_I_7_0_2),
    .I_8_0_0(n88_I_8_0_0),
    .I_8_0_1(n88_I_8_0_1),
    .I_8_0_2(n88_I_8_0_2),
    .I_9_0_0(n88_I_9_0_0),
    .I_9_0_1(n88_I_9_0_1),
    .I_9_0_2(n88_I_9_0_2),
    .I_10_0_0(n88_I_10_0_0),
    .I_10_0_1(n88_I_10_0_1),
    .I_10_0_2(n88_I_10_0_2),
    .I_11_0_0(n88_I_11_0_0),
    .I_11_0_1(n88_I_11_0_1),
    .I_11_0_2(n88_I_11_0_2),
    .I_12_0_0(n88_I_12_0_0),
    .I_12_0_1(n88_I_12_0_1),
    .I_12_0_2(n88_I_12_0_2),
    .I_13_0_0(n88_I_13_0_0),
    .I_13_0_1(n88_I_13_0_1),
    .I_13_0_2(n88_I_13_0_2),
    .I_14_0_0(n88_I_14_0_0),
    .I_14_0_1(n88_I_14_0_1),
    .I_14_0_2(n88_I_14_0_2),
    .I_15_0_0(n88_I_15_0_0),
    .I_15_0_1(n88_I_15_0_1),
    .I_15_0_2(n88_I_15_0_2),
    .O_0_0(n88_O_0_0),
    .O_0_1(n88_O_0_1),
    .O_0_2(n88_O_0_2),
    .O_1_0(n88_O_1_0),
    .O_1_1(n88_O_1_1),
    .O_1_2(n88_O_1_2),
    .O_2_0(n88_O_2_0),
    .O_2_1(n88_O_2_1),
    .O_2_2(n88_O_2_2),
    .O_3_0(n88_O_3_0),
    .O_3_1(n88_O_3_1),
    .O_3_2(n88_O_3_2),
    .O_4_0(n88_O_4_0),
    .O_4_1(n88_O_4_1),
    .O_4_2(n88_O_4_2),
    .O_5_0(n88_O_5_0),
    .O_5_1(n88_O_5_1),
    .O_5_2(n88_O_5_2),
    .O_6_0(n88_O_6_0),
    .O_6_1(n88_O_6_1),
    .O_6_2(n88_O_6_2),
    .O_7_0(n88_O_7_0),
    .O_7_1(n88_O_7_1),
    .O_7_2(n88_O_7_2),
    .O_8_0(n88_O_8_0),
    .O_8_1(n88_O_8_1),
    .O_8_2(n88_O_8_2),
    .O_9_0(n88_O_9_0),
    .O_9_1(n88_O_9_1),
    .O_9_2(n88_O_9_2),
    .O_10_0(n88_O_10_0),
    .O_10_1(n88_O_10_1),
    .O_10_2(n88_O_10_2),
    .O_11_0(n88_O_11_0),
    .O_11_1(n88_O_11_1),
    .O_11_2(n88_O_11_2),
    .O_12_0(n88_O_12_0),
    .O_12_1(n88_O_12_1),
    .O_12_2(n88_O_12_2),
    .O_13_0(n88_O_13_0),
    .O_13_1(n88_O_13_1),
    .O_13_2(n88_O_13_2),
    .O_14_0(n88_O_14_0),
    .O_14_1(n88_O_14_1),
    .O_14_2(n88_O_14_2),
    .O_15_0(n88_O_15_0),
    .O_15_1(n88_O_15_1),
    .O_15_2(n88_O_15_2)
  );
  Map2T_7 n89 ( // @[Top.scala 430:21]
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I0_0_0_0(n89_I0_0_0_0),
    .I0_0_0_1(n89_I0_0_0_1),
    .I0_0_0_2(n89_I0_0_0_2),
    .I0_0_1_0(n89_I0_0_1_0),
    .I0_0_1_1(n89_I0_0_1_1),
    .I0_0_1_2(n89_I0_0_1_2),
    .I0_1_0_0(n89_I0_1_0_0),
    .I0_1_0_1(n89_I0_1_0_1),
    .I0_1_0_2(n89_I0_1_0_2),
    .I0_1_1_0(n89_I0_1_1_0),
    .I0_1_1_1(n89_I0_1_1_1),
    .I0_1_1_2(n89_I0_1_1_2),
    .I0_2_0_0(n89_I0_2_0_0),
    .I0_2_0_1(n89_I0_2_0_1),
    .I0_2_0_2(n89_I0_2_0_2),
    .I0_2_1_0(n89_I0_2_1_0),
    .I0_2_1_1(n89_I0_2_1_1),
    .I0_2_1_2(n89_I0_2_1_2),
    .I0_3_0_0(n89_I0_3_0_0),
    .I0_3_0_1(n89_I0_3_0_1),
    .I0_3_0_2(n89_I0_3_0_2),
    .I0_3_1_0(n89_I0_3_1_0),
    .I0_3_1_1(n89_I0_3_1_1),
    .I0_3_1_2(n89_I0_3_1_2),
    .I0_4_0_0(n89_I0_4_0_0),
    .I0_4_0_1(n89_I0_4_0_1),
    .I0_4_0_2(n89_I0_4_0_2),
    .I0_4_1_0(n89_I0_4_1_0),
    .I0_4_1_1(n89_I0_4_1_1),
    .I0_4_1_2(n89_I0_4_1_2),
    .I0_5_0_0(n89_I0_5_0_0),
    .I0_5_0_1(n89_I0_5_0_1),
    .I0_5_0_2(n89_I0_5_0_2),
    .I0_5_1_0(n89_I0_5_1_0),
    .I0_5_1_1(n89_I0_5_1_1),
    .I0_5_1_2(n89_I0_5_1_2),
    .I0_6_0_0(n89_I0_6_0_0),
    .I0_6_0_1(n89_I0_6_0_1),
    .I0_6_0_2(n89_I0_6_0_2),
    .I0_6_1_0(n89_I0_6_1_0),
    .I0_6_1_1(n89_I0_6_1_1),
    .I0_6_1_2(n89_I0_6_1_2),
    .I0_7_0_0(n89_I0_7_0_0),
    .I0_7_0_1(n89_I0_7_0_1),
    .I0_7_0_2(n89_I0_7_0_2),
    .I0_7_1_0(n89_I0_7_1_0),
    .I0_7_1_1(n89_I0_7_1_1),
    .I0_7_1_2(n89_I0_7_1_2),
    .I0_8_0_0(n89_I0_8_0_0),
    .I0_8_0_1(n89_I0_8_0_1),
    .I0_8_0_2(n89_I0_8_0_2),
    .I0_8_1_0(n89_I0_8_1_0),
    .I0_8_1_1(n89_I0_8_1_1),
    .I0_8_1_2(n89_I0_8_1_2),
    .I0_9_0_0(n89_I0_9_0_0),
    .I0_9_0_1(n89_I0_9_0_1),
    .I0_9_0_2(n89_I0_9_0_2),
    .I0_9_1_0(n89_I0_9_1_0),
    .I0_9_1_1(n89_I0_9_1_1),
    .I0_9_1_2(n89_I0_9_1_2),
    .I0_10_0_0(n89_I0_10_0_0),
    .I0_10_0_1(n89_I0_10_0_1),
    .I0_10_0_2(n89_I0_10_0_2),
    .I0_10_1_0(n89_I0_10_1_0),
    .I0_10_1_1(n89_I0_10_1_1),
    .I0_10_1_2(n89_I0_10_1_2),
    .I0_11_0_0(n89_I0_11_0_0),
    .I0_11_0_1(n89_I0_11_0_1),
    .I0_11_0_2(n89_I0_11_0_2),
    .I0_11_1_0(n89_I0_11_1_0),
    .I0_11_1_1(n89_I0_11_1_1),
    .I0_11_1_2(n89_I0_11_1_2),
    .I0_12_0_0(n89_I0_12_0_0),
    .I0_12_0_1(n89_I0_12_0_1),
    .I0_12_0_2(n89_I0_12_0_2),
    .I0_12_1_0(n89_I0_12_1_0),
    .I0_12_1_1(n89_I0_12_1_1),
    .I0_12_1_2(n89_I0_12_1_2),
    .I0_13_0_0(n89_I0_13_0_0),
    .I0_13_0_1(n89_I0_13_0_1),
    .I0_13_0_2(n89_I0_13_0_2),
    .I0_13_1_0(n89_I0_13_1_0),
    .I0_13_1_1(n89_I0_13_1_1),
    .I0_13_1_2(n89_I0_13_1_2),
    .I0_14_0_0(n89_I0_14_0_0),
    .I0_14_0_1(n89_I0_14_0_1),
    .I0_14_0_2(n89_I0_14_0_2),
    .I0_14_1_0(n89_I0_14_1_0),
    .I0_14_1_1(n89_I0_14_1_1),
    .I0_14_1_2(n89_I0_14_1_2),
    .I0_15_0_0(n89_I0_15_0_0),
    .I0_15_0_1(n89_I0_15_0_1),
    .I0_15_0_2(n89_I0_15_0_2),
    .I0_15_1_0(n89_I0_15_1_0),
    .I0_15_1_1(n89_I0_15_1_1),
    .I0_15_1_2(n89_I0_15_1_2),
    .I1_0_0(n89_I1_0_0),
    .I1_0_1(n89_I1_0_1),
    .I1_0_2(n89_I1_0_2),
    .I1_1_0(n89_I1_1_0),
    .I1_1_1(n89_I1_1_1),
    .I1_1_2(n89_I1_1_2),
    .I1_2_0(n89_I1_2_0),
    .I1_2_1(n89_I1_2_1),
    .I1_2_2(n89_I1_2_2),
    .I1_3_0(n89_I1_3_0),
    .I1_3_1(n89_I1_3_1),
    .I1_3_2(n89_I1_3_2),
    .I1_4_0(n89_I1_4_0),
    .I1_4_1(n89_I1_4_1),
    .I1_4_2(n89_I1_4_2),
    .I1_5_0(n89_I1_5_0),
    .I1_5_1(n89_I1_5_1),
    .I1_5_2(n89_I1_5_2),
    .I1_6_0(n89_I1_6_0),
    .I1_6_1(n89_I1_6_1),
    .I1_6_2(n89_I1_6_2),
    .I1_7_0(n89_I1_7_0),
    .I1_7_1(n89_I1_7_1),
    .I1_7_2(n89_I1_7_2),
    .I1_8_0(n89_I1_8_0),
    .I1_8_1(n89_I1_8_1),
    .I1_8_2(n89_I1_8_2),
    .I1_9_0(n89_I1_9_0),
    .I1_9_1(n89_I1_9_1),
    .I1_9_2(n89_I1_9_2),
    .I1_10_0(n89_I1_10_0),
    .I1_10_1(n89_I1_10_1),
    .I1_10_2(n89_I1_10_2),
    .I1_11_0(n89_I1_11_0),
    .I1_11_1(n89_I1_11_1),
    .I1_11_2(n89_I1_11_2),
    .I1_12_0(n89_I1_12_0),
    .I1_12_1(n89_I1_12_1),
    .I1_12_2(n89_I1_12_2),
    .I1_13_0(n89_I1_13_0),
    .I1_13_1(n89_I1_13_1),
    .I1_13_2(n89_I1_13_2),
    .I1_14_0(n89_I1_14_0),
    .I1_14_1(n89_I1_14_1),
    .I1_14_2(n89_I1_14_2),
    .I1_15_0(n89_I1_15_0),
    .I1_15_1(n89_I1_15_1),
    .I1_15_2(n89_I1_15_2),
    .O_0_0_0(n89_O_0_0_0),
    .O_0_0_1(n89_O_0_0_1),
    .O_0_0_2(n89_O_0_0_2),
    .O_0_1_0(n89_O_0_1_0),
    .O_0_1_1(n89_O_0_1_1),
    .O_0_1_2(n89_O_0_1_2),
    .O_0_2_0(n89_O_0_2_0),
    .O_0_2_1(n89_O_0_2_1),
    .O_0_2_2(n89_O_0_2_2),
    .O_1_0_0(n89_O_1_0_0),
    .O_1_0_1(n89_O_1_0_1),
    .O_1_0_2(n89_O_1_0_2),
    .O_1_1_0(n89_O_1_1_0),
    .O_1_1_1(n89_O_1_1_1),
    .O_1_1_2(n89_O_1_1_2),
    .O_1_2_0(n89_O_1_2_0),
    .O_1_2_1(n89_O_1_2_1),
    .O_1_2_2(n89_O_1_2_2),
    .O_2_0_0(n89_O_2_0_0),
    .O_2_0_1(n89_O_2_0_1),
    .O_2_0_2(n89_O_2_0_2),
    .O_2_1_0(n89_O_2_1_0),
    .O_2_1_1(n89_O_2_1_1),
    .O_2_1_2(n89_O_2_1_2),
    .O_2_2_0(n89_O_2_2_0),
    .O_2_2_1(n89_O_2_2_1),
    .O_2_2_2(n89_O_2_2_2),
    .O_3_0_0(n89_O_3_0_0),
    .O_3_0_1(n89_O_3_0_1),
    .O_3_0_2(n89_O_3_0_2),
    .O_3_1_0(n89_O_3_1_0),
    .O_3_1_1(n89_O_3_1_1),
    .O_3_1_2(n89_O_3_1_2),
    .O_3_2_0(n89_O_3_2_0),
    .O_3_2_1(n89_O_3_2_1),
    .O_3_2_2(n89_O_3_2_2),
    .O_4_0_0(n89_O_4_0_0),
    .O_4_0_1(n89_O_4_0_1),
    .O_4_0_2(n89_O_4_0_2),
    .O_4_1_0(n89_O_4_1_0),
    .O_4_1_1(n89_O_4_1_1),
    .O_4_1_2(n89_O_4_1_2),
    .O_4_2_0(n89_O_4_2_0),
    .O_4_2_1(n89_O_4_2_1),
    .O_4_2_2(n89_O_4_2_2),
    .O_5_0_0(n89_O_5_0_0),
    .O_5_0_1(n89_O_5_0_1),
    .O_5_0_2(n89_O_5_0_2),
    .O_5_1_0(n89_O_5_1_0),
    .O_5_1_1(n89_O_5_1_1),
    .O_5_1_2(n89_O_5_1_2),
    .O_5_2_0(n89_O_5_2_0),
    .O_5_2_1(n89_O_5_2_1),
    .O_5_2_2(n89_O_5_2_2),
    .O_6_0_0(n89_O_6_0_0),
    .O_6_0_1(n89_O_6_0_1),
    .O_6_0_2(n89_O_6_0_2),
    .O_6_1_0(n89_O_6_1_0),
    .O_6_1_1(n89_O_6_1_1),
    .O_6_1_2(n89_O_6_1_2),
    .O_6_2_0(n89_O_6_2_0),
    .O_6_2_1(n89_O_6_2_1),
    .O_6_2_2(n89_O_6_2_2),
    .O_7_0_0(n89_O_7_0_0),
    .O_7_0_1(n89_O_7_0_1),
    .O_7_0_2(n89_O_7_0_2),
    .O_7_1_0(n89_O_7_1_0),
    .O_7_1_1(n89_O_7_1_1),
    .O_7_1_2(n89_O_7_1_2),
    .O_7_2_0(n89_O_7_2_0),
    .O_7_2_1(n89_O_7_2_1),
    .O_7_2_2(n89_O_7_2_2),
    .O_8_0_0(n89_O_8_0_0),
    .O_8_0_1(n89_O_8_0_1),
    .O_8_0_2(n89_O_8_0_2),
    .O_8_1_0(n89_O_8_1_0),
    .O_8_1_1(n89_O_8_1_1),
    .O_8_1_2(n89_O_8_1_2),
    .O_8_2_0(n89_O_8_2_0),
    .O_8_2_1(n89_O_8_2_1),
    .O_8_2_2(n89_O_8_2_2),
    .O_9_0_0(n89_O_9_0_0),
    .O_9_0_1(n89_O_9_0_1),
    .O_9_0_2(n89_O_9_0_2),
    .O_9_1_0(n89_O_9_1_0),
    .O_9_1_1(n89_O_9_1_1),
    .O_9_1_2(n89_O_9_1_2),
    .O_9_2_0(n89_O_9_2_0),
    .O_9_2_1(n89_O_9_2_1),
    .O_9_2_2(n89_O_9_2_2),
    .O_10_0_0(n89_O_10_0_0),
    .O_10_0_1(n89_O_10_0_1),
    .O_10_0_2(n89_O_10_0_2),
    .O_10_1_0(n89_O_10_1_0),
    .O_10_1_1(n89_O_10_1_1),
    .O_10_1_2(n89_O_10_1_2),
    .O_10_2_0(n89_O_10_2_0),
    .O_10_2_1(n89_O_10_2_1),
    .O_10_2_2(n89_O_10_2_2),
    .O_11_0_0(n89_O_11_0_0),
    .O_11_0_1(n89_O_11_0_1),
    .O_11_0_2(n89_O_11_0_2),
    .O_11_1_0(n89_O_11_1_0),
    .O_11_1_1(n89_O_11_1_1),
    .O_11_1_2(n89_O_11_1_2),
    .O_11_2_0(n89_O_11_2_0),
    .O_11_2_1(n89_O_11_2_1),
    .O_11_2_2(n89_O_11_2_2),
    .O_12_0_0(n89_O_12_0_0),
    .O_12_0_1(n89_O_12_0_1),
    .O_12_0_2(n89_O_12_0_2),
    .O_12_1_0(n89_O_12_1_0),
    .O_12_1_1(n89_O_12_1_1),
    .O_12_1_2(n89_O_12_1_2),
    .O_12_2_0(n89_O_12_2_0),
    .O_12_2_1(n89_O_12_2_1),
    .O_12_2_2(n89_O_12_2_2),
    .O_13_0_0(n89_O_13_0_0),
    .O_13_0_1(n89_O_13_0_1),
    .O_13_0_2(n89_O_13_0_2),
    .O_13_1_0(n89_O_13_1_0),
    .O_13_1_1(n89_O_13_1_1),
    .O_13_1_2(n89_O_13_1_2),
    .O_13_2_0(n89_O_13_2_0),
    .O_13_2_1(n89_O_13_2_1),
    .O_13_2_2(n89_O_13_2_2),
    .O_14_0_0(n89_O_14_0_0),
    .O_14_0_1(n89_O_14_0_1),
    .O_14_0_2(n89_O_14_0_2),
    .O_14_1_0(n89_O_14_1_0),
    .O_14_1_1(n89_O_14_1_1),
    .O_14_1_2(n89_O_14_1_2),
    .O_14_2_0(n89_O_14_2_0),
    .O_14_2_1(n89_O_14_2_1),
    .O_14_2_2(n89_O_14_2_2),
    .O_15_0_0(n89_O_15_0_0),
    .O_15_0_1(n89_O_15_0_1),
    .O_15_0_2(n89_O_15_0_2),
    .O_15_1_0(n89_O_15_1_0),
    .O_15_1_1(n89_O_15_1_1),
    .O_15_1_2(n89_O_15_1_2),
    .O_15_2_0(n89_O_15_2_0),
    .O_15_2_1(n89_O_15_2_1),
    .O_15_2_2(n89_O_15_2_2)
  );
  MapT_6 n98 ( // @[Top.scala 434:21]
    .valid_up(n98_valid_up),
    .valid_down(n98_valid_down),
    .I_0_0_0(n98_I_0_0_0),
    .I_0_0_1(n98_I_0_0_1),
    .I_0_0_2(n98_I_0_0_2),
    .I_0_1_0(n98_I_0_1_0),
    .I_0_1_1(n98_I_0_1_1),
    .I_0_1_2(n98_I_0_1_2),
    .I_0_2_0(n98_I_0_2_0),
    .I_0_2_1(n98_I_0_2_1),
    .I_0_2_2(n98_I_0_2_2),
    .I_1_0_0(n98_I_1_0_0),
    .I_1_0_1(n98_I_1_0_1),
    .I_1_0_2(n98_I_1_0_2),
    .I_1_1_0(n98_I_1_1_0),
    .I_1_1_1(n98_I_1_1_1),
    .I_1_1_2(n98_I_1_1_2),
    .I_1_2_0(n98_I_1_2_0),
    .I_1_2_1(n98_I_1_2_1),
    .I_1_2_2(n98_I_1_2_2),
    .I_2_0_0(n98_I_2_0_0),
    .I_2_0_1(n98_I_2_0_1),
    .I_2_0_2(n98_I_2_0_2),
    .I_2_1_0(n98_I_2_1_0),
    .I_2_1_1(n98_I_2_1_1),
    .I_2_1_2(n98_I_2_1_2),
    .I_2_2_0(n98_I_2_2_0),
    .I_2_2_1(n98_I_2_2_1),
    .I_2_2_2(n98_I_2_2_2),
    .I_3_0_0(n98_I_3_0_0),
    .I_3_0_1(n98_I_3_0_1),
    .I_3_0_2(n98_I_3_0_2),
    .I_3_1_0(n98_I_3_1_0),
    .I_3_1_1(n98_I_3_1_1),
    .I_3_1_2(n98_I_3_1_2),
    .I_3_2_0(n98_I_3_2_0),
    .I_3_2_1(n98_I_3_2_1),
    .I_3_2_2(n98_I_3_2_2),
    .I_4_0_0(n98_I_4_0_0),
    .I_4_0_1(n98_I_4_0_1),
    .I_4_0_2(n98_I_4_0_2),
    .I_4_1_0(n98_I_4_1_0),
    .I_4_1_1(n98_I_4_1_1),
    .I_4_1_2(n98_I_4_1_2),
    .I_4_2_0(n98_I_4_2_0),
    .I_4_2_1(n98_I_4_2_1),
    .I_4_2_2(n98_I_4_2_2),
    .I_5_0_0(n98_I_5_0_0),
    .I_5_0_1(n98_I_5_0_1),
    .I_5_0_2(n98_I_5_0_2),
    .I_5_1_0(n98_I_5_1_0),
    .I_5_1_1(n98_I_5_1_1),
    .I_5_1_2(n98_I_5_1_2),
    .I_5_2_0(n98_I_5_2_0),
    .I_5_2_1(n98_I_5_2_1),
    .I_5_2_2(n98_I_5_2_2),
    .I_6_0_0(n98_I_6_0_0),
    .I_6_0_1(n98_I_6_0_1),
    .I_6_0_2(n98_I_6_0_2),
    .I_6_1_0(n98_I_6_1_0),
    .I_6_1_1(n98_I_6_1_1),
    .I_6_1_2(n98_I_6_1_2),
    .I_6_2_0(n98_I_6_2_0),
    .I_6_2_1(n98_I_6_2_1),
    .I_6_2_2(n98_I_6_2_2),
    .I_7_0_0(n98_I_7_0_0),
    .I_7_0_1(n98_I_7_0_1),
    .I_7_0_2(n98_I_7_0_2),
    .I_7_1_0(n98_I_7_1_0),
    .I_7_1_1(n98_I_7_1_1),
    .I_7_1_2(n98_I_7_1_2),
    .I_7_2_0(n98_I_7_2_0),
    .I_7_2_1(n98_I_7_2_1),
    .I_7_2_2(n98_I_7_2_2),
    .I_8_0_0(n98_I_8_0_0),
    .I_8_0_1(n98_I_8_0_1),
    .I_8_0_2(n98_I_8_0_2),
    .I_8_1_0(n98_I_8_1_0),
    .I_8_1_1(n98_I_8_1_1),
    .I_8_1_2(n98_I_8_1_2),
    .I_8_2_0(n98_I_8_2_0),
    .I_8_2_1(n98_I_8_2_1),
    .I_8_2_2(n98_I_8_2_2),
    .I_9_0_0(n98_I_9_0_0),
    .I_9_0_1(n98_I_9_0_1),
    .I_9_0_2(n98_I_9_0_2),
    .I_9_1_0(n98_I_9_1_0),
    .I_9_1_1(n98_I_9_1_1),
    .I_9_1_2(n98_I_9_1_2),
    .I_9_2_0(n98_I_9_2_0),
    .I_9_2_1(n98_I_9_2_1),
    .I_9_2_2(n98_I_9_2_2),
    .I_10_0_0(n98_I_10_0_0),
    .I_10_0_1(n98_I_10_0_1),
    .I_10_0_2(n98_I_10_0_2),
    .I_10_1_0(n98_I_10_1_0),
    .I_10_1_1(n98_I_10_1_1),
    .I_10_1_2(n98_I_10_1_2),
    .I_10_2_0(n98_I_10_2_0),
    .I_10_2_1(n98_I_10_2_1),
    .I_10_2_2(n98_I_10_2_2),
    .I_11_0_0(n98_I_11_0_0),
    .I_11_0_1(n98_I_11_0_1),
    .I_11_0_2(n98_I_11_0_2),
    .I_11_1_0(n98_I_11_1_0),
    .I_11_1_1(n98_I_11_1_1),
    .I_11_1_2(n98_I_11_1_2),
    .I_11_2_0(n98_I_11_2_0),
    .I_11_2_1(n98_I_11_2_1),
    .I_11_2_2(n98_I_11_2_2),
    .I_12_0_0(n98_I_12_0_0),
    .I_12_0_1(n98_I_12_0_1),
    .I_12_0_2(n98_I_12_0_2),
    .I_12_1_0(n98_I_12_1_0),
    .I_12_1_1(n98_I_12_1_1),
    .I_12_1_2(n98_I_12_1_2),
    .I_12_2_0(n98_I_12_2_0),
    .I_12_2_1(n98_I_12_2_1),
    .I_12_2_2(n98_I_12_2_2),
    .I_13_0_0(n98_I_13_0_0),
    .I_13_0_1(n98_I_13_0_1),
    .I_13_0_2(n98_I_13_0_2),
    .I_13_1_0(n98_I_13_1_0),
    .I_13_1_1(n98_I_13_1_1),
    .I_13_1_2(n98_I_13_1_2),
    .I_13_2_0(n98_I_13_2_0),
    .I_13_2_1(n98_I_13_2_1),
    .I_13_2_2(n98_I_13_2_2),
    .I_14_0_0(n98_I_14_0_0),
    .I_14_0_1(n98_I_14_0_1),
    .I_14_0_2(n98_I_14_0_2),
    .I_14_1_0(n98_I_14_1_0),
    .I_14_1_1(n98_I_14_1_1),
    .I_14_1_2(n98_I_14_1_2),
    .I_14_2_0(n98_I_14_2_0),
    .I_14_2_1(n98_I_14_2_1),
    .I_14_2_2(n98_I_14_2_2),
    .I_15_0_0(n98_I_15_0_0),
    .I_15_0_1(n98_I_15_0_1),
    .I_15_0_2(n98_I_15_0_2),
    .I_15_1_0(n98_I_15_1_0),
    .I_15_1_1(n98_I_15_1_1),
    .I_15_1_2(n98_I_15_1_2),
    .I_15_2_0(n98_I_15_2_0),
    .I_15_2_1(n98_I_15_2_1),
    .I_15_2_2(n98_I_15_2_2),
    .O_0_0_0_0(n98_O_0_0_0_0),
    .O_0_0_0_1(n98_O_0_0_0_1),
    .O_0_0_0_2(n98_O_0_0_0_2),
    .O_0_0_1_0(n98_O_0_0_1_0),
    .O_0_0_1_1(n98_O_0_0_1_1),
    .O_0_0_1_2(n98_O_0_0_1_2),
    .O_0_0_2_0(n98_O_0_0_2_0),
    .O_0_0_2_1(n98_O_0_0_2_1),
    .O_0_0_2_2(n98_O_0_0_2_2),
    .O_1_0_0_0(n98_O_1_0_0_0),
    .O_1_0_0_1(n98_O_1_0_0_1),
    .O_1_0_0_2(n98_O_1_0_0_2),
    .O_1_0_1_0(n98_O_1_0_1_0),
    .O_1_0_1_1(n98_O_1_0_1_1),
    .O_1_0_1_2(n98_O_1_0_1_2),
    .O_1_0_2_0(n98_O_1_0_2_0),
    .O_1_0_2_1(n98_O_1_0_2_1),
    .O_1_0_2_2(n98_O_1_0_2_2),
    .O_2_0_0_0(n98_O_2_0_0_0),
    .O_2_0_0_1(n98_O_2_0_0_1),
    .O_2_0_0_2(n98_O_2_0_0_2),
    .O_2_0_1_0(n98_O_2_0_1_0),
    .O_2_0_1_1(n98_O_2_0_1_1),
    .O_2_0_1_2(n98_O_2_0_1_2),
    .O_2_0_2_0(n98_O_2_0_2_0),
    .O_2_0_2_1(n98_O_2_0_2_1),
    .O_2_0_2_2(n98_O_2_0_2_2),
    .O_3_0_0_0(n98_O_3_0_0_0),
    .O_3_0_0_1(n98_O_3_0_0_1),
    .O_3_0_0_2(n98_O_3_0_0_2),
    .O_3_0_1_0(n98_O_3_0_1_0),
    .O_3_0_1_1(n98_O_3_0_1_1),
    .O_3_0_1_2(n98_O_3_0_1_2),
    .O_3_0_2_0(n98_O_3_0_2_0),
    .O_3_0_2_1(n98_O_3_0_2_1),
    .O_3_0_2_2(n98_O_3_0_2_2),
    .O_4_0_0_0(n98_O_4_0_0_0),
    .O_4_0_0_1(n98_O_4_0_0_1),
    .O_4_0_0_2(n98_O_4_0_0_2),
    .O_4_0_1_0(n98_O_4_0_1_0),
    .O_4_0_1_1(n98_O_4_0_1_1),
    .O_4_0_1_2(n98_O_4_0_1_2),
    .O_4_0_2_0(n98_O_4_0_2_0),
    .O_4_0_2_1(n98_O_4_0_2_1),
    .O_4_0_2_2(n98_O_4_0_2_2),
    .O_5_0_0_0(n98_O_5_0_0_0),
    .O_5_0_0_1(n98_O_5_0_0_1),
    .O_5_0_0_2(n98_O_5_0_0_2),
    .O_5_0_1_0(n98_O_5_0_1_0),
    .O_5_0_1_1(n98_O_5_0_1_1),
    .O_5_0_1_2(n98_O_5_0_1_2),
    .O_5_0_2_0(n98_O_5_0_2_0),
    .O_5_0_2_1(n98_O_5_0_2_1),
    .O_5_0_2_2(n98_O_5_0_2_2),
    .O_6_0_0_0(n98_O_6_0_0_0),
    .O_6_0_0_1(n98_O_6_0_0_1),
    .O_6_0_0_2(n98_O_6_0_0_2),
    .O_6_0_1_0(n98_O_6_0_1_0),
    .O_6_0_1_1(n98_O_6_0_1_1),
    .O_6_0_1_2(n98_O_6_0_1_2),
    .O_6_0_2_0(n98_O_6_0_2_0),
    .O_6_0_2_1(n98_O_6_0_2_1),
    .O_6_0_2_2(n98_O_6_0_2_2),
    .O_7_0_0_0(n98_O_7_0_0_0),
    .O_7_0_0_1(n98_O_7_0_0_1),
    .O_7_0_0_2(n98_O_7_0_0_2),
    .O_7_0_1_0(n98_O_7_0_1_0),
    .O_7_0_1_1(n98_O_7_0_1_1),
    .O_7_0_1_2(n98_O_7_0_1_2),
    .O_7_0_2_0(n98_O_7_0_2_0),
    .O_7_0_2_1(n98_O_7_0_2_1),
    .O_7_0_2_2(n98_O_7_0_2_2),
    .O_8_0_0_0(n98_O_8_0_0_0),
    .O_8_0_0_1(n98_O_8_0_0_1),
    .O_8_0_0_2(n98_O_8_0_0_2),
    .O_8_0_1_0(n98_O_8_0_1_0),
    .O_8_0_1_1(n98_O_8_0_1_1),
    .O_8_0_1_2(n98_O_8_0_1_2),
    .O_8_0_2_0(n98_O_8_0_2_0),
    .O_8_0_2_1(n98_O_8_0_2_1),
    .O_8_0_2_2(n98_O_8_0_2_2),
    .O_9_0_0_0(n98_O_9_0_0_0),
    .O_9_0_0_1(n98_O_9_0_0_1),
    .O_9_0_0_2(n98_O_9_0_0_2),
    .O_9_0_1_0(n98_O_9_0_1_0),
    .O_9_0_1_1(n98_O_9_0_1_1),
    .O_9_0_1_2(n98_O_9_0_1_2),
    .O_9_0_2_0(n98_O_9_0_2_0),
    .O_9_0_2_1(n98_O_9_0_2_1),
    .O_9_0_2_2(n98_O_9_0_2_2),
    .O_10_0_0_0(n98_O_10_0_0_0),
    .O_10_0_0_1(n98_O_10_0_0_1),
    .O_10_0_0_2(n98_O_10_0_0_2),
    .O_10_0_1_0(n98_O_10_0_1_0),
    .O_10_0_1_1(n98_O_10_0_1_1),
    .O_10_0_1_2(n98_O_10_0_1_2),
    .O_10_0_2_0(n98_O_10_0_2_0),
    .O_10_0_2_1(n98_O_10_0_2_1),
    .O_10_0_2_2(n98_O_10_0_2_2),
    .O_11_0_0_0(n98_O_11_0_0_0),
    .O_11_0_0_1(n98_O_11_0_0_1),
    .O_11_0_0_2(n98_O_11_0_0_2),
    .O_11_0_1_0(n98_O_11_0_1_0),
    .O_11_0_1_1(n98_O_11_0_1_1),
    .O_11_0_1_2(n98_O_11_0_1_2),
    .O_11_0_2_0(n98_O_11_0_2_0),
    .O_11_0_2_1(n98_O_11_0_2_1),
    .O_11_0_2_2(n98_O_11_0_2_2),
    .O_12_0_0_0(n98_O_12_0_0_0),
    .O_12_0_0_1(n98_O_12_0_0_1),
    .O_12_0_0_2(n98_O_12_0_0_2),
    .O_12_0_1_0(n98_O_12_0_1_0),
    .O_12_0_1_1(n98_O_12_0_1_1),
    .O_12_0_1_2(n98_O_12_0_1_2),
    .O_12_0_2_0(n98_O_12_0_2_0),
    .O_12_0_2_1(n98_O_12_0_2_1),
    .O_12_0_2_2(n98_O_12_0_2_2),
    .O_13_0_0_0(n98_O_13_0_0_0),
    .O_13_0_0_1(n98_O_13_0_0_1),
    .O_13_0_0_2(n98_O_13_0_0_2),
    .O_13_0_1_0(n98_O_13_0_1_0),
    .O_13_0_1_1(n98_O_13_0_1_1),
    .O_13_0_1_2(n98_O_13_0_1_2),
    .O_13_0_2_0(n98_O_13_0_2_0),
    .O_13_0_2_1(n98_O_13_0_2_1),
    .O_13_0_2_2(n98_O_13_0_2_2),
    .O_14_0_0_0(n98_O_14_0_0_0),
    .O_14_0_0_1(n98_O_14_0_0_1),
    .O_14_0_0_2(n98_O_14_0_0_2),
    .O_14_0_1_0(n98_O_14_0_1_0),
    .O_14_0_1_1(n98_O_14_0_1_1),
    .O_14_0_1_2(n98_O_14_0_1_2),
    .O_14_0_2_0(n98_O_14_0_2_0),
    .O_14_0_2_1(n98_O_14_0_2_1),
    .O_14_0_2_2(n98_O_14_0_2_2),
    .O_15_0_0_0(n98_O_15_0_0_0),
    .O_15_0_0_1(n98_O_15_0_0_1),
    .O_15_0_0_2(n98_O_15_0_0_2),
    .O_15_0_1_0(n98_O_15_0_1_0),
    .O_15_0_1_1(n98_O_15_0_1_1),
    .O_15_0_1_2(n98_O_15_0_1_2),
    .O_15_0_2_0(n98_O_15_0_2_0),
    .O_15_0_2_1(n98_O_15_0_2_1),
    .O_15_0_2_2(n98_O_15_0_2_2)
  );
  MapT_7 n105 ( // @[Top.scala 437:22]
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0_0(n105_I_0_0_0_0),
    .I_0_0_0_1(n105_I_0_0_0_1),
    .I_0_0_0_2(n105_I_0_0_0_2),
    .I_0_0_1_0(n105_I_0_0_1_0),
    .I_0_0_1_1(n105_I_0_0_1_1),
    .I_0_0_1_2(n105_I_0_0_1_2),
    .I_0_0_2_0(n105_I_0_0_2_0),
    .I_0_0_2_1(n105_I_0_0_2_1),
    .I_0_0_2_2(n105_I_0_0_2_2),
    .I_1_0_0_0(n105_I_1_0_0_0),
    .I_1_0_0_1(n105_I_1_0_0_1),
    .I_1_0_0_2(n105_I_1_0_0_2),
    .I_1_0_1_0(n105_I_1_0_1_0),
    .I_1_0_1_1(n105_I_1_0_1_1),
    .I_1_0_1_2(n105_I_1_0_1_2),
    .I_1_0_2_0(n105_I_1_0_2_0),
    .I_1_0_2_1(n105_I_1_0_2_1),
    .I_1_0_2_2(n105_I_1_0_2_2),
    .I_2_0_0_0(n105_I_2_0_0_0),
    .I_2_0_0_1(n105_I_2_0_0_1),
    .I_2_0_0_2(n105_I_2_0_0_2),
    .I_2_0_1_0(n105_I_2_0_1_0),
    .I_2_0_1_1(n105_I_2_0_1_1),
    .I_2_0_1_2(n105_I_2_0_1_2),
    .I_2_0_2_0(n105_I_2_0_2_0),
    .I_2_0_2_1(n105_I_2_0_2_1),
    .I_2_0_2_2(n105_I_2_0_2_2),
    .I_3_0_0_0(n105_I_3_0_0_0),
    .I_3_0_0_1(n105_I_3_0_0_1),
    .I_3_0_0_2(n105_I_3_0_0_2),
    .I_3_0_1_0(n105_I_3_0_1_0),
    .I_3_0_1_1(n105_I_3_0_1_1),
    .I_3_0_1_2(n105_I_3_0_1_2),
    .I_3_0_2_0(n105_I_3_0_2_0),
    .I_3_0_2_1(n105_I_3_0_2_1),
    .I_3_0_2_2(n105_I_3_0_2_2),
    .I_4_0_0_0(n105_I_4_0_0_0),
    .I_4_0_0_1(n105_I_4_0_0_1),
    .I_4_0_0_2(n105_I_4_0_0_2),
    .I_4_0_1_0(n105_I_4_0_1_0),
    .I_4_0_1_1(n105_I_4_0_1_1),
    .I_4_0_1_2(n105_I_4_0_1_2),
    .I_4_0_2_0(n105_I_4_0_2_0),
    .I_4_0_2_1(n105_I_4_0_2_1),
    .I_4_0_2_2(n105_I_4_0_2_2),
    .I_5_0_0_0(n105_I_5_0_0_0),
    .I_5_0_0_1(n105_I_5_0_0_1),
    .I_5_0_0_2(n105_I_5_0_0_2),
    .I_5_0_1_0(n105_I_5_0_1_0),
    .I_5_0_1_1(n105_I_5_0_1_1),
    .I_5_0_1_2(n105_I_5_0_1_2),
    .I_5_0_2_0(n105_I_5_0_2_0),
    .I_5_0_2_1(n105_I_5_0_2_1),
    .I_5_0_2_2(n105_I_5_0_2_2),
    .I_6_0_0_0(n105_I_6_0_0_0),
    .I_6_0_0_1(n105_I_6_0_0_1),
    .I_6_0_0_2(n105_I_6_0_0_2),
    .I_6_0_1_0(n105_I_6_0_1_0),
    .I_6_0_1_1(n105_I_6_0_1_1),
    .I_6_0_1_2(n105_I_6_0_1_2),
    .I_6_0_2_0(n105_I_6_0_2_0),
    .I_6_0_2_1(n105_I_6_0_2_1),
    .I_6_0_2_2(n105_I_6_0_2_2),
    .I_7_0_0_0(n105_I_7_0_0_0),
    .I_7_0_0_1(n105_I_7_0_0_1),
    .I_7_0_0_2(n105_I_7_0_0_2),
    .I_7_0_1_0(n105_I_7_0_1_0),
    .I_7_0_1_1(n105_I_7_0_1_1),
    .I_7_0_1_2(n105_I_7_0_1_2),
    .I_7_0_2_0(n105_I_7_0_2_0),
    .I_7_0_2_1(n105_I_7_0_2_1),
    .I_7_0_2_2(n105_I_7_0_2_2),
    .I_8_0_0_0(n105_I_8_0_0_0),
    .I_8_0_0_1(n105_I_8_0_0_1),
    .I_8_0_0_2(n105_I_8_0_0_2),
    .I_8_0_1_0(n105_I_8_0_1_0),
    .I_8_0_1_1(n105_I_8_0_1_1),
    .I_8_0_1_2(n105_I_8_0_1_2),
    .I_8_0_2_0(n105_I_8_0_2_0),
    .I_8_0_2_1(n105_I_8_0_2_1),
    .I_8_0_2_2(n105_I_8_0_2_2),
    .I_9_0_0_0(n105_I_9_0_0_0),
    .I_9_0_0_1(n105_I_9_0_0_1),
    .I_9_0_0_2(n105_I_9_0_0_2),
    .I_9_0_1_0(n105_I_9_0_1_0),
    .I_9_0_1_1(n105_I_9_0_1_1),
    .I_9_0_1_2(n105_I_9_0_1_2),
    .I_9_0_2_0(n105_I_9_0_2_0),
    .I_9_0_2_1(n105_I_9_0_2_1),
    .I_9_0_2_2(n105_I_9_0_2_2),
    .I_10_0_0_0(n105_I_10_0_0_0),
    .I_10_0_0_1(n105_I_10_0_0_1),
    .I_10_0_0_2(n105_I_10_0_0_2),
    .I_10_0_1_0(n105_I_10_0_1_0),
    .I_10_0_1_1(n105_I_10_0_1_1),
    .I_10_0_1_2(n105_I_10_0_1_2),
    .I_10_0_2_0(n105_I_10_0_2_0),
    .I_10_0_2_1(n105_I_10_0_2_1),
    .I_10_0_2_2(n105_I_10_0_2_2),
    .I_11_0_0_0(n105_I_11_0_0_0),
    .I_11_0_0_1(n105_I_11_0_0_1),
    .I_11_0_0_2(n105_I_11_0_0_2),
    .I_11_0_1_0(n105_I_11_0_1_0),
    .I_11_0_1_1(n105_I_11_0_1_1),
    .I_11_0_1_2(n105_I_11_0_1_2),
    .I_11_0_2_0(n105_I_11_0_2_0),
    .I_11_0_2_1(n105_I_11_0_2_1),
    .I_11_0_2_2(n105_I_11_0_2_2),
    .I_12_0_0_0(n105_I_12_0_0_0),
    .I_12_0_0_1(n105_I_12_0_0_1),
    .I_12_0_0_2(n105_I_12_0_0_2),
    .I_12_0_1_0(n105_I_12_0_1_0),
    .I_12_0_1_1(n105_I_12_0_1_1),
    .I_12_0_1_2(n105_I_12_0_1_2),
    .I_12_0_2_0(n105_I_12_0_2_0),
    .I_12_0_2_1(n105_I_12_0_2_1),
    .I_12_0_2_2(n105_I_12_0_2_2),
    .I_13_0_0_0(n105_I_13_0_0_0),
    .I_13_0_0_1(n105_I_13_0_0_1),
    .I_13_0_0_2(n105_I_13_0_0_2),
    .I_13_0_1_0(n105_I_13_0_1_0),
    .I_13_0_1_1(n105_I_13_0_1_1),
    .I_13_0_1_2(n105_I_13_0_1_2),
    .I_13_0_2_0(n105_I_13_0_2_0),
    .I_13_0_2_1(n105_I_13_0_2_1),
    .I_13_0_2_2(n105_I_13_0_2_2),
    .I_14_0_0_0(n105_I_14_0_0_0),
    .I_14_0_0_1(n105_I_14_0_0_1),
    .I_14_0_0_2(n105_I_14_0_0_2),
    .I_14_0_1_0(n105_I_14_0_1_0),
    .I_14_0_1_1(n105_I_14_0_1_1),
    .I_14_0_1_2(n105_I_14_0_1_2),
    .I_14_0_2_0(n105_I_14_0_2_0),
    .I_14_0_2_1(n105_I_14_0_2_1),
    .I_14_0_2_2(n105_I_14_0_2_2),
    .I_15_0_0_0(n105_I_15_0_0_0),
    .I_15_0_0_1(n105_I_15_0_0_1),
    .I_15_0_0_2(n105_I_15_0_0_2),
    .I_15_0_1_0(n105_I_15_0_1_0),
    .I_15_0_1_1(n105_I_15_0_1_1),
    .I_15_0_1_2(n105_I_15_0_1_2),
    .I_15_0_2_0(n105_I_15_0_2_0),
    .I_15_0_2_1(n105_I_15_0_2_1),
    .I_15_0_2_2(n105_I_15_0_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_0_0_1(n105_O_0_0_1),
    .O_0_0_2(n105_O_0_0_2),
    .O_0_1_0(n105_O_0_1_0),
    .O_0_1_1(n105_O_0_1_1),
    .O_0_1_2(n105_O_0_1_2),
    .O_0_2_0(n105_O_0_2_0),
    .O_0_2_1(n105_O_0_2_1),
    .O_0_2_2(n105_O_0_2_2),
    .O_1_0_0(n105_O_1_0_0),
    .O_1_0_1(n105_O_1_0_1),
    .O_1_0_2(n105_O_1_0_2),
    .O_1_1_0(n105_O_1_1_0),
    .O_1_1_1(n105_O_1_1_1),
    .O_1_1_2(n105_O_1_1_2),
    .O_1_2_0(n105_O_1_2_0),
    .O_1_2_1(n105_O_1_2_1),
    .O_1_2_2(n105_O_1_2_2),
    .O_2_0_0(n105_O_2_0_0),
    .O_2_0_1(n105_O_2_0_1),
    .O_2_0_2(n105_O_2_0_2),
    .O_2_1_0(n105_O_2_1_0),
    .O_2_1_1(n105_O_2_1_1),
    .O_2_1_2(n105_O_2_1_2),
    .O_2_2_0(n105_O_2_2_0),
    .O_2_2_1(n105_O_2_2_1),
    .O_2_2_2(n105_O_2_2_2),
    .O_3_0_0(n105_O_3_0_0),
    .O_3_0_1(n105_O_3_0_1),
    .O_3_0_2(n105_O_3_0_2),
    .O_3_1_0(n105_O_3_1_0),
    .O_3_1_1(n105_O_3_1_1),
    .O_3_1_2(n105_O_3_1_2),
    .O_3_2_0(n105_O_3_2_0),
    .O_3_2_1(n105_O_3_2_1),
    .O_3_2_2(n105_O_3_2_2),
    .O_4_0_0(n105_O_4_0_0),
    .O_4_0_1(n105_O_4_0_1),
    .O_4_0_2(n105_O_4_0_2),
    .O_4_1_0(n105_O_4_1_0),
    .O_4_1_1(n105_O_4_1_1),
    .O_4_1_2(n105_O_4_1_2),
    .O_4_2_0(n105_O_4_2_0),
    .O_4_2_1(n105_O_4_2_1),
    .O_4_2_2(n105_O_4_2_2),
    .O_5_0_0(n105_O_5_0_0),
    .O_5_0_1(n105_O_5_0_1),
    .O_5_0_2(n105_O_5_0_2),
    .O_5_1_0(n105_O_5_1_0),
    .O_5_1_1(n105_O_5_1_1),
    .O_5_1_2(n105_O_5_1_2),
    .O_5_2_0(n105_O_5_2_0),
    .O_5_2_1(n105_O_5_2_1),
    .O_5_2_2(n105_O_5_2_2),
    .O_6_0_0(n105_O_6_0_0),
    .O_6_0_1(n105_O_6_0_1),
    .O_6_0_2(n105_O_6_0_2),
    .O_6_1_0(n105_O_6_1_0),
    .O_6_1_1(n105_O_6_1_1),
    .O_6_1_2(n105_O_6_1_2),
    .O_6_2_0(n105_O_6_2_0),
    .O_6_2_1(n105_O_6_2_1),
    .O_6_2_2(n105_O_6_2_2),
    .O_7_0_0(n105_O_7_0_0),
    .O_7_0_1(n105_O_7_0_1),
    .O_7_0_2(n105_O_7_0_2),
    .O_7_1_0(n105_O_7_1_0),
    .O_7_1_1(n105_O_7_1_1),
    .O_7_1_2(n105_O_7_1_2),
    .O_7_2_0(n105_O_7_2_0),
    .O_7_2_1(n105_O_7_2_1),
    .O_7_2_2(n105_O_7_2_2),
    .O_8_0_0(n105_O_8_0_0),
    .O_8_0_1(n105_O_8_0_1),
    .O_8_0_2(n105_O_8_0_2),
    .O_8_1_0(n105_O_8_1_0),
    .O_8_1_1(n105_O_8_1_1),
    .O_8_1_2(n105_O_8_1_2),
    .O_8_2_0(n105_O_8_2_0),
    .O_8_2_1(n105_O_8_2_1),
    .O_8_2_2(n105_O_8_2_2),
    .O_9_0_0(n105_O_9_0_0),
    .O_9_0_1(n105_O_9_0_1),
    .O_9_0_2(n105_O_9_0_2),
    .O_9_1_0(n105_O_9_1_0),
    .O_9_1_1(n105_O_9_1_1),
    .O_9_1_2(n105_O_9_1_2),
    .O_9_2_0(n105_O_9_2_0),
    .O_9_2_1(n105_O_9_2_1),
    .O_9_2_2(n105_O_9_2_2),
    .O_10_0_0(n105_O_10_0_0),
    .O_10_0_1(n105_O_10_0_1),
    .O_10_0_2(n105_O_10_0_2),
    .O_10_1_0(n105_O_10_1_0),
    .O_10_1_1(n105_O_10_1_1),
    .O_10_1_2(n105_O_10_1_2),
    .O_10_2_0(n105_O_10_2_0),
    .O_10_2_1(n105_O_10_2_1),
    .O_10_2_2(n105_O_10_2_2),
    .O_11_0_0(n105_O_11_0_0),
    .O_11_0_1(n105_O_11_0_1),
    .O_11_0_2(n105_O_11_0_2),
    .O_11_1_0(n105_O_11_1_0),
    .O_11_1_1(n105_O_11_1_1),
    .O_11_1_2(n105_O_11_1_2),
    .O_11_2_0(n105_O_11_2_0),
    .O_11_2_1(n105_O_11_2_1),
    .O_11_2_2(n105_O_11_2_2),
    .O_12_0_0(n105_O_12_0_0),
    .O_12_0_1(n105_O_12_0_1),
    .O_12_0_2(n105_O_12_0_2),
    .O_12_1_0(n105_O_12_1_0),
    .O_12_1_1(n105_O_12_1_1),
    .O_12_1_2(n105_O_12_1_2),
    .O_12_2_0(n105_O_12_2_0),
    .O_12_2_1(n105_O_12_2_1),
    .O_12_2_2(n105_O_12_2_2),
    .O_13_0_0(n105_O_13_0_0),
    .O_13_0_1(n105_O_13_0_1),
    .O_13_0_2(n105_O_13_0_2),
    .O_13_1_0(n105_O_13_1_0),
    .O_13_1_1(n105_O_13_1_1),
    .O_13_1_2(n105_O_13_1_2),
    .O_13_2_0(n105_O_13_2_0),
    .O_13_2_1(n105_O_13_2_1),
    .O_13_2_2(n105_O_13_2_2),
    .O_14_0_0(n105_O_14_0_0),
    .O_14_0_1(n105_O_14_0_1),
    .O_14_0_2(n105_O_14_0_2),
    .O_14_1_0(n105_O_14_1_0),
    .O_14_1_1(n105_O_14_1_1),
    .O_14_1_2(n105_O_14_1_2),
    .O_14_2_0(n105_O_14_2_0),
    .O_14_2_1(n105_O_14_2_1),
    .O_14_2_2(n105_O_14_2_2),
    .O_15_0_0(n105_O_15_0_0),
    .O_15_0_1(n105_O_15_0_1),
    .O_15_0_2(n105_O_15_0_2),
    .O_15_1_0(n105_O_15_1_0),
    .O_15_1_1(n105_O_15_1_1),
    .O_15_1_2(n105_O_15_1_2),
    .O_15_2_0(n105_O_15_2_0),
    .O_15_2_1(n105_O_15_2_1),
    .O_15_2_2(n105_O_15_2_2)
  );
  Passthrough n106 ( // @[Top.scala 440:22]
    .valid_up(n106_valid_up),
    .valid_down(n106_valid_down),
    .I_0_0_0(n106_I_0_0_0),
    .I_0_0_1(n106_I_0_0_1),
    .I_0_0_2(n106_I_0_0_2),
    .I_0_1_0(n106_I_0_1_0),
    .I_0_1_1(n106_I_0_1_1),
    .I_0_1_2(n106_I_0_1_2),
    .I_0_2_0(n106_I_0_2_0),
    .I_0_2_1(n106_I_0_2_1),
    .I_0_2_2(n106_I_0_2_2),
    .I_1_0_0(n106_I_1_0_0),
    .I_1_0_1(n106_I_1_0_1),
    .I_1_0_2(n106_I_1_0_2),
    .I_1_1_0(n106_I_1_1_0),
    .I_1_1_1(n106_I_1_1_1),
    .I_1_1_2(n106_I_1_1_2),
    .I_1_2_0(n106_I_1_2_0),
    .I_1_2_1(n106_I_1_2_1),
    .I_1_2_2(n106_I_1_2_2),
    .I_2_0_0(n106_I_2_0_0),
    .I_2_0_1(n106_I_2_0_1),
    .I_2_0_2(n106_I_2_0_2),
    .I_2_1_0(n106_I_2_1_0),
    .I_2_1_1(n106_I_2_1_1),
    .I_2_1_2(n106_I_2_1_2),
    .I_2_2_0(n106_I_2_2_0),
    .I_2_2_1(n106_I_2_2_1),
    .I_2_2_2(n106_I_2_2_2),
    .I_3_0_0(n106_I_3_0_0),
    .I_3_0_1(n106_I_3_0_1),
    .I_3_0_2(n106_I_3_0_2),
    .I_3_1_0(n106_I_3_1_0),
    .I_3_1_1(n106_I_3_1_1),
    .I_3_1_2(n106_I_3_1_2),
    .I_3_2_0(n106_I_3_2_0),
    .I_3_2_1(n106_I_3_2_1),
    .I_3_2_2(n106_I_3_2_2),
    .I_4_0_0(n106_I_4_0_0),
    .I_4_0_1(n106_I_4_0_1),
    .I_4_0_2(n106_I_4_0_2),
    .I_4_1_0(n106_I_4_1_0),
    .I_4_1_1(n106_I_4_1_1),
    .I_4_1_2(n106_I_4_1_2),
    .I_4_2_0(n106_I_4_2_0),
    .I_4_2_1(n106_I_4_2_1),
    .I_4_2_2(n106_I_4_2_2),
    .I_5_0_0(n106_I_5_0_0),
    .I_5_0_1(n106_I_5_0_1),
    .I_5_0_2(n106_I_5_0_2),
    .I_5_1_0(n106_I_5_1_0),
    .I_5_1_1(n106_I_5_1_1),
    .I_5_1_2(n106_I_5_1_2),
    .I_5_2_0(n106_I_5_2_0),
    .I_5_2_1(n106_I_5_2_1),
    .I_5_2_2(n106_I_5_2_2),
    .I_6_0_0(n106_I_6_0_0),
    .I_6_0_1(n106_I_6_0_1),
    .I_6_0_2(n106_I_6_0_2),
    .I_6_1_0(n106_I_6_1_0),
    .I_6_1_1(n106_I_6_1_1),
    .I_6_1_2(n106_I_6_1_2),
    .I_6_2_0(n106_I_6_2_0),
    .I_6_2_1(n106_I_6_2_1),
    .I_6_2_2(n106_I_6_2_2),
    .I_7_0_0(n106_I_7_0_0),
    .I_7_0_1(n106_I_7_0_1),
    .I_7_0_2(n106_I_7_0_2),
    .I_7_1_0(n106_I_7_1_0),
    .I_7_1_1(n106_I_7_1_1),
    .I_7_1_2(n106_I_7_1_2),
    .I_7_2_0(n106_I_7_2_0),
    .I_7_2_1(n106_I_7_2_1),
    .I_7_2_2(n106_I_7_2_2),
    .I_8_0_0(n106_I_8_0_0),
    .I_8_0_1(n106_I_8_0_1),
    .I_8_0_2(n106_I_8_0_2),
    .I_8_1_0(n106_I_8_1_0),
    .I_8_1_1(n106_I_8_1_1),
    .I_8_1_2(n106_I_8_1_2),
    .I_8_2_0(n106_I_8_2_0),
    .I_8_2_1(n106_I_8_2_1),
    .I_8_2_2(n106_I_8_2_2),
    .I_9_0_0(n106_I_9_0_0),
    .I_9_0_1(n106_I_9_0_1),
    .I_9_0_2(n106_I_9_0_2),
    .I_9_1_0(n106_I_9_1_0),
    .I_9_1_1(n106_I_9_1_1),
    .I_9_1_2(n106_I_9_1_2),
    .I_9_2_0(n106_I_9_2_0),
    .I_9_2_1(n106_I_9_2_1),
    .I_9_2_2(n106_I_9_2_2),
    .I_10_0_0(n106_I_10_0_0),
    .I_10_0_1(n106_I_10_0_1),
    .I_10_0_2(n106_I_10_0_2),
    .I_10_1_0(n106_I_10_1_0),
    .I_10_1_1(n106_I_10_1_1),
    .I_10_1_2(n106_I_10_1_2),
    .I_10_2_0(n106_I_10_2_0),
    .I_10_2_1(n106_I_10_2_1),
    .I_10_2_2(n106_I_10_2_2),
    .I_11_0_0(n106_I_11_0_0),
    .I_11_0_1(n106_I_11_0_1),
    .I_11_0_2(n106_I_11_0_2),
    .I_11_1_0(n106_I_11_1_0),
    .I_11_1_1(n106_I_11_1_1),
    .I_11_1_2(n106_I_11_1_2),
    .I_11_2_0(n106_I_11_2_0),
    .I_11_2_1(n106_I_11_2_1),
    .I_11_2_2(n106_I_11_2_2),
    .I_12_0_0(n106_I_12_0_0),
    .I_12_0_1(n106_I_12_0_1),
    .I_12_0_2(n106_I_12_0_2),
    .I_12_1_0(n106_I_12_1_0),
    .I_12_1_1(n106_I_12_1_1),
    .I_12_1_2(n106_I_12_1_2),
    .I_12_2_0(n106_I_12_2_0),
    .I_12_2_1(n106_I_12_2_1),
    .I_12_2_2(n106_I_12_2_2),
    .I_13_0_0(n106_I_13_0_0),
    .I_13_0_1(n106_I_13_0_1),
    .I_13_0_2(n106_I_13_0_2),
    .I_13_1_0(n106_I_13_1_0),
    .I_13_1_1(n106_I_13_1_1),
    .I_13_1_2(n106_I_13_1_2),
    .I_13_2_0(n106_I_13_2_0),
    .I_13_2_1(n106_I_13_2_1),
    .I_13_2_2(n106_I_13_2_2),
    .I_14_0_0(n106_I_14_0_0),
    .I_14_0_1(n106_I_14_0_1),
    .I_14_0_2(n106_I_14_0_2),
    .I_14_1_0(n106_I_14_1_0),
    .I_14_1_1(n106_I_14_1_1),
    .I_14_1_2(n106_I_14_1_2),
    .I_14_2_0(n106_I_14_2_0),
    .I_14_2_1(n106_I_14_2_1),
    .I_14_2_2(n106_I_14_2_2),
    .I_15_0_0(n106_I_15_0_0),
    .I_15_0_1(n106_I_15_0_1),
    .I_15_0_2(n106_I_15_0_2),
    .I_15_1_0(n106_I_15_1_0),
    .I_15_1_1(n106_I_15_1_1),
    .I_15_1_2(n106_I_15_1_2),
    .I_15_2_0(n106_I_15_2_0),
    .I_15_2_1(n106_I_15_2_1),
    .I_15_2_2(n106_I_15_2_2),
    .O_0_0_0(n106_O_0_0_0),
    .O_0_0_1(n106_O_0_0_1),
    .O_0_0_2(n106_O_0_0_2),
    .O_0_1_0(n106_O_0_1_0),
    .O_0_1_1(n106_O_0_1_1),
    .O_0_1_2(n106_O_0_1_2),
    .O_0_2_0(n106_O_0_2_0),
    .O_0_2_1(n106_O_0_2_1),
    .O_0_2_2(n106_O_0_2_2),
    .O_1_0_0(n106_O_1_0_0),
    .O_1_0_1(n106_O_1_0_1),
    .O_1_0_2(n106_O_1_0_2),
    .O_1_1_0(n106_O_1_1_0),
    .O_1_1_1(n106_O_1_1_1),
    .O_1_1_2(n106_O_1_1_2),
    .O_1_2_0(n106_O_1_2_0),
    .O_1_2_1(n106_O_1_2_1),
    .O_1_2_2(n106_O_1_2_2),
    .O_2_0_0(n106_O_2_0_0),
    .O_2_0_1(n106_O_2_0_1),
    .O_2_0_2(n106_O_2_0_2),
    .O_2_1_0(n106_O_2_1_0),
    .O_2_1_1(n106_O_2_1_1),
    .O_2_1_2(n106_O_2_1_2),
    .O_2_2_0(n106_O_2_2_0),
    .O_2_2_1(n106_O_2_2_1),
    .O_2_2_2(n106_O_2_2_2),
    .O_3_0_0(n106_O_3_0_0),
    .O_3_0_1(n106_O_3_0_1),
    .O_3_0_2(n106_O_3_0_2),
    .O_3_1_0(n106_O_3_1_0),
    .O_3_1_1(n106_O_3_1_1),
    .O_3_1_2(n106_O_3_1_2),
    .O_3_2_0(n106_O_3_2_0),
    .O_3_2_1(n106_O_3_2_1),
    .O_3_2_2(n106_O_3_2_2),
    .O_4_0_0(n106_O_4_0_0),
    .O_4_0_1(n106_O_4_0_1),
    .O_4_0_2(n106_O_4_0_2),
    .O_4_1_0(n106_O_4_1_0),
    .O_4_1_1(n106_O_4_1_1),
    .O_4_1_2(n106_O_4_1_2),
    .O_4_2_0(n106_O_4_2_0),
    .O_4_2_1(n106_O_4_2_1),
    .O_4_2_2(n106_O_4_2_2),
    .O_5_0_0(n106_O_5_0_0),
    .O_5_0_1(n106_O_5_0_1),
    .O_5_0_2(n106_O_5_0_2),
    .O_5_1_0(n106_O_5_1_0),
    .O_5_1_1(n106_O_5_1_1),
    .O_5_1_2(n106_O_5_1_2),
    .O_5_2_0(n106_O_5_2_0),
    .O_5_2_1(n106_O_5_2_1),
    .O_5_2_2(n106_O_5_2_2),
    .O_6_0_0(n106_O_6_0_0),
    .O_6_0_1(n106_O_6_0_1),
    .O_6_0_2(n106_O_6_0_2),
    .O_6_1_0(n106_O_6_1_0),
    .O_6_1_1(n106_O_6_1_1),
    .O_6_1_2(n106_O_6_1_2),
    .O_6_2_0(n106_O_6_2_0),
    .O_6_2_1(n106_O_6_2_1),
    .O_6_2_2(n106_O_6_2_2),
    .O_7_0_0(n106_O_7_0_0),
    .O_7_0_1(n106_O_7_0_1),
    .O_7_0_2(n106_O_7_0_2),
    .O_7_1_0(n106_O_7_1_0),
    .O_7_1_1(n106_O_7_1_1),
    .O_7_1_2(n106_O_7_1_2),
    .O_7_2_0(n106_O_7_2_0),
    .O_7_2_1(n106_O_7_2_1),
    .O_7_2_2(n106_O_7_2_2),
    .O_8_0_0(n106_O_8_0_0),
    .O_8_0_1(n106_O_8_0_1),
    .O_8_0_2(n106_O_8_0_2),
    .O_8_1_0(n106_O_8_1_0),
    .O_8_1_1(n106_O_8_1_1),
    .O_8_1_2(n106_O_8_1_2),
    .O_8_2_0(n106_O_8_2_0),
    .O_8_2_1(n106_O_8_2_1),
    .O_8_2_2(n106_O_8_2_2),
    .O_9_0_0(n106_O_9_0_0),
    .O_9_0_1(n106_O_9_0_1),
    .O_9_0_2(n106_O_9_0_2),
    .O_9_1_0(n106_O_9_1_0),
    .O_9_1_1(n106_O_9_1_1),
    .O_9_1_2(n106_O_9_1_2),
    .O_9_2_0(n106_O_9_2_0),
    .O_9_2_1(n106_O_9_2_1),
    .O_9_2_2(n106_O_9_2_2),
    .O_10_0_0(n106_O_10_0_0),
    .O_10_0_1(n106_O_10_0_1),
    .O_10_0_2(n106_O_10_0_2),
    .O_10_1_0(n106_O_10_1_0),
    .O_10_1_1(n106_O_10_1_1),
    .O_10_1_2(n106_O_10_1_2),
    .O_10_2_0(n106_O_10_2_0),
    .O_10_2_1(n106_O_10_2_1),
    .O_10_2_2(n106_O_10_2_2),
    .O_11_0_0(n106_O_11_0_0),
    .O_11_0_1(n106_O_11_0_1),
    .O_11_0_2(n106_O_11_0_2),
    .O_11_1_0(n106_O_11_1_0),
    .O_11_1_1(n106_O_11_1_1),
    .O_11_1_2(n106_O_11_1_2),
    .O_11_2_0(n106_O_11_2_0),
    .O_11_2_1(n106_O_11_2_1),
    .O_11_2_2(n106_O_11_2_2),
    .O_12_0_0(n106_O_12_0_0),
    .O_12_0_1(n106_O_12_0_1),
    .O_12_0_2(n106_O_12_0_2),
    .O_12_1_0(n106_O_12_1_0),
    .O_12_1_1(n106_O_12_1_1),
    .O_12_1_2(n106_O_12_1_2),
    .O_12_2_0(n106_O_12_2_0),
    .O_12_2_1(n106_O_12_2_1),
    .O_12_2_2(n106_O_12_2_2),
    .O_13_0_0(n106_O_13_0_0),
    .O_13_0_1(n106_O_13_0_1),
    .O_13_0_2(n106_O_13_0_2),
    .O_13_1_0(n106_O_13_1_0),
    .O_13_1_1(n106_O_13_1_1),
    .O_13_1_2(n106_O_13_1_2),
    .O_13_2_0(n106_O_13_2_0),
    .O_13_2_1(n106_O_13_2_1),
    .O_13_2_2(n106_O_13_2_2),
    .O_14_0_0(n106_O_14_0_0),
    .O_14_0_1(n106_O_14_0_1),
    .O_14_0_2(n106_O_14_0_2),
    .O_14_1_0(n106_O_14_1_0),
    .O_14_1_1(n106_O_14_1_1),
    .O_14_1_2(n106_O_14_1_2),
    .O_14_2_0(n106_O_14_2_0),
    .O_14_2_1(n106_O_14_2_1),
    .O_14_2_2(n106_O_14_2_2),
    .O_15_0_0(n106_O_15_0_0),
    .O_15_0_1(n106_O_15_0_1),
    .O_15_0_2(n106_O_15_0_2),
    .O_15_1_0(n106_O_15_1_0),
    .O_15_1_1(n106_O_15_1_1),
    .O_15_1_2(n106_O_15_1_2),
    .O_15_2_0(n106_O_15_2_0),
    .O_15_2_1(n106_O_15_2_1),
    .O_15_2_2(n106_O_15_2_2)
  );
  MapT_12 n443 ( // @[Top.scala 443:22]
    .clock(n443_clock),
    .reset(n443_reset),
    .valid_up(n443_valid_up),
    .valid_down(n443_valid_down),
    .I_0_0_0(n443_I_0_0_0),
    .I_0_0_1(n443_I_0_0_1),
    .I_0_0_2(n443_I_0_0_2),
    .I_0_1_0(n443_I_0_1_0),
    .I_0_1_1(n443_I_0_1_1),
    .I_0_1_2(n443_I_0_1_2),
    .I_0_2_0(n443_I_0_2_0),
    .I_0_2_1(n443_I_0_2_1),
    .I_0_2_2(n443_I_0_2_2),
    .I_1_0_0(n443_I_1_0_0),
    .I_1_0_1(n443_I_1_0_1),
    .I_1_0_2(n443_I_1_0_2),
    .I_1_1_0(n443_I_1_1_0),
    .I_1_1_1(n443_I_1_1_1),
    .I_1_1_2(n443_I_1_1_2),
    .I_1_2_0(n443_I_1_2_0),
    .I_1_2_1(n443_I_1_2_1),
    .I_1_2_2(n443_I_1_2_2),
    .I_2_0_0(n443_I_2_0_0),
    .I_2_0_1(n443_I_2_0_1),
    .I_2_0_2(n443_I_2_0_2),
    .I_2_1_0(n443_I_2_1_0),
    .I_2_1_1(n443_I_2_1_1),
    .I_2_1_2(n443_I_2_1_2),
    .I_2_2_0(n443_I_2_2_0),
    .I_2_2_1(n443_I_2_2_1),
    .I_2_2_2(n443_I_2_2_2),
    .I_3_0_0(n443_I_3_0_0),
    .I_3_0_1(n443_I_3_0_1),
    .I_3_0_2(n443_I_3_0_2),
    .I_3_1_0(n443_I_3_1_0),
    .I_3_1_1(n443_I_3_1_1),
    .I_3_1_2(n443_I_3_1_2),
    .I_3_2_0(n443_I_3_2_0),
    .I_3_2_1(n443_I_3_2_1),
    .I_3_2_2(n443_I_3_2_2),
    .I_4_0_0(n443_I_4_0_0),
    .I_4_0_1(n443_I_4_0_1),
    .I_4_0_2(n443_I_4_0_2),
    .I_4_1_0(n443_I_4_1_0),
    .I_4_1_1(n443_I_4_1_1),
    .I_4_1_2(n443_I_4_1_2),
    .I_4_2_0(n443_I_4_2_0),
    .I_4_2_1(n443_I_4_2_1),
    .I_4_2_2(n443_I_4_2_2),
    .I_5_0_0(n443_I_5_0_0),
    .I_5_0_1(n443_I_5_0_1),
    .I_5_0_2(n443_I_5_0_2),
    .I_5_1_0(n443_I_5_1_0),
    .I_5_1_1(n443_I_5_1_1),
    .I_5_1_2(n443_I_5_1_2),
    .I_5_2_0(n443_I_5_2_0),
    .I_5_2_1(n443_I_5_2_1),
    .I_5_2_2(n443_I_5_2_2),
    .I_6_0_0(n443_I_6_0_0),
    .I_6_0_1(n443_I_6_0_1),
    .I_6_0_2(n443_I_6_0_2),
    .I_6_1_0(n443_I_6_1_0),
    .I_6_1_1(n443_I_6_1_1),
    .I_6_1_2(n443_I_6_1_2),
    .I_6_2_0(n443_I_6_2_0),
    .I_6_2_1(n443_I_6_2_1),
    .I_6_2_2(n443_I_6_2_2),
    .I_7_0_0(n443_I_7_0_0),
    .I_7_0_1(n443_I_7_0_1),
    .I_7_0_2(n443_I_7_0_2),
    .I_7_1_0(n443_I_7_1_0),
    .I_7_1_1(n443_I_7_1_1),
    .I_7_1_2(n443_I_7_1_2),
    .I_7_2_0(n443_I_7_2_0),
    .I_7_2_1(n443_I_7_2_1),
    .I_7_2_2(n443_I_7_2_2),
    .I_8_0_0(n443_I_8_0_0),
    .I_8_0_1(n443_I_8_0_1),
    .I_8_0_2(n443_I_8_0_2),
    .I_8_1_0(n443_I_8_1_0),
    .I_8_1_1(n443_I_8_1_1),
    .I_8_1_2(n443_I_8_1_2),
    .I_8_2_0(n443_I_8_2_0),
    .I_8_2_1(n443_I_8_2_1),
    .I_8_2_2(n443_I_8_2_2),
    .I_9_0_0(n443_I_9_0_0),
    .I_9_0_1(n443_I_9_0_1),
    .I_9_0_2(n443_I_9_0_2),
    .I_9_1_0(n443_I_9_1_0),
    .I_9_1_1(n443_I_9_1_1),
    .I_9_1_2(n443_I_9_1_2),
    .I_9_2_0(n443_I_9_2_0),
    .I_9_2_1(n443_I_9_2_1),
    .I_9_2_2(n443_I_9_2_2),
    .I_10_0_0(n443_I_10_0_0),
    .I_10_0_1(n443_I_10_0_1),
    .I_10_0_2(n443_I_10_0_2),
    .I_10_1_0(n443_I_10_1_0),
    .I_10_1_1(n443_I_10_1_1),
    .I_10_1_2(n443_I_10_1_2),
    .I_10_2_0(n443_I_10_2_0),
    .I_10_2_1(n443_I_10_2_1),
    .I_10_2_2(n443_I_10_2_2),
    .I_11_0_0(n443_I_11_0_0),
    .I_11_0_1(n443_I_11_0_1),
    .I_11_0_2(n443_I_11_0_2),
    .I_11_1_0(n443_I_11_1_0),
    .I_11_1_1(n443_I_11_1_1),
    .I_11_1_2(n443_I_11_1_2),
    .I_11_2_0(n443_I_11_2_0),
    .I_11_2_1(n443_I_11_2_1),
    .I_11_2_2(n443_I_11_2_2),
    .I_12_0_0(n443_I_12_0_0),
    .I_12_0_1(n443_I_12_0_1),
    .I_12_0_2(n443_I_12_0_2),
    .I_12_1_0(n443_I_12_1_0),
    .I_12_1_1(n443_I_12_1_1),
    .I_12_1_2(n443_I_12_1_2),
    .I_12_2_0(n443_I_12_2_0),
    .I_12_2_1(n443_I_12_2_1),
    .I_12_2_2(n443_I_12_2_2),
    .I_13_0_0(n443_I_13_0_0),
    .I_13_0_1(n443_I_13_0_1),
    .I_13_0_2(n443_I_13_0_2),
    .I_13_1_0(n443_I_13_1_0),
    .I_13_1_1(n443_I_13_1_1),
    .I_13_1_2(n443_I_13_1_2),
    .I_13_2_0(n443_I_13_2_0),
    .I_13_2_1(n443_I_13_2_1),
    .I_13_2_2(n443_I_13_2_2),
    .I_14_0_0(n443_I_14_0_0),
    .I_14_0_1(n443_I_14_0_1),
    .I_14_0_2(n443_I_14_0_2),
    .I_14_1_0(n443_I_14_1_0),
    .I_14_1_1(n443_I_14_1_1),
    .I_14_1_2(n443_I_14_1_2),
    .I_14_2_0(n443_I_14_2_0),
    .I_14_2_1(n443_I_14_2_1),
    .I_14_2_2(n443_I_14_2_2),
    .I_15_0_0(n443_I_15_0_0),
    .I_15_0_1(n443_I_15_0_1),
    .I_15_0_2(n443_I_15_0_2),
    .I_15_1_0(n443_I_15_1_0),
    .I_15_1_1(n443_I_15_1_1),
    .I_15_1_2(n443_I_15_1_2),
    .I_15_2_0(n443_I_15_2_0),
    .I_15_2_1(n443_I_15_2_1),
    .I_15_2_2(n443_I_15_2_2),
    .O_0_0_0_t0b(n443_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(n443_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(n443_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(n443_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(n443_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(n443_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(n443_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(n443_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(n443_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(n443_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(n443_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(n443_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(n443_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(n443_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(n443_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(n443_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(n443_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(n443_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(n443_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(n443_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(n443_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(n443_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(n443_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(n443_O_7_0_0_t1b_t1b),
    .O_8_0_0_t0b(n443_O_8_0_0_t0b),
    .O_8_0_0_t1b_t0b(n443_O_8_0_0_t1b_t0b),
    .O_8_0_0_t1b_t1b(n443_O_8_0_0_t1b_t1b),
    .O_9_0_0_t0b(n443_O_9_0_0_t0b),
    .O_9_0_0_t1b_t0b(n443_O_9_0_0_t1b_t0b),
    .O_9_0_0_t1b_t1b(n443_O_9_0_0_t1b_t1b),
    .O_10_0_0_t0b(n443_O_10_0_0_t0b),
    .O_10_0_0_t1b_t0b(n443_O_10_0_0_t1b_t0b),
    .O_10_0_0_t1b_t1b(n443_O_10_0_0_t1b_t1b),
    .O_11_0_0_t0b(n443_O_11_0_0_t0b),
    .O_11_0_0_t1b_t0b(n443_O_11_0_0_t1b_t0b),
    .O_11_0_0_t1b_t1b(n443_O_11_0_0_t1b_t1b),
    .O_12_0_0_t0b(n443_O_12_0_0_t0b),
    .O_12_0_0_t1b_t0b(n443_O_12_0_0_t1b_t0b),
    .O_12_0_0_t1b_t1b(n443_O_12_0_0_t1b_t1b),
    .O_13_0_0_t0b(n443_O_13_0_0_t0b),
    .O_13_0_0_t1b_t0b(n443_O_13_0_0_t1b_t0b),
    .O_13_0_0_t1b_t1b(n443_O_13_0_0_t1b_t1b),
    .O_14_0_0_t0b(n443_O_14_0_0_t0b),
    .O_14_0_0_t1b_t0b(n443_O_14_0_0_t1b_t0b),
    .O_14_0_0_t1b_t1b(n443_O_14_0_0_t1b_t1b),
    .O_15_0_0_t0b(n443_O_15_0_0_t0b),
    .O_15_0_0_t1b_t0b(n443_O_15_0_0_t1b_t0b),
    .O_15_0_0_t1b_t1b(n443_O_15_0_0_t1b_t1b)
  );
  Passthrough_1 n444 ( // @[Top.scala 446:22]
    .valid_up(n444_valid_up),
    .valid_down(n444_valid_down),
    .I_0_0_0_t0b(n444_I_0_0_0_t0b),
    .I_0_0_0_t1b_t0b(n444_I_0_0_0_t1b_t0b),
    .I_0_0_0_t1b_t1b(n444_I_0_0_0_t1b_t1b),
    .I_1_0_0_t0b(n444_I_1_0_0_t0b),
    .I_1_0_0_t1b_t0b(n444_I_1_0_0_t1b_t0b),
    .I_1_0_0_t1b_t1b(n444_I_1_0_0_t1b_t1b),
    .I_2_0_0_t0b(n444_I_2_0_0_t0b),
    .I_2_0_0_t1b_t0b(n444_I_2_0_0_t1b_t0b),
    .I_2_0_0_t1b_t1b(n444_I_2_0_0_t1b_t1b),
    .I_3_0_0_t0b(n444_I_3_0_0_t0b),
    .I_3_0_0_t1b_t0b(n444_I_3_0_0_t1b_t0b),
    .I_3_0_0_t1b_t1b(n444_I_3_0_0_t1b_t1b),
    .I_4_0_0_t0b(n444_I_4_0_0_t0b),
    .I_4_0_0_t1b_t0b(n444_I_4_0_0_t1b_t0b),
    .I_4_0_0_t1b_t1b(n444_I_4_0_0_t1b_t1b),
    .I_5_0_0_t0b(n444_I_5_0_0_t0b),
    .I_5_0_0_t1b_t0b(n444_I_5_0_0_t1b_t0b),
    .I_5_0_0_t1b_t1b(n444_I_5_0_0_t1b_t1b),
    .I_6_0_0_t0b(n444_I_6_0_0_t0b),
    .I_6_0_0_t1b_t0b(n444_I_6_0_0_t1b_t0b),
    .I_6_0_0_t1b_t1b(n444_I_6_0_0_t1b_t1b),
    .I_7_0_0_t0b(n444_I_7_0_0_t0b),
    .I_7_0_0_t1b_t0b(n444_I_7_0_0_t1b_t0b),
    .I_7_0_0_t1b_t1b(n444_I_7_0_0_t1b_t1b),
    .I_8_0_0_t0b(n444_I_8_0_0_t0b),
    .I_8_0_0_t1b_t0b(n444_I_8_0_0_t1b_t0b),
    .I_8_0_0_t1b_t1b(n444_I_8_0_0_t1b_t1b),
    .I_9_0_0_t0b(n444_I_9_0_0_t0b),
    .I_9_0_0_t1b_t0b(n444_I_9_0_0_t1b_t0b),
    .I_9_0_0_t1b_t1b(n444_I_9_0_0_t1b_t1b),
    .I_10_0_0_t0b(n444_I_10_0_0_t0b),
    .I_10_0_0_t1b_t0b(n444_I_10_0_0_t1b_t0b),
    .I_10_0_0_t1b_t1b(n444_I_10_0_0_t1b_t1b),
    .I_11_0_0_t0b(n444_I_11_0_0_t0b),
    .I_11_0_0_t1b_t0b(n444_I_11_0_0_t1b_t0b),
    .I_11_0_0_t1b_t1b(n444_I_11_0_0_t1b_t1b),
    .I_12_0_0_t0b(n444_I_12_0_0_t0b),
    .I_12_0_0_t1b_t0b(n444_I_12_0_0_t1b_t0b),
    .I_12_0_0_t1b_t1b(n444_I_12_0_0_t1b_t1b),
    .I_13_0_0_t0b(n444_I_13_0_0_t0b),
    .I_13_0_0_t1b_t0b(n444_I_13_0_0_t1b_t0b),
    .I_13_0_0_t1b_t1b(n444_I_13_0_0_t1b_t1b),
    .I_14_0_0_t0b(n444_I_14_0_0_t0b),
    .I_14_0_0_t1b_t0b(n444_I_14_0_0_t1b_t0b),
    .I_14_0_0_t1b_t1b(n444_I_14_0_0_t1b_t1b),
    .I_15_0_0_t0b(n444_I_15_0_0_t0b),
    .I_15_0_0_t1b_t0b(n444_I_15_0_0_t1b_t0b),
    .I_15_0_0_t1b_t1b(n444_I_15_0_0_t1b_t1b),
    .O_0_0_0_t0b(n444_O_0_0_0_t0b),
    .O_0_0_0_t1b_t0b(n444_O_0_0_0_t1b_t0b),
    .O_0_0_0_t1b_t1b(n444_O_0_0_0_t1b_t1b),
    .O_1_0_0_t0b(n444_O_1_0_0_t0b),
    .O_1_0_0_t1b_t0b(n444_O_1_0_0_t1b_t0b),
    .O_1_0_0_t1b_t1b(n444_O_1_0_0_t1b_t1b),
    .O_2_0_0_t0b(n444_O_2_0_0_t0b),
    .O_2_0_0_t1b_t0b(n444_O_2_0_0_t1b_t0b),
    .O_2_0_0_t1b_t1b(n444_O_2_0_0_t1b_t1b),
    .O_3_0_0_t0b(n444_O_3_0_0_t0b),
    .O_3_0_0_t1b_t0b(n444_O_3_0_0_t1b_t0b),
    .O_3_0_0_t1b_t1b(n444_O_3_0_0_t1b_t1b),
    .O_4_0_0_t0b(n444_O_4_0_0_t0b),
    .O_4_0_0_t1b_t0b(n444_O_4_0_0_t1b_t0b),
    .O_4_0_0_t1b_t1b(n444_O_4_0_0_t1b_t1b),
    .O_5_0_0_t0b(n444_O_5_0_0_t0b),
    .O_5_0_0_t1b_t0b(n444_O_5_0_0_t1b_t0b),
    .O_5_0_0_t1b_t1b(n444_O_5_0_0_t1b_t1b),
    .O_6_0_0_t0b(n444_O_6_0_0_t0b),
    .O_6_0_0_t1b_t0b(n444_O_6_0_0_t1b_t0b),
    .O_6_0_0_t1b_t1b(n444_O_6_0_0_t1b_t1b),
    .O_7_0_0_t0b(n444_O_7_0_0_t0b),
    .O_7_0_0_t1b_t0b(n444_O_7_0_0_t1b_t0b),
    .O_7_0_0_t1b_t1b(n444_O_7_0_0_t1b_t1b),
    .O_8_0_0_t0b(n444_O_8_0_0_t0b),
    .O_8_0_0_t1b_t0b(n444_O_8_0_0_t1b_t0b),
    .O_8_0_0_t1b_t1b(n444_O_8_0_0_t1b_t1b),
    .O_9_0_0_t0b(n444_O_9_0_0_t0b),
    .O_9_0_0_t1b_t0b(n444_O_9_0_0_t1b_t0b),
    .O_9_0_0_t1b_t1b(n444_O_9_0_0_t1b_t1b),
    .O_10_0_0_t0b(n444_O_10_0_0_t0b),
    .O_10_0_0_t1b_t0b(n444_O_10_0_0_t1b_t0b),
    .O_10_0_0_t1b_t1b(n444_O_10_0_0_t1b_t1b),
    .O_11_0_0_t0b(n444_O_11_0_0_t0b),
    .O_11_0_0_t1b_t0b(n444_O_11_0_0_t1b_t0b),
    .O_11_0_0_t1b_t1b(n444_O_11_0_0_t1b_t1b),
    .O_12_0_0_t0b(n444_O_12_0_0_t0b),
    .O_12_0_0_t1b_t0b(n444_O_12_0_0_t1b_t0b),
    .O_12_0_0_t1b_t1b(n444_O_12_0_0_t1b_t1b),
    .O_13_0_0_t0b(n444_O_13_0_0_t0b),
    .O_13_0_0_t1b_t0b(n444_O_13_0_0_t1b_t0b),
    .O_13_0_0_t1b_t1b(n444_O_13_0_0_t1b_t1b),
    .O_14_0_0_t0b(n444_O_14_0_0_t0b),
    .O_14_0_0_t1b_t0b(n444_O_14_0_0_t1b_t0b),
    .O_14_0_0_t1b_t1b(n444_O_14_0_0_t1b_t1b),
    .O_15_0_0_t0b(n444_O_15_0_0_t0b),
    .O_15_0_0_t1b_t0b(n444_O_15_0_0_t1b_t0b),
    .O_15_0_0_t1b_t1b(n444_O_15_0_0_t1b_t1b)
  );
  Passthrough_2 n445 ( // @[Top.scala 449:22]
    .valid_up(n445_valid_up),
    .valid_down(n445_valid_down),
    .I_0_0_0_t0b(n445_I_0_0_0_t0b),
    .I_0_0_0_t1b_t0b(n445_I_0_0_0_t1b_t0b),
    .I_0_0_0_t1b_t1b(n445_I_0_0_0_t1b_t1b),
    .I_1_0_0_t0b(n445_I_1_0_0_t0b),
    .I_1_0_0_t1b_t0b(n445_I_1_0_0_t1b_t0b),
    .I_1_0_0_t1b_t1b(n445_I_1_0_0_t1b_t1b),
    .I_2_0_0_t0b(n445_I_2_0_0_t0b),
    .I_2_0_0_t1b_t0b(n445_I_2_0_0_t1b_t0b),
    .I_2_0_0_t1b_t1b(n445_I_2_0_0_t1b_t1b),
    .I_3_0_0_t0b(n445_I_3_0_0_t0b),
    .I_3_0_0_t1b_t0b(n445_I_3_0_0_t1b_t0b),
    .I_3_0_0_t1b_t1b(n445_I_3_0_0_t1b_t1b),
    .I_4_0_0_t0b(n445_I_4_0_0_t0b),
    .I_4_0_0_t1b_t0b(n445_I_4_0_0_t1b_t0b),
    .I_4_0_0_t1b_t1b(n445_I_4_0_0_t1b_t1b),
    .I_5_0_0_t0b(n445_I_5_0_0_t0b),
    .I_5_0_0_t1b_t0b(n445_I_5_0_0_t1b_t0b),
    .I_5_0_0_t1b_t1b(n445_I_5_0_0_t1b_t1b),
    .I_6_0_0_t0b(n445_I_6_0_0_t0b),
    .I_6_0_0_t1b_t0b(n445_I_6_0_0_t1b_t0b),
    .I_6_0_0_t1b_t1b(n445_I_6_0_0_t1b_t1b),
    .I_7_0_0_t0b(n445_I_7_0_0_t0b),
    .I_7_0_0_t1b_t0b(n445_I_7_0_0_t1b_t0b),
    .I_7_0_0_t1b_t1b(n445_I_7_0_0_t1b_t1b),
    .I_8_0_0_t0b(n445_I_8_0_0_t0b),
    .I_8_0_0_t1b_t0b(n445_I_8_0_0_t1b_t0b),
    .I_8_0_0_t1b_t1b(n445_I_8_0_0_t1b_t1b),
    .I_9_0_0_t0b(n445_I_9_0_0_t0b),
    .I_9_0_0_t1b_t0b(n445_I_9_0_0_t1b_t0b),
    .I_9_0_0_t1b_t1b(n445_I_9_0_0_t1b_t1b),
    .I_10_0_0_t0b(n445_I_10_0_0_t0b),
    .I_10_0_0_t1b_t0b(n445_I_10_0_0_t1b_t0b),
    .I_10_0_0_t1b_t1b(n445_I_10_0_0_t1b_t1b),
    .I_11_0_0_t0b(n445_I_11_0_0_t0b),
    .I_11_0_0_t1b_t0b(n445_I_11_0_0_t1b_t0b),
    .I_11_0_0_t1b_t1b(n445_I_11_0_0_t1b_t1b),
    .I_12_0_0_t0b(n445_I_12_0_0_t0b),
    .I_12_0_0_t1b_t0b(n445_I_12_0_0_t1b_t0b),
    .I_12_0_0_t1b_t1b(n445_I_12_0_0_t1b_t1b),
    .I_13_0_0_t0b(n445_I_13_0_0_t0b),
    .I_13_0_0_t1b_t0b(n445_I_13_0_0_t1b_t0b),
    .I_13_0_0_t1b_t1b(n445_I_13_0_0_t1b_t1b),
    .I_14_0_0_t0b(n445_I_14_0_0_t0b),
    .I_14_0_0_t1b_t0b(n445_I_14_0_0_t1b_t0b),
    .I_14_0_0_t1b_t1b(n445_I_14_0_0_t1b_t1b),
    .I_15_0_0_t0b(n445_I_15_0_0_t0b),
    .I_15_0_0_t1b_t0b(n445_I_15_0_0_t1b_t0b),
    .I_15_0_0_t1b_t1b(n445_I_15_0_0_t1b_t1b),
    .O_0_0_t0b(n445_O_0_0_t0b),
    .O_0_0_t1b_t0b(n445_O_0_0_t1b_t0b),
    .O_0_0_t1b_t1b(n445_O_0_0_t1b_t1b),
    .O_1_0_t0b(n445_O_1_0_t0b),
    .O_1_0_t1b_t0b(n445_O_1_0_t1b_t0b),
    .O_1_0_t1b_t1b(n445_O_1_0_t1b_t1b),
    .O_2_0_t0b(n445_O_2_0_t0b),
    .O_2_0_t1b_t0b(n445_O_2_0_t1b_t0b),
    .O_2_0_t1b_t1b(n445_O_2_0_t1b_t1b),
    .O_3_0_t0b(n445_O_3_0_t0b),
    .O_3_0_t1b_t0b(n445_O_3_0_t1b_t0b),
    .O_3_0_t1b_t1b(n445_O_3_0_t1b_t1b),
    .O_4_0_t0b(n445_O_4_0_t0b),
    .O_4_0_t1b_t0b(n445_O_4_0_t1b_t0b),
    .O_4_0_t1b_t1b(n445_O_4_0_t1b_t1b),
    .O_5_0_t0b(n445_O_5_0_t0b),
    .O_5_0_t1b_t0b(n445_O_5_0_t1b_t0b),
    .O_5_0_t1b_t1b(n445_O_5_0_t1b_t1b),
    .O_6_0_t0b(n445_O_6_0_t0b),
    .O_6_0_t1b_t0b(n445_O_6_0_t1b_t0b),
    .O_6_0_t1b_t1b(n445_O_6_0_t1b_t1b),
    .O_7_0_t0b(n445_O_7_0_t0b),
    .O_7_0_t1b_t0b(n445_O_7_0_t1b_t0b),
    .O_7_0_t1b_t1b(n445_O_7_0_t1b_t1b),
    .O_8_0_t0b(n445_O_8_0_t0b),
    .O_8_0_t1b_t0b(n445_O_8_0_t1b_t0b),
    .O_8_0_t1b_t1b(n445_O_8_0_t1b_t1b),
    .O_9_0_t0b(n445_O_9_0_t0b),
    .O_9_0_t1b_t0b(n445_O_9_0_t1b_t0b),
    .O_9_0_t1b_t1b(n445_O_9_0_t1b_t1b),
    .O_10_0_t0b(n445_O_10_0_t0b),
    .O_10_0_t1b_t0b(n445_O_10_0_t1b_t0b),
    .O_10_0_t1b_t1b(n445_O_10_0_t1b_t1b),
    .O_11_0_t0b(n445_O_11_0_t0b),
    .O_11_0_t1b_t0b(n445_O_11_0_t1b_t0b),
    .O_11_0_t1b_t1b(n445_O_11_0_t1b_t1b),
    .O_12_0_t0b(n445_O_12_0_t0b),
    .O_12_0_t1b_t0b(n445_O_12_0_t1b_t0b),
    .O_12_0_t1b_t1b(n445_O_12_0_t1b_t1b),
    .O_13_0_t0b(n445_O_13_0_t0b),
    .O_13_0_t1b_t0b(n445_O_13_0_t1b_t0b),
    .O_13_0_t1b_t1b(n445_O_13_0_t1b_t1b),
    .O_14_0_t0b(n445_O_14_0_t0b),
    .O_14_0_t1b_t0b(n445_O_14_0_t1b_t0b),
    .O_14_0_t1b_t1b(n445_O_14_0_t1b_t1b),
    .O_15_0_t0b(n445_O_15_0_t0b),
    .O_15_0_t1b_t0b(n445_O_15_0_t1b_t0b),
    .O_15_0_t1b_t1b(n445_O_15_0_t1b_t1b)
  );
  Passthrough_3 n446 ( // @[Top.scala 452:22]
    .valid_up(n446_valid_up),
    .valid_down(n446_valid_down),
    .I_0_0_t0b(n446_I_0_0_t0b),
    .I_0_0_t1b_t0b(n446_I_0_0_t1b_t0b),
    .I_0_0_t1b_t1b(n446_I_0_0_t1b_t1b),
    .I_1_0_t0b(n446_I_1_0_t0b),
    .I_1_0_t1b_t0b(n446_I_1_0_t1b_t0b),
    .I_1_0_t1b_t1b(n446_I_1_0_t1b_t1b),
    .I_2_0_t0b(n446_I_2_0_t0b),
    .I_2_0_t1b_t0b(n446_I_2_0_t1b_t0b),
    .I_2_0_t1b_t1b(n446_I_2_0_t1b_t1b),
    .I_3_0_t0b(n446_I_3_0_t0b),
    .I_3_0_t1b_t0b(n446_I_3_0_t1b_t0b),
    .I_3_0_t1b_t1b(n446_I_3_0_t1b_t1b),
    .I_4_0_t0b(n446_I_4_0_t0b),
    .I_4_0_t1b_t0b(n446_I_4_0_t1b_t0b),
    .I_4_0_t1b_t1b(n446_I_4_0_t1b_t1b),
    .I_5_0_t0b(n446_I_5_0_t0b),
    .I_5_0_t1b_t0b(n446_I_5_0_t1b_t0b),
    .I_5_0_t1b_t1b(n446_I_5_0_t1b_t1b),
    .I_6_0_t0b(n446_I_6_0_t0b),
    .I_6_0_t1b_t0b(n446_I_6_0_t1b_t0b),
    .I_6_0_t1b_t1b(n446_I_6_0_t1b_t1b),
    .I_7_0_t0b(n446_I_7_0_t0b),
    .I_7_0_t1b_t0b(n446_I_7_0_t1b_t0b),
    .I_7_0_t1b_t1b(n446_I_7_0_t1b_t1b),
    .I_8_0_t0b(n446_I_8_0_t0b),
    .I_8_0_t1b_t0b(n446_I_8_0_t1b_t0b),
    .I_8_0_t1b_t1b(n446_I_8_0_t1b_t1b),
    .I_9_0_t0b(n446_I_9_0_t0b),
    .I_9_0_t1b_t0b(n446_I_9_0_t1b_t0b),
    .I_9_0_t1b_t1b(n446_I_9_0_t1b_t1b),
    .I_10_0_t0b(n446_I_10_0_t0b),
    .I_10_0_t1b_t0b(n446_I_10_0_t1b_t0b),
    .I_10_0_t1b_t1b(n446_I_10_0_t1b_t1b),
    .I_11_0_t0b(n446_I_11_0_t0b),
    .I_11_0_t1b_t0b(n446_I_11_0_t1b_t0b),
    .I_11_0_t1b_t1b(n446_I_11_0_t1b_t1b),
    .I_12_0_t0b(n446_I_12_0_t0b),
    .I_12_0_t1b_t0b(n446_I_12_0_t1b_t0b),
    .I_12_0_t1b_t1b(n446_I_12_0_t1b_t1b),
    .I_13_0_t0b(n446_I_13_0_t0b),
    .I_13_0_t1b_t0b(n446_I_13_0_t1b_t0b),
    .I_13_0_t1b_t1b(n446_I_13_0_t1b_t1b),
    .I_14_0_t0b(n446_I_14_0_t0b),
    .I_14_0_t1b_t0b(n446_I_14_0_t1b_t0b),
    .I_14_0_t1b_t1b(n446_I_14_0_t1b_t1b),
    .I_15_0_t0b(n446_I_15_0_t0b),
    .I_15_0_t1b_t0b(n446_I_15_0_t1b_t0b),
    .I_15_0_t1b_t1b(n446_I_15_0_t1b_t1b),
    .O_0_t0b(n446_O_0_t0b),
    .O_0_t1b_t0b(n446_O_0_t1b_t0b),
    .O_0_t1b_t1b(n446_O_0_t1b_t1b),
    .O_1_t0b(n446_O_1_t0b),
    .O_1_t1b_t0b(n446_O_1_t1b_t0b),
    .O_1_t1b_t1b(n446_O_1_t1b_t1b),
    .O_2_t0b(n446_O_2_t0b),
    .O_2_t1b_t0b(n446_O_2_t1b_t0b),
    .O_2_t1b_t1b(n446_O_2_t1b_t1b),
    .O_3_t0b(n446_O_3_t0b),
    .O_3_t1b_t0b(n446_O_3_t1b_t0b),
    .O_3_t1b_t1b(n446_O_3_t1b_t1b),
    .O_4_t0b(n446_O_4_t0b),
    .O_4_t1b_t0b(n446_O_4_t1b_t0b),
    .O_4_t1b_t1b(n446_O_4_t1b_t1b),
    .O_5_t0b(n446_O_5_t0b),
    .O_5_t1b_t0b(n446_O_5_t1b_t0b),
    .O_5_t1b_t1b(n446_O_5_t1b_t1b),
    .O_6_t0b(n446_O_6_t0b),
    .O_6_t1b_t0b(n446_O_6_t1b_t0b),
    .O_6_t1b_t1b(n446_O_6_t1b_t1b),
    .O_7_t0b(n446_O_7_t0b),
    .O_7_t1b_t0b(n446_O_7_t1b_t0b),
    .O_7_t1b_t1b(n446_O_7_t1b_t1b),
    .O_8_t0b(n446_O_8_t0b),
    .O_8_t1b_t0b(n446_O_8_t1b_t0b),
    .O_8_t1b_t1b(n446_O_8_t1b_t1b),
    .O_9_t0b(n446_O_9_t0b),
    .O_9_t1b_t0b(n446_O_9_t1b_t0b),
    .O_9_t1b_t1b(n446_O_9_t1b_t1b),
    .O_10_t0b(n446_O_10_t0b),
    .O_10_t1b_t0b(n446_O_10_t1b_t0b),
    .O_10_t1b_t1b(n446_O_10_t1b_t1b),
    .O_11_t0b(n446_O_11_t0b),
    .O_11_t1b_t0b(n446_O_11_t1b_t0b),
    .O_11_t1b_t1b(n446_O_11_t1b_t1b),
    .O_12_t0b(n446_O_12_t0b),
    .O_12_t1b_t0b(n446_O_12_t1b_t0b),
    .O_12_t1b_t1b(n446_O_12_t1b_t1b),
    .O_13_t0b(n446_O_13_t0b),
    .O_13_t1b_t0b(n446_O_13_t1b_t0b),
    .O_13_t1b_t1b(n446_O_13_t1b_t1b),
    .O_14_t0b(n446_O_14_t0b),
    .O_14_t1b_t0b(n446_O_14_t1b_t0b),
    .O_14_t1b_t1b(n446_O_14_t1b_t1b),
    .O_15_t0b(n446_O_15_t0b),
    .O_15_t1b_t0b(n446_O_15_t1b_t0b),
    .O_15_t1b_t1b(n446_O_15_t1b_t1b)
  );
  FIFO_9 n447 ( // @[Top.scala 455:22]
    .clock(n447_clock),
    .reset(n447_reset),
    .valid_up(n447_valid_up),
    .valid_down(n447_valid_down),
    .I_0_t0b(n447_I_0_t0b),
    .I_0_t1b_t0b(n447_I_0_t1b_t0b),
    .I_0_t1b_t1b(n447_I_0_t1b_t1b),
    .I_1_t0b(n447_I_1_t0b),
    .I_1_t1b_t0b(n447_I_1_t1b_t0b),
    .I_1_t1b_t1b(n447_I_1_t1b_t1b),
    .I_2_t0b(n447_I_2_t0b),
    .I_2_t1b_t0b(n447_I_2_t1b_t0b),
    .I_2_t1b_t1b(n447_I_2_t1b_t1b),
    .I_3_t0b(n447_I_3_t0b),
    .I_3_t1b_t0b(n447_I_3_t1b_t0b),
    .I_3_t1b_t1b(n447_I_3_t1b_t1b),
    .I_4_t0b(n447_I_4_t0b),
    .I_4_t1b_t0b(n447_I_4_t1b_t0b),
    .I_4_t1b_t1b(n447_I_4_t1b_t1b),
    .I_5_t0b(n447_I_5_t0b),
    .I_5_t1b_t0b(n447_I_5_t1b_t0b),
    .I_5_t1b_t1b(n447_I_5_t1b_t1b),
    .I_6_t0b(n447_I_6_t0b),
    .I_6_t1b_t0b(n447_I_6_t1b_t0b),
    .I_6_t1b_t1b(n447_I_6_t1b_t1b),
    .I_7_t0b(n447_I_7_t0b),
    .I_7_t1b_t0b(n447_I_7_t1b_t0b),
    .I_7_t1b_t1b(n447_I_7_t1b_t1b),
    .I_8_t0b(n447_I_8_t0b),
    .I_8_t1b_t0b(n447_I_8_t1b_t0b),
    .I_8_t1b_t1b(n447_I_8_t1b_t1b),
    .I_9_t0b(n447_I_9_t0b),
    .I_9_t1b_t0b(n447_I_9_t1b_t0b),
    .I_9_t1b_t1b(n447_I_9_t1b_t1b),
    .I_10_t0b(n447_I_10_t0b),
    .I_10_t1b_t0b(n447_I_10_t1b_t0b),
    .I_10_t1b_t1b(n447_I_10_t1b_t1b),
    .I_11_t0b(n447_I_11_t0b),
    .I_11_t1b_t0b(n447_I_11_t1b_t0b),
    .I_11_t1b_t1b(n447_I_11_t1b_t1b),
    .I_12_t0b(n447_I_12_t0b),
    .I_12_t1b_t0b(n447_I_12_t1b_t0b),
    .I_12_t1b_t1b(n447_I_12_t1b_t1b),
    .I_13_t0b(n447_I_13_t0b),
    .I_13_t1b_t0b(n447_I_13_t1b_t0b),
    .I_13_t1b_t1b(n447_I_13_t1b_t1b),
    .I_14_t0b(n447_I_14_t0b),
    .I_14_t1b_t0b(n447_I_14_t1b_t0b),
    .I_14_t1b_t1b(n447_I_14_t1b_t1b),
    .I_15_t0b(n447_I_15_t0b),
    .I_15_t1b_t0b(n447_I_15_t1b_t0b),
    .I_15_t1b_t1b(n447_I_15_t1b_t1b),
    .O_0_t0b(n447_O_0_t0b),
    .O_0_t1b_t0b(n447_O_0_t1b_t0b),
    .O_0_t1b_t1b(n447_O_0_t1b_t1b),
    .O_1_t0b(n447_O_1_t0b),
    .O_1_t1b_t0b(n447_O_1_t1b_t0b),
    .O_1_t1b_t1b(n447_O_1_t1b_t1b),
    .O_2_t0b(n447_O_2_t0b),
    .O_2_t1b_t0b(n447_O_2_t1b_t0b),
    .O_2_t1b_t1b(n447_O_2_t1b_t1b),
    .O_3_t0b(n447_O_3_t0b),
    .O_3_t1b_t0b(n447_O_3_t1b_t0b),
    .O_3_t1b_t1b(n447_O_3_t1b_t1b),
    .O_4_t0b(n447_O_4_t0b),
    .O_4_t1b_t0b(n447_O_4_t1b_t0b),
    .O_4_t1b_t1b(n447_O_4_t1b_t1b),
    .O_5_t0b(n447_O_5_t0b),
    .O_5_t1b_t0b(n447_O_5_t1b_t0b),
    .O_5_t1b_t1b(n447_O_5_t1b_t1b),
    .O_6_t0b(n447_O_6_t0b),
    .O_6_t1b_t0b(n447_O_6_t1b_t0b),
    .O_6_t1b_t1b(n447_O_6_t1b_t1b),
    .O_7_t0b(n447_O_7_t0b),
    .O_7_t1b_t0b(n447_O_7_t1b_t0b),
    .O_7_t1b_t1b(n447_O_7_t1b_t1b),
    .O_8_t0b(n447_O_8_t0b),
    .O_8_t1b_t0b(n447_O_8_t1b_t0b),
    .O_8_t1b_t1b(n447_O_8_t1b_t1b),
    .O_9_t0b(n447_O_9_t0b),
    .O_9_t1b_t0b(n447_O_9_t1b_t0b),
    .O_9_t1b_t1b(n447_O_9_t1b_t1b),
    .O_10_t0b(n447_O_10_t0b),
    .O_10_t1b_t0b(n447_O_10_t1b_t0b),
    .O_10_t1b_t1b(n447_O_10_t1b_t1b),
    .O_11_t0b(n447_O_11_t0b),
    .O_11_t1b_t0b(n447_O_11_t1b_t0b),
    .O_11_t1b_t1b(n447_O_11_t1b_t1b),
    .O_12_t0b(n447_O_12_t0b),
    .O_12_t1b_t0b(n447_O_12_t1b_t0b),
    .O_12_t1b_t1b(n447_O_12_t1b_t1b),
    .O_13_t0b(n447_O_13_t0b),
    .O_13_t1b_t0b(n447_O_13_t1b_t0b),
    .O_13_t1b_t1b(n447_O_13_t1b_t1b),
    .O_14_t0b(n447_O_14_t0b),
    .O_14_t1b_t0b(n447_O_14_t1b_t0b),
    .O_14_t1b_t1b(n447_O_14_t1b_t1b),
    .O_15_t0b(n447_O_15_t0b),
    .O_15_t1b_t0b(n447_O_15_t1b_t0b),
    .O_15_t1b_t1b(n447_O_15_t1b_t1b)
  );
  FIFO_9 n448 ( // @[Top.scala 458:22]
    .clock(n448_clock),
    .reset(n448_reset),
    .valid_up(n448_valid_up),
    .valid_down(n448_valid_down),
    .I_0_t0b(n448_I_0_t0b),
    .I_0_t1b_t0b(n448_I_0_t1b_t0b),
    .I_0_t1b_t1b(n448_I_0_t1b_t1b),
    .I_1_t0b(n448_I_1_t0b),
    .I_1_t1b_t0b(n448_I_1_t1b_t0b),
    .I_1_t1b_t1b(n448_I_1_t1b_t1b),
    .I_2_t0b(n448_I_2_t0b),
    .I_2_t1b_t0b(n448_I_2_t1b_t0b),
    .I_2_t1b_t1b(n448_I_2_t1b_t1b),
    .I_3_t0b(n448_I_3_t0b),
    .I_3_t1b_t0b(n448_I_3_t1b_t0b),
    .I_3_t1b_t1b(n448_I_3_t1b_t1b),
    .I_4_t0b(n448_I_4_t0b),
    .I_4_t1b_t0b(n448_I_4_t1b_t0b),
    .I_4_t1b_t1b(n448_I_4_t1b_t1b),
    .I_5_t0b(n448_I_5_t0b),
    .I_5_t1b_t0b(n448_I_5_t1b_t0b),
    .I_5_t1b_t1b(n448_I_5_t1b_t1b),
    .I_6_t0b(n448_I_6_t0b),
    .I_6_t1b_t0b(n448_I_6_t1b_t0b),
    .I_6_t1b_t1b(n448_I_6_t1b_t1b),
    .I_7_t0b(n448_I_7_t0b),
    .I_7_t1b_t0b(n448_I_7_t1b_t0b),
    .I_7_t1b_t1b(n448_I_7_t1b_t1b),
    .I_8_t0b(n448_I_8_t0b),
    .I_8_t1b_t0b(n448_I_8_t1b_t0b),
    .I_8_t1b_t1b(n448_I_8_t1b_t1b),
    .I_9_t0b(n448_I_9_t0b),
    .I_9_t1b_t0b(n448_I_9_t1b_t0b),
    .I_9_t1b_t1b(n448_I_9_t1b_t1b),
    .I_10_t0b(n448_I_10_t0b),
    .I_10_t1b_t0b(n448_I_10_t1b_t0b),
    .I_10_t1b_t1b(n448_I_10_t1b_t1b),
    .I_11_t0b(n448_I_11_t0b),
    .I_11_t1b_t0b(n448_I_11_t1b_t0b),
    .I_11_t1b_t1b(n448_I_11_t1b_t1b),
    .I_12_t0b(n448_I_12_t0b),
    .I_12_t1b_t0b(n448_I_12_t1b_t0b),
    .I_12_t1b_t1b(n448_I_12_t1b_t1b),
    .I_13_t0b(n448_I_13_t0b),
    .I_13_t1b_t0b(n448_I_13_t1b_t0b),
    .I_13_t1b_t1b(n448_I_13_t1b_t1b),
    .I_14_t0b(n448_I_14_t0b),
    .I_14_t1b_t0b(n448_I_14_t1b_t0b),
    .I_14_t1b_t1b(n448_I_14_t1b_t1b),
    .I_15_t0b(n448_I_15_t0b),
    .I_15_t1b_t0b(n448_I_15_t1b_t0b),
    .I_15_t1b_t1b(n448_I_15_t1b_t1b),
    .O_0_t0b(n448_O_0_t0b),
    .O_0_t1b_t0b(n448_O_0_t1b_t0b),
    .O_0_t1b_t1b(n448_O_0_t1b_t1b),
    .O_1_t0b(n448_O_1_t0b),
    .O_1_t1b_t0b(n448_O_1_t1b_t0b),
    .O_1_t1b_t1b(n448_O_1_t1b_t1b),
    .O_2_t0b(n448_O_2_t0b),
    .O_2_t1b_t0b(n448_O_2_t1b_t0b),
    .O_2_t1b_t1b(n448_O_2_t1b_t1b),
    .O_3_t0b(n448_O_3_t0b),
    .O_3_t1b_t0b(n448_O_3_t1b_t0b),
    .O_3_t1b_t1b(n448_O_3_t1b_t1b),
    .O_4_t0b(n448_O_4_t0b),
    .O_4_t1b_t0b(n448_O_4_t1b_t0b),
    .O_4_t1b_t1b(n448_O_4_t1b_t1b),
    .O_5_t0b(n448_O_5_t0b),
    .O_5_t1b_t0b(n448_O_5_t1b_t0b),
    .O_5_t1b_t1b(n448_O_5_t1b_t1b),
    .O_6_t0b(n448_O_6_t0b),
    .O_6_t1b_t0b(n448_O_6_t1b_t0b),
    .O_6_t1b_t1b(n448_O_6_t1b_t1b),
    .O_7_t0b(n448_O_7_t0b),
    .O_7_t1b_t0b(n448_O_7_t1b_t0b),
    .O_7_t1b_t1b(n448_O_7_t1b_t1b),
    .O_8_t0b(n448_O_8_t0b),
    .O_8_t1b_t0b(n448_O_8_t1b_t0b),
    .O_8_t1b_t1b(n448_O_8_t1b_t1b),
    .O_9_t0b(n448_O_9_t0b),
    .O_9_t1b_t0b(n448_O_9_t1b_t0b),
    .O_9_t1b_t1b(n448_O_9_t1b_t1b),
    .O_10_t0b(n448_O_10_t0b),
    .O_10_t1b_t0b(n448_O_10_t1b_t0b),
    .O_10_t1b_t1b(n448_O_10_t1b_t1b),
    .O_11_t0b(n448_O_11_t0b),
    .O_11_t1b_t0b(n448_O_11_t1b_t0b),
    .O_11_t1b_t1b(n448_O_11_t1b_t1b),
    .O_12_t0b(n448_O_12_t0b),
    .O_12_t1b_t0b(n448_O_12_t1b_t0b),
    .O_12_t1b_t1b(n448_O_12_t1b_t1b),
    .O_13_t0b(n448_O_13_t0b),
    .O_13_t1b_t0b(n448_O_13_t1b_t0b),
    .O_13_t1b_t1b(n448_O_13_t1b_t1b),
    .O_14_t0b(n448_O_14_t0b),
    .O_14_t1b_t0b(n448_O_14_t1b_t0b),
    .O_14_t1b_t1b(n448_O_14_t1b_t1b),
    .O_15_t0b(n448_O_15_t0b),
    .O_15_t1b_t0b(n448_O_15_t1b_t0b),
    .O_15_t1b_t1b(n448_O_15_t1b_t1b)
  );
  FIFO_9 n449 ( // @[Top.scala 461:22]
    .clock(n449_clock),
    .reset(n449_reset),
    .valid_up(n449_valid_up),
    .valid_down(n449_valid_down),
    .I_0_t0b(n449_I_0_t0b),
    .I_0_t1b_t0b(n449_I_0_t1b_t0b),
    .I_0_t1b_t1b(n449_I_0_t1b_t1b),
    .I_1_t0b(n449_I_1_t0b),
    .I_1_t1b_t0b(n449_I_1_t1b_t0b),
    .I_1_t1b_t1b(n449_I_1_t1b_t1b),
    .I_2_t0b(n449_I_2_t0b),
    .I_2_t1b_t0b(n449_I_2_t1b_t0b),
    .I_2_t1b_t1b(n449_I_2_t1b_t1b),
    .I_3_t0b(n449_I_3_t0b),
    .I_3_t1b_t0b(n449_I_3_t1b_t0b),
    .I_3_t1b_t1b(n449_I_3_t1b_t1b),
    .I_4_t0b(n449_I_4_t0b),
    .I_4_t1b_t0b(n449_I_4_t1b_t0b),
    .I_4_t1b_t1b(n449_I_4_t1b_t1b),
    .I_5_t0b(n449_I_5_t0b),
    .I_5_t1b_t0b(n449_I_5_t1b_t0b),
    .I_5_t1b_t1b(n449_I_5_t1b_t1b),
    .I_6_t0b(n449_I_6_t0b),
    .I_6_t1b_t0b(n449_I_6_t1b_t0b),
    .I_6_t1b_t1b(n449_I_6_t1b_t1b),
    .I_7_t0b(n449_I_7_t0b),
    .I_7_t1b_t0b(n449_I_7_t1b_t0b),
    .I_7_t1b_t1b(n449_I_7_t1b_t1b),
    .I_8_t0b(n449_I_8_t0b),
    .I_8_t1b_t0b(n449_I_8_t1b_t0b),
    .I_8_t1b_t1b(n449_I_8_t1b_t1b),
    .I_9_t0b(n449_I_9_t0b),
    .I_9_t1b_t0b(n449_I_9_t1b_t0b),
    .I_9_t1b_t1b(n449_I_9_t1b_t1b),
    .I_10_t0b(n449_I_10_t0b),
    .I_10_t1b_t0b(n449_I_10_t1b_t0b),
    .I_10_t1b_t1b(n449_I_10_t1b_t1b),
    .I_11_t0b(n449_I_11_t0b),
    .I_11_t1b_t0b(n449_I_11_t1b_t0b),
    .I_11_t1b_t1b(n449_I_11_t1b_t1b),
    .I_12_t0b(n449_I_12_t0b),
    .I_12_t1b_t0b(n449_I_12_t1b_t0b),
    .I_12_t1b_t1b(n449_I_12_t1b_t1b),
    .I_13_t0b(n449_I_13_t0b),
    .I_13_t1b_t0b(n449_I_13_t1b_t0b),
    .I_13_t1b_t1b(n449_I_13_t1b_t1b),
    .I_14_t0b(n449_I_14_t0b),
    .I_14_t1b_t0b(n449_I_14_t1b_t0b),
    .I_14_t1b_t1b(n449_I_14_t1b_t1b),
    .I_15_t0b(n449_I_15_t0b),
    .I_15_t1b_t0b(n449_I_15_t1b_t0b),
    .I_15_t1b_t1b(n449_I_15_t1b_t1b),
    .O_0_t0b(n449_O_0_t0b),
    .O_0_t1b_t0b(n449_O_0_t1b_t0b),
    .O_0_t1b_t1b(n449_O_0_t1b_t1b),
    .O_1_t0b(n449_O_1_t0b),
    .O_1_t1b_t0b(n449_O_1_t1b_t0b),
    .O_1_t1b_t1b(n449_O_1_t1b_t1b),
    .O_2_t0b(n449_O_2_t0b),
    .O_2_t1b_t0b(n449_O_2_t1b_t0b),
    .O_2_t1b_t1b(n449_O_2_t1b_t1b),
    .O_3_t0b(n449_O_3_t0b),
    .O_3_t1b_t0b(n449_O_3_t1b_t0b),
    .O_3_t1b_t1b(n449_O_3_t1b_t1b),
    .O_4_t0b(n449_O_4_t0b),
    .O_4_t1b_t0b(n449_O_4_t1b_t0b),
    .O_4_t1b_t1b(n449_O_4_t1b_t1b),
    .O_5_t0b(n449_O_5_t0b),
    .O_5_t1b_t0b(n449_O_5_t1b_t0b),
    .O_5_t1b_t1b(n449_O_5_t1b_t1b),
    .O_6_t0b(n449_O_6_t0b),
    .O_6_t1b_t0b(n449_O_6_t1b_t0b),
    .O_6_t1b_t1b(n449_O_6_t1b_t1b),
    .O_7_t0b(n449_O_7_t0b),
    .O_7_t1b_t0b(n449_O_7_t1b_t0b),
    .O_7_t1b_t1b(n449_O_7_t1b_t1b),
    .O_8_t0b(n449_O_8_t0b),
    .O_8_t1b_t0b(n449_O_8_t1b_t0b),
    .O_8_t1b_t1b(n449_O_8_t1b_t1b),
    .O_9_t0b(n449_O_9_t0b),
    .O_9_t1b_t0b(n449_O_9_t1b_t0b),
    .O_9_t1b_t1b(n449_O_9_t1b_t1b),
    .O_10_t0b(n449_O_10_t0b),
    .O_10_t1b_t0b(n449_O_10_t1b_t0b),
    .O_10_t1b_t1b(n449_O_10_t1b_t1b),
    .O_11_t0b(n449_O_11_t0b),
    .O_11_t1b_t0b(n449_O_11_t1b_t0b),
    .O_11_t1b_t1b(n449_O_11_t1b_t1b),
    .O_12_t0b(n449_O_12_t0b),
    .O_12_t1b_t0b(n449_O_12_t1b_t0b),
    .O_12_t1b_t1b(n449_O_12_t1b_t1b),
    .O_13_t0b(n449_O_13_t0b),
    .O_13_t1b_t0b(n449_O_13_t1b_t0b),
    .O_13_t1b_t1b(n449_O_13_t1b_t1b),
    .O_14_t0b(n449_O_14_t0b),
    .O_14_t1b_t0b(n449_O_14_t1b_t0b),
    .O_14_t1b_t1b(n449_O_14_t1b_t1b),
    .O_15_t0b(n449_O_15_t0b),
    .O_15_t1b_t0b(n449_O_15_t1b_t0b),
    .O_15_t1b_t1b(n449_O_15_t1b_t1b)
  );
  assign valid_down = n449_valid_down; // @[Top.scala 465:16]
  assign O_0_t0b = n449_O_0_t0b; // @[Top.scala 464:7]
  assign O_0_t1b_t0b = n449_O_0_t1b_t0b; // @[Top.scala 464:7]
  assign O_0_t1b_t1b = n449_O_0_t1b_t1b; // @[Top.scala 464:7]
  assign O_1_t0b = n449_O_1_t0b; // @[Top.scala 464:7]
  assign O_1_t1b_t0b = n449_O_1_t1b_t0b; // @[Top.scala 464:7]
  assign O_1_t1b_t1b = n449_O_1_t1b_t1b; // @[Top.scala 464:7]
  assign O_2_t0b = n449_O_2_t0b; // @[Top.scala 464:7]
  assign O_2_t1b_t0b = n449_O_2_t1b_t0b; // @[Top.scala 464:7]
  assign O_2_t1b_t1b = n449_O_2_t1b_t1b; // @[Top.scala 464:7]
  assign O_3_t0b = n449_O_3_t0b; // @[Top.scala 464:7]
  assign O_3_t1b_t0b = n449_O_3_t1b_t0b; // @[Top.scala 464:7]
  assign O_3_t1b_t1b = n449_O_3_t1b_t1b; // @[Top.scala 464:7]
  assign O_4_t0b = n449_O_4_t0b; // @[Top.scala 464:7]
  assign O_4_t1b_t0b = n449_O_4_t1b_t0b; // @[Top.scala 464:7]
  assign O_4_t1b_t1b = n449_O_4_t1b_t1b; // @[Top.scala 464:7]
  assign O_5_t0b = n449_O_5_t0b; // @[Top.scala 464:7]
  assign O_5_t1b_t0b = n449_O_5_t1b_t0b; // @[Top.scala 464:7]
  assign O_5_t1b_t1b = n449_O_5_t1b_t1b; // @[Top.scala 464:7]
  assign O_6_t0b = n449_O_6_t0b; // @[Top.scala 464:7]
  assign O_6_t1b_t0b = n449_O_6_t1b_t0b; // @[Top.scala 464:7]
  assign O_6_t1b_t1b = n449_O_6_t1b_t1b; // @[Top.scala 464:7]
  assign O_7_t0b = n449_O_7_t0b; // @[Top.scala 464:7]
  assign O_7_t1b_t0b = n449_O_7_t1b_t0b; // @[Top.scala 464:7]
  assign O_7_t1b_t1b = n449_O_7_t1b_t1b; // @[Top.scala 464:7]
  assign O_8_t0b = n449_O_8_t0b; // @[Top.scala 464:7]
  assign O_8_t1b_t0b = n449_O_8_t1b_t0b; // @[Top.scala 464:7]
  assign O_8_t1b_t1b = n449_O_8_t1b_t1b; // @[Top.scala 464:7]
  assign O_9_t0b = n449_O_9_t0b; // @[Top.scala 464:7]
  assign O_9_t1b_t0b = n449_O_9_t1b_t0b; // @[Top.scala 464:7]
  assign O_9_t1b_t1b = n449_O_9_t1b_t1b; // @[Top.scala 464:7]
  assign O_10_t0b = n449_O_10_t0b; // @[Top.scala 464:7]
  assign O_10_t1b_t0b = n449_O_10_t1b_t0b; // @[Top.scala 464:7]
  assign O_10_t1b_t1b = n449_O_10_t1b_t1b; // @[Top.scala 464:7]
  assign O_11_t0b = n449_O_11_t0b; // @[Top.scala 464:7]
  assign O_11_t1b_t0b = n449_O_11_t1b_t0b; // @[Top.scala 464:7]
  assign O_11_t1b_t1b = n449_O_11_t1b_t1b; // @[Top.scala 464:7]
  assign O_12_t0b = n449_O_12_t0b; // @[Top.scala 464:7]
  assign O_12_t1b_t0b = n449_O_12_t1b_t0b; // @[Top.scala 464:7]
  assign O_12_t1b_t1b = n449_O_12_t1b_t1b; // @[Top.scala 464:7]
  assign O_13_t0b = n449_O_13_t0b; // @[Top.scala 464:7]
  assign O_13_t1b_t0b = n449_O_13_t1b_t0b; // @[Top.scala 464:7]
  assign O_13_t1b_t1b = n449_O_13_t1b_t1b; // @[Top.scala 464:7]
  assign O_14_t0b = n449_O_14_t0b; // @[Top.scala 464:7]
  assign O_14_t1b_t0b = n449_O_14_t1b_t0b; // @[Top.scala 464:7]
  assign O_14_t1b_t1b = n449_O_14_t1b_t1b; // @[Top.scala 464:7]
  assign O_15_t0b = n449_O_15_t0b; // @[Top.scala 464:7]
  assign O_15_t1b_t0b = n449_O_15_t1b_t0b; // @[Top.scala 464:7]
  assign O_15_t1b_t1b = n449_O_15_t1b_t1b; // @[Top.scala 464:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 359:17]
  assign n1_I_0 = I_0; // @[Top.scala 358:10]
  assign n1_I_1 = I_1; // @[Top.scala 358:10]
  assign n1_I_2 = I_2; // @[Top.scala 358:10]
  assign n1_I_3 = I_3; // @[Top.scala 358:10]
  assign n1_I_4 = I_4; // @[Top.scala 358:10]
  assign n1_I_5 = I_5; // @[Top.scala 358:10]
  assign n1_I_6 = I_6; // @[Top.scala 358:10]
  assign n1_I_7 = I_7; // @[Top.scala 358:10]
  assign n1_I_8 = I_8; // @[Top.scala 358:10]
  assign n1_I_9 = I_9; // @[Top.scala 358:10]
  assign n1_I_10 = I_10; // @[Top.scala 358:10]
  assign n1_I_11 = I_11; // @[Top.scala 358:10]
  assign n1_I_12 = I_12; // @[Top.scala 358:10]
  assign n1_I_13 = I_13; // @[Top.scala 358:10]
  assign n1_I_14 = I_14; // @[Top.scala 358:10]
  assign n1_I_15 = I_15; // @[Top.scala 358:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 362:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 361:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 361:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 361:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 361:10]
  assign n2_I_4 = n1_O_4; // @[Top.scala 361:10]
  assign n2_I_5 = n1_O_5; // @[Top.scala 361:10]
  assign n2_I_6 = n1_O_6; // @[Top.scala 361:10]
  assign n2_I_7 = n1_O_7; // @[Top.scala 361:10]
  assign n2_I_8 = n1_O_8; // @[Top.scala 361:10]
  assign n2_I_9 = n1_O_9; // @[Top.scala 361:10]
  assign n2_I_10 = n1_O_10; // @[Top.scala 361:10]
  assign n2_I_11 = n1_O_11; // @[Top.scala 361:10]
  assign n2_I_12 = n1_O_12; // @[Top.scala 361:10]
  assign n2_I_13 = n1_O_13; // @[Top.scala 361:10]
  assign n2_I_14 = n1_O_14; // @[Top.scala 361:10]
  assign n2_I_15 = n1_O_15; // @[Top.scala 361:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 365:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 364:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 364:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 364:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 364:10]
  assign n3_I_4 = n2_O_4; // @[Top.scala 364:10]
  assign n3_I_5 = n2_O_5; // @[Top.scala 364:10]
  assign n3_I_6 = n2_O_6; // @[Top.scala 364:10]
  assign n3_I_7 = n2_O_7; // @[Top.scala 364:10]
  assign n3_I_8 = n2_O_8; // @[Top.scala 364:10]
  assign n3_I_9 = n2_O_9; // @[Top.scala 364:10]
  assign n3_I_10 = n2_O_10; // @[Top.scala 364:10]
  assign n3_I_11 = n2_O_11; // @[Top.scala 364:10]
  assign n3_I_12 = n2_O_12; // @[Top.scala 364:10]
  assign n3_I_13 = n2_O_13; // @[Top.scala 364:10]
  assign n3_I_14 = n2_O_14; // @[Top.scala 364:10]
  assign n3_I_15 = n2_O_15; // @[Top.scala 364:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 368:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 367:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 367:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 367:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 367:10]
  assign n4_I_4 = n3_O_4; // @[Top.scala 367:10]
  assign n4_I_5 = n3_O_5; // @[Top.scala 367:10]
  assign n4_I_6 = n3_O_6; // @[Top.scala 367:10]
  assign n4_I_7 = n3_O_7; // @[Top.scala 367:10]
  assign n4_I_8 = n3_O_8; // @[Top.scala 367:10]
  assign n4_I_9 = n3_O_9; // @[Top.scala 367:10]
  assign n4_I_10 = n3_O_10; // @[Top.scala 367:10]
  assign n4_I_11 = n3_O_11; // @[Top.scala 367:10]
  assign n4_I_12 = n3_O_12; // @[Top.scala 367:10]
  assign n4_I_13 = n3_O_13; // @[Top.scala 367:10]
  assign n4_I_14 = n3_O_14; // @[Top.scala 367:10]
  assign n4_I_15 = n3_O_15; // @[Top.scala 367:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 371:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 370:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 370:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 370:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 370:10]
  assign n5_I_4 = n4_O_4; // @[Top.scala 370:10]
  assign n5_I_5 = n4_O_5; // @[Top.scala 370:10]
  assign n5_I_6 = n4_O_6; // @[Top.scala 370:10]
  assign n5_I_7 = n4_O_7; // @[Top.scala 370:10]
  assign n5_I_8 = n4_O_8; // @[Top.scala 370:10]
  assign n5_I_9 = n4_O_9; // @[Top.scala 370:10]
  assign n5_I_10 = n4_O_10; // @[Top.scala 370:10]
  assign n5_I_11 = n4_O_11; // @[Top.scala 370:10]
  assign n5_I_12 = n4_O_12; // @[Top.scala 370:10]
  assign n5_I_13 = n4_O_13; // @[Top.scala 370:10]
  assign n5_I_14 = n4_O_14; // @[Top.scala 370:10]
  assign n5_I_15 = n4_O_15; // @[Top.scala 370:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 375:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 373:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 373:11]
  assign n6_I0_2 = n5_O_2; // @[Top.scala 373:11]
  assign n6_I0_3 = n5_O_3; // @[Top.scala 373:11]
  assign n6_I0_4 = n5_O_4; // @[Top.scala 373:11]
  assign n6_I0_5 = n5_O_5; // @[Top.scala 373:11]
  assign n6_I0_6 = n5_O_6; // @[Top.scala 373:11]
  assign n6_I0_7 = n5_O_7; // @[Top.scala 373:11]
  assign n6_I0_8 = n5_O_8; // @[Top.scala 373:11]
  assign n6_I0_9 = n5_O_9; // @[Top.scala 373:11]
  assign n6_I0_10 = n5_O_10; // @[Top.scala 373:11]
  assign n6_I0_11 = n5_O_11; // @[Top.scala 373:11]
  assign n6_I0_12 = n5_O_12; // @[Top.scala 373:11]
  assign n6_I0_13 = n5_O_13; // @[Top.scala 373:11]
  assign n6_I0_14 = n5_O_14; // @[Top.scala 373:11]
  assign n6_I0_15 = n5_O_15; // @[Top.scala 373:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 374:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 374:11]
  assign n6_I1_2 = n4_O_2; // @[Top.scala 374:11]
  assign n6_I1_3 = n4_O_3; // @[Top.scala 374:11]
  assign n6_I1_4 = n4_O_4; // @[Top.scala 374:11]
  assign n6_I1_5 = n4_O_5; // @[Top.scala 374:11]
  assign n6_I1_6 = n4_O_6; // @[Top.scala 374:11]
  assign n6_I1_7 = n4_O_7; // @[Top.scala 374:11]
  assign n6_I1_8 = n4_O_8; // @[Top.scala 374:11]
  assign n6_I1_9 = n4_O_9; // @[Top.scala 374:11]
  assign n6_I1_10 = n4_O_10; // @[Top.scala 374:11]
  assign n6_I1_11 = n4_O_11; // @[Top.scala 374:11]
  assign n6_I1_12 = n4_O_12; // @[Top.scala 374:11]
  assign n6_I1_13 = n4_O_13; // @[Top.scala 374:11]
  assign n6_I1_14 = n4_O_14; // @[Top.scala 374:11]
  assign n6_I1_15 = n4_O_15; // @[Top.scala 374:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 379:18]
  assign n13_I0_0_0 = n6_O_0_0; // @[Top.scala 377:12]
  assign n13_I0_0_1 = n6_O_0_1; // @[Top.scala 377:12]
  assign n13_I0_1_0 = n6_O_1_0; // @[Top.scala 377:12]
  assign n13_I0_1_1 = n6_O_1_1; // @[Top.scala 377:12]
  assign n13_I0_2_0 = n6_O_2_0; // @[Top.scala 377:12]
  assign n13_I0_2_1 = n6_O_2_1; // @[Top.scala 377:12]
  assign n13_I0_3_0 = n6_O_3_0; // @[Top.scala 377:12]
  assign n13_I0_3_1 = n6_O_3_1; // @[Top.scala 377:12]
  assign n13_I0_4_0 = n6_O_4_0; // @[Top.scala 377:12]
  assign n13_I0_4_1 = n6_O_4_1; // @[Top.scala 377:12]
  assign n13_I0_5_0 = n6_O_5_0; // @[Top.scala 377:12]
  assign n13_I0_5_1 = n6_O_5_1; // @[Top.scala 377:12]
  assign n13_I0_6_0 = n6_O_6_0; // @[Top.scala 377:12]
  assign n13_I0_6_1 = n6_O_6_1; // @[Top.scala 377:12]
  assign n13_I0_7_0 = n6_O_7_0; // @[Top.scala 377:12]
  assign n13_I0_7_1 = n6_O_7_1; // @[Top.scala 377:12]
  assign n13_I0_8_0 = n6_O_8_0; // @[Top.scala 377:12]
  assign n13_I0_8_1 = n6_O_8_1; // @[Top.scala 377:12]
  assign n13_I0_9_0 = n6_O_9_0; // @[Top.scala 377:12]
  assign n13_I0_9_1 = n6_O_9_1; // @[Top.scala 377:12]
  assign n13_I0_10_0 = n6_O_10_0; // @[Top.scala 377:12]
  assign n13_I0_10_1 = n6_O_10_1; // @[Top.scala 377:12]
  assign n13_I0_11_0 = n6_O_11_0; // @[Top.scala 377:12]
  assign n13_I0_11_1 = n6_O_11_1; // @[Top.scala 377:12]
  assign n13_I0_12_0 = n6_O_12_0; // @[Top.scala 377:12]
  assign n13_I0_12_1 = n6_O_12_1; // @[Top.scala 377:12]
  assign n13_I0_13_0 = n6_O_13_0; // @[Top.scala 377:12]
  assign n13_I0_13_1 = n6_O_13_1; // @[Top.scala 377:12]
  assign n13_I0_14_0 = n6_O_14_0; // @[Top.scala 377:12]
  assign n13_I0_14_1 = n6_O_14_1; // @[Top.scala 377:12]
  assign n13_I0_15_0 = n6_O_15_0; // @[Top.scala 377:12]
  assign n13_I0_15_1 = n6_O_15_1; // @[Top.scala 377:12]
  assign n13_I1_0 = n3_O_0; // @[Top.scala 378:12]
  assign n13_I1_1 = n3_O_1; // @[Top.scala 378:12]
  assign n13_I1_2 = n3_O_2; // @[Top.scala 378:12]
  assign n13_I1_3 = n3_O_3; // @[Top.scala 378:12]
  assign n13_I1_4 = n3_O_4; // @[Top.scala 378:12]
  assign n13_I1_5 = n3_O_5; // @[Top.scala 378:12]
  assign n13_I1_6 = n3_O_6; // @[Top.scala 378:12]
  assign n13_I1_7 = n3_O_7; // @[Top.scala 378:12]
  assign n13_I1_8 = n3_O_8; // @[Top.scala 378:12]
  assign n13_I1_9 = n3_O_9; // @[Top.scala 378:12]
  assign n13_I1_10 = n3_O_10; // @[Top.scala 378:12]
  assign n13_I1_11 = n3_O_11; // @[Top.scala 378:12]
  assign n13_I1_12 = n3_O_12; // @[Top.scala 378:12]
  assign n13_I1_13 = n3_O_13; // @[Top.scala 378:12]
  assign n13_I1_14 = n3_O_14; // @[Top.scala 378:12]
  assign n13_I1_15 = n3_O_15; // @[Top.scala 378:12]
  assign n22_valid_up = n13_valid_down; // @[Top.scala 382:18]
  assign n22_I_0_0 = n13_O_0_0; // @[Top.scala 381:11]
  assign n22_I_0_1 = n13_O_0_1; // @[Top.scala 381:11]
  assign n22_I_0_2 = n13_O_0_2; // @[Top.scala 381:11]
  assign n22_I_1_0 = n13_O_1_0; // @[Top.scala 381:11]
  assign n22_I_1_1 = n13_O_1_1; // @[Top.scala 381:11]
  assign n22_I_1_2 = n13_O_1_2; // @[Top.scala 381:11]
  assign n22_I_2_0 = n13_O_2_0; // @[Top.scala 381:11]
  assign n22_I_2_1 = n13_O_2_1; // @[Top.scala 381:11]
  assign n22_I_2_2 = n13_O_2_2; // @[Top.scala 381:11]
  assign n22_I_3_0 = n13_O_3_0; // @[Top.scala 381:11]
  assign n22_I_3_1 = n13_O_3_1; // @[Top.scala 381:11]
  assign n22_I_3_2 = n13_O_3_2; // @[Top.scala 381:11]
  assign n22_I_4_0 = n13_O_4_0; // @[Top.scala 381:11]
  assign n22_I_4_1 = n13_O_4_1; // @[Top.scala 381:11]
  assign n22_I_4_2 = n13_O_4_2; // @[Top.scala 381:11]
  assign n22_I_5_0 = n13_O_5_0; // @[Top.scala 381:11]
  assign n22_I_5_1 = n13_O_5_1; // @[Top.scala 381:11]
  assign n22_I_5_2 = n13_O_5_2; // @[Top.scala 381:11]
  assign n22_I_6_0 = n13_O_6_0; // @[Top.scala 381:11]
  assign n22_I_6_1 = n13_O_6_1; // @[Top.scala 381:11]
  assign n22_I_6_2 = n13_O_6_2; // @[Top.scala 381:11]
  assign n22_I_7_0 = n13_O_7_0; // @[Top.scala 381:11]
  assign n22_I_7_1 = n13_O_7_1; // @[Top.scala 381:11]
  assign n22_I_7_2 = n13_O_7_2; // @[Top.scala 381:11]
  assign n22_I_8_0 = n13_O_8_0; // @[Top.scala 381:11]
  assign n22_I_8_1 = n13_O_8_1; // @[Top.scala 381:11]
  assign n22_I_8_2 = n13_O_8_2; // @[Top.scala 381:11]
  assign n22_I_9_0 = n13_O_9_0; // @[Top.scala 381:11]
  assign n22_I_9_1 = n13_O_9_1; // @[Top.scala 381:11]
  assign n22_I_9_2 = n13_O_9_2; // @[Top.scala 381:11]
  assign n22_I_10_0 = n13_O_10_0; // @[Top.scala 381:11]
  assign n22_I_10_1 = n13_O_10_1; // @[Top.scala 381:11]
  assign n22_I_10_2 = n13_O_10_2; // @[Top.scala 381:11]
  assign n22_I_11_0 = n13_O_11_0; // @[Top.scala 381:11]
  assign n22_I_11_1 = n13_O_11_1; // @[Top.scala 381:11]
  assign n22_I_11_2 = n13_O_11_2; // @[Top.scala 381:11]
  assign n22_I_12_0 = n13_O_12_0; // @[Top.scala 381:11]
  assign n22_I_12_1 = n13_O_12_1; // @[Top.scala 381:11]
  assign n22_I_12_2 = n13_O_12_2; // @[Top.scala 381:11]
  assign n22_I_13_0 = n13_O_13_0; // @[Top.scala 381:11]
  assign n22_I_13_1 = n13_O_13_1; // @[Top.scala 381:11]
  assign n22_I_13_2 = n13_O_13_2; // @[Top.scala 381:11]
  assign n22_I_14_0 = n13_O_14_0; // @[Top.scala 381:11]
  assign n22_I_14_1 = n13_O_14_1; // @[Top.scala 381:11]
  assign n22_I_14_2 = n13_O_14_2; // @[Top.scala 381:11]
  assign n22_I_15_0 = n13_O_15_0; // @[Top.scala 381:11]
  assign n22_I_15_1 = n13_O_15_1; // @[Top.scala 381:11]
  assign n22_I_15_2 = n13_O_15_2; // @[Top.scala 381:11]
  assign n29_valid_up = n22_valid_down; // @[Top.scala 385:18]
  assign n29_I_0_0_0 = n22_O_0_0_0; // @[Top.scala 384:11]
  assign n29_I_0_0_1 = n22_O_0_0_1; // @[Top.scala 384:11]
  assign n29_I_0_0_2 = n22_O_0_0_2; // @[Top.scala 384:11]
  assign n29_I_1_0_0 = n22_O_1_0_0; // @[Top.scala 384:11]
  assign n29_I_1_0_1 = n22_O_1_0_1; // @[Top.scala 384:11]
  assign n29_I_1_0_2 = n22_O_1_0_2; // @[Top.scala 384:11]
  assign n29_I_2_0_0 = n22_O_2_0_0; // @[Top.scala 384:11]
  assign n29_I_2_0_1 = n22_O_2_0_1; // @[Top.scala 384:11]
  assign n29_I_2_0_2 = n22_O_2_0_2; // @[Top.scala 384:11]
  assign n29_I_3_0_0 = n22_O_3_0_0; // @[Top.scala 384:11]
  assign n29_I_3_0_1 = n22_O_3_0_1; // @[Top.scala 384:11]
  assign n29_I_3_0_2 = n22_O_3_0_2; // @[Top.scala 384:11]
  assign n29_I_4_0_0 = n22_O_4_0_0; // @[Top.scala 384:11]
  assign n29_I_4_0_1 = n22_O_4_0_1; // @[Top.scala 384:11]
  assign n29_I_4_0_2 = n22_O_4_0_2; // @[Top.scala 384:11]
  assign n29_I_5_0_0 = n22_O_5_0_0; // @[Top.scala 384:11]
  assign n29_I_5_0_1 = n22_O_5_0_1; // @[Top.scala 384:11]
  assign n29_I_5_0_2 = n22_O_5_0_2; // @[Top.scala 384:11]
  assign n29_I_6_0_0 = n22_O_6_0_0; // @[Top.scala 384:11]
  assign n29_I_6_0_1 = n22_O_6_0_1; // @[Top.scala 384:11]
  assign n29_I_6_0_2 = n22_O_6_0_2; // @[Top.scala 384:11]
  assign n29_I_7_0_0 = n22_O_7_0_0; // @[Top.scala 384:11]
  assign n29_I_7_0_1 = n22_O_7_0_1; // @[Top.scala 384:11]
  assign n29_I_7_0_2 = n22_O_7_0_2; // @[Top.scala 384:11]
  assign n29_I_8_0_0 = n22_O_8_0_0; // @[Top.scala 384:11]
  assign n29_I_8_0_1 = n22_O_8_0_1; // @[Top.scala 384:11]
  assign n29_I_8_0_2 = n22_O_8_0_2; // @[Top.scala 384:11]
  assign n29_I_9_0_0 = n22_O_9_0_0; // @[Top.scala 384:11]
  assign n29_I_9_0_1 = n22_O_9_0_1; // @[Top.scala 384:11]
  assign n29_I_9_0_2 = n22_O_9_0_2; // @[Top.scala 384:11]
  assign n29_I_10_0_0 = n22_O_10_0_0; // @[Top.scala 384:11]
  assign n29_I_10_0_1 = n22_O_10_0_1; // @[Top.scala 384:11]
  assign n29_I_10_0_2 = n22_O_10_0_2; // @[Top.scala 384:11]
  assign n29_I_11_0_0 = n22_O_11_0_0; // @[Top.scala 384:11]
  assign n29_I_11_0_1 = n22_O_11_0_1; // @[Top.scala 384:11]
  assign n29_I_11_0_2 = n22_O_11_0_2; // @[Top.scala 384:11]
  assign n29_I_12_0_0 = n22_O_12_0_0; // @[Top.scala 384:11]
  assign n29_I_12_0_1 = n22_O_12_0_1; // @[Top.scala 384:11]
  assign n29_I_12_0_2 = n22_O_12_0_2; // @[Top.scala 384:11]
  assign n29_I_13_0_0 = n22_O_13_0_0; // @[Top.scala 384:11]
  assign n29_I_13_0_1 = n22_O_13_0_1; // @[Top.scala 384:11]
  assign n29_I_13_0_2 = n22_O_13_0_2; // @[Top.scala 384:11]
  assign n29_I_14_0_0 = n22_O_14_0_0; // @[Top.scala 384:11]
  assign n29_I_14_0_1 = n22_O_14_0_1; // @[Top.scala 384:11]
  assign n29_I_14_0_2 = n22_O_14_0_2; // @[Top.scala 384:11]
  assign n29_I_15_0_0 = n22_O_15_0_0; // @[Top.scala 384:11]
  assign n29_I_15_0_1 = n22_O_15_0_1; // @[Top.scala 384:11]
  assign n29_I_15_0_2 = n22_O_15_0_2; // @[Top.scala 384:11]
  assign n30_clock = clock;
  assign n30_valid_up = n2_valid_down; // @[Top.scala 388:18]
  assign n30_I_0 = n2_O_0; // @[Top.scala 387:11]
  assign n30_I_1 = n2_O_1; // @[Top.scala 387:11]
  assign n30_I_2 = n2_O_2; // @[Top.scala 387:11]
  assign n30_I_3 = n2_O_3; // @[Top.scala 387:11]
  assign n30_I_4 = n2_O_4; // @[Top.scala 387:11]
  assign n30_I_5 = n2_O_5; // @[Top.scala 387:11]
  assign n30_I_6 = n2_O_6; // @[Top.scala 387:11]
  assign n30_I_7 = n2_O_7; // @[Top.scala 387:11]
  assign n30_I_8 = n2_O_8; // @[Top.scala 387:11]
  assign n30_I_9 = n2_O_9; // @[Top.scala 387:11]
  assign n30_I_10 = n2_O_10; // @[Top.scala 387:11]
  assign n30_I_11 = n2_O_11; // @[Top.scala 387:11]
  assign n30_I_12 = n2_O_12; // @[Top.scala 387:11]
  assign n30_I_13 = n2_O_13; // @[Top.scala 387:11]
  assign n30_I_14 = n2_O_14; // @[Top.scala 387:11]
  assign n30_I_15 = n2_O_15; // @[Top.scala 387:11]
  assign n31_clock = clock;
  assign n31_valid_up = n30_valid_down; // @[Top.scala 391:18]
  assign n31_I_0 = n30_O_0; // @[Top.scala 390:11]
  assign n31_I_1 = n30_O_1; // @[Top.scala 390:11]
  assign n31_I_2 = n30_O_2; // @[Top.scala 390:11]
  assign n31_I_3 = n30_O_3; // @[Top.scala 390:11]
  assign n31_I_4 = n30_O_4; // @[Top.scala 390:11]
  assign n31_I_5 = n30_O_5; // @[Top.scala 390:11]
  assign n31_I_6 = n30_O_6; // @[Top.scala 390:11]
  assign n31_I_7 = n30_O_7; // @[Top.scala 390:11]
  assign n31_I_8 = n30_O_8; // @[Top.scala 390:11]
  assign n31_I_9 = n30_O_9; // @[Top.scala 390:11]
  assign n31_I_10 = n30_O_10; // @[Top.scala 390:11]
  assign n31_I_11 = n30_O_11; // @[Top.scala 390:11]
  assign n31_I_12 = n30_O_12; // @[Top.scala 390:11]
  assign n31_I_13 = n30_O_13; // @[Top.scala 390:11]
  assign n31_I_14 = n30_O_14; // @[Top.scala 390:11]
  assign n31_I_15 = n30_O_15; // @[Top.scala 390:11]
  assign n32_valid_up = n31_valid_down & n30_valid_down; // @[Top.scala 395:18]
  assign n32_I0_0 = n31_O_0; // @[Top.scala 393:12]
  assign n32_I0_1 = n31_O_1; // @[Top.scala 393:12]
  assign n32_I0_2 = n31_O_2; // @[Top.scala 393:12]
  assign n32_I0_3 = n31_O_3; // @[Top.scala 393:12]
  assign n32_I0_4 = n31_O_4; // @[Top.scala 393:12]
  assign n32_I0_5 = n31_O_5; // @[Top.scala 393:12]
  assign n32_I0_6 = n31_O_6; // @[Top.scala 393:12]
  assign n32_I0_7 = n31_O_7; // @[Top.scala 393:12]
  assign n32_I0_8 = n31_O_8; // @[Top.scala 393:12]
  assign n32_I0_9 = n31_O_9; // @[Top.scala 393:12]
  assign n32_I0_10 = n31_O_10; // @[Top.scala 393:12]
  assign n32_I0_11 = n31_O_11; // @[Top.scala 393:12]
  assign n32_I0_12 = n31_O_12; // @[Top.scala 393:12]
  assign n32_I0_13 = n31_O_13; // @[Top.scala 393:12]
  assign n32_I0_14 = n31_O_14; // @[Top.scala 393:12]
  assign n32_I0_15 = n31_O_15; // @[Top.scala 393:12]
  assign n32_I1_0 = n30_O_0; // @[Top.scala 394:12]
  assign n32_I1_1 = n30_O_1; // @[Top.scala 394:12]
  assign n32_I1_2 = n30_O_2; // @[Top.scala 394:12]
  assign n32_I1_3 = n30_O_3; // @[Top.scala 394:12]
  assign n32_I1_4 = n30_O_4; // @[Top.scala 394:12]
  assign n32_I1_5 = n30_O_5; // @[Top.scala 394:12]
  assign n32_I1_6 = n30_O_6; // @[Top.scala 394:12]
  assign n32_I1_7 = n30_O_7; // @[Top.scala 394:12]
  assign n32_I1_8 = n30_O_8; // @[Top.scala 394:12]
  assign n32_I1_9 = n30_O_9; // @[Top.scala 394:12]
  assign n32_I1_10 = n30_O_10; // @[Top.scala 394:12]
  assign n32_I1_11 = n30_O_11; // @[Top.scala 394:12]
  assign n32_I1_12 = n30_O_12; // @[Top.scala 394:12]
  assign n32_I1_13 = n30_O_13; // @[Top.scala 394:12]
  assign n32_I1_14 = n30_O_14; // @[Top.scala 394:12]
  assign n32_I1_15 = n30_O_15; // @[Top.scala 394:12]
  assign n39_valid_up = n32_valid_down & n2_valid_down; // @[Top.scala 399:18]
  assign n39_I0_0_0 = n32_O_0_0; // @[Top.scala 397:12]
  assign n39_I0_0_1 = n32_O_0_1; // @[Top.scala 397:12]
  assign n39_I0_1_0 = n32_O_1_0; // @[Top.scala 397:12]
  assign n39_I0_1_1 = n32_O_1_1; // @[Top.scala 397:12]
  assign n39_I0_2_0 = n32_O_2_0; // @[Top.scala 397:12]
  assign n39_I0_2_1 = n32_O_2_1; // @[Top.scala 397:12]
  assign n39_I0_3_0 = n32_O_3_0; // @[Top.scala 397:12]
  assign n39_I0_3_1 = n32_O_3_1; // @[Top.scala 397:12]
  assign n39_I0_4_0 = n32_O_4_0; // @[Top.scala 397:12]
  assign n39_I0_4_1 = n32_O_4_1; // @[Top.scala 397:12]
  assign n39_I0_5_0 = n32_O_5_0; // @[Top.scala 397:12]
  assign n39_I0_5_1 = n32_O_5_1; // @[Top.scala 397:12]
  assign n39_I0_6_0 = n32_O_6_0; // @[Top.scala 397:12]
  assign n39_I0_6_1 = n32_O_6_1; // @[Top.scala 397:12]
  assign n39_I0_7_0 = n32_O_7_0; // @[Top.scala 397:12]
  assign n39_I0_7_1 = n32_O_7_1; // @[Top.scala 397:12]
  assign n39_I0_8_0 = n32_O_8_0; // @[Top.scala 397:12]
  assign n39_I0_8_1 = n32_O_8_1; // @[Top.scala 397:12]
  assign n39_I0_9_0 = n32_O_9_0; // @[Top.scala 397:12]
  assign n39_I0_9_1 = n32_O_9_1; // @[Top.scala 397:12]
  assign n39_I0_10_0 = n32_O_10_0; // @[Top.scala 397:12]
  assign n39_I0_10_1 = n32_O_10_1; // @[Top.scala 397:12]
  assign n39_I0_11_0 = n32_O_11_0; // @[Top.scala 397:12]
  assign n39_I0_11_1 = n32_O_11_1; // @[Top.scala 397:12]
  assign n39_I0_12_0 = n32_O_12_0; // @[Top.scala 397:12]
  assign n39_I0_12_1 = n32_O_12_1; // @[Top.scala 397:12]
  assign n39_I0_13_0 = n32_O_13_0; // @[Top.scala 397:12]
  assign n39_I0_13_1 = n32_O_13_1; // @[Top.scala 397:12]
  assign n39_I0_14_0 = n32_O_14_0; // @[Top.scala 397:12]
  assign n39_I0_14_1 = n32_O_14_1; // @[Top.scala 397:12]
  assign n39_I0_15_0 = n32_O_15_0; // @[Top.scala 397:12]
  assign n39_I0_15_1 = n32_O_15_1; // @[Top.scala 397:12]
  assign n39_I1_0 = n2_O_0; // @[Top.scala 398:12]
  assign n39_I1_1 = n2_O_1; // @[Top.scala 398:12]
  assign n39_I1_2 = n2_O_2; // @[Top.scala 398:12]
  assign n39_I1_3 = n2_O_3; // @[Top.scala 398:12]
  assign n39_I1_4 = n2_O_4; // @[Top.scala 398:12]
  assign n39_I1_5 = n2_O_5; // @[Top.scala 398:12]
  assign n39_I1_6 = n2_O_6; // @[Top.scala 398:12]
  assign n39_I1_7 = n2_O_7; // @[Top.scala 398:12]
  assign n39_I1_8 = n2_O_8; // @[Top.scala 398:12]
  assign n39_I1_9 = n2_O_9; // @[Top.scala 398:12]
  assign n39_I1_10 = n2_O_10; // @[Top.scala 398:12]
  assign n39_I1_11 = n2_O_11; // @[Top.scala 398:12]
  assign n39_I1_12 = n2_O_12; // @[Top.scala 398:12]
  assign n39_I1_13 = n2_O_13; // @[Top.scala 398:12]
  assign n39_I1_14 = n2_O_14; // @[Top.scala 398:12]
  assign n39_I1_15 = n2_O_15; // @[Top.scala 398:12]
  assign n48_valid_up = n39_valid_down; // @[Top.scala 402:18]
  assign n48_I_0_0 = n39_O_0_0; // @[Top.scala 401:11]
  assign n48_I_0_1 = n39_O_0_1; // @[Top.scala 401:11]
  assign n48_I_0_2 = n39_O_0_2; // @[Top.scala 401:11]
  assign n48_I_1_0 = n39_O_1_0; // @[Top.scala 401:11]
  assign n48_I_1_1 = n39_O_1_1; // @[Top.scala 401:11]
  assign n48_I_1_2 = n39_O_1_2; // @[Top.scala 401:11]
  assign n48_I_2_0 = n39_O_2_0; // @[Top.scala 401:11]
  assign n48_I_2_1 = n39_O_2_1; // @[Top.scala 401:11]
  assign n48_I_2_2 = n39_O_2_2; // @[Top.scala 401:11]
  assign n48_I_3_0 = n39_O_3_0; // @[Top.scala 401:11]
  assign n48_I_3_1 = n39_O_3_1; // @[Top.scala 401:11]
  assign n48_I_3_2 = n39_O_3_2; // @[Top.scala 401:11]
  assign n48_I_4_0 = n39_O_4_0; // @[Top.scala 401:11]
  assign n48_I_4_1 = n39_O_4_1; // @[Top.scala 401:11]
  assign n48_I_4_2 = n39_O_4_2; // @[Top.scala 401:11]
  assign n48_I_5_0 = n39_O_5_0; // @[Top.scala 401:11]
  assign n48_I_5_1 = n39_O_5_1; // @[Top.scala 401:11]
  assign n48_I_5_2 = n39_O_5_2; // @[Top.scala 401:11]
  assign n48_I_6_0 = n39_O_6_0; // @[Top.scala 401:11]
  assign n48_I_6_1 = n39_O_6_1; // @[Top.scala 401:11]
  assign n48_I_6_2 = n39_O_6_2; // @[Top.scala 401:11]
  assign n48_I_7_0 = n39_O_7_0; // @[Top.scala 401:11]
  assign n48_I_7_1 = n39_O_7_1; // @[Top.scala 401:11]
  assign n48_I_7_2 = n39_O_7_2; // @[Top.scala 401:11]
  assign n48_I_8_0 = n39_O_8_0; // @[Top.scala 401:11]
  assign n48_I_8_1 = n39_O_8_1; // @[Top.scala 401:11]
  assign n48_I_8_2 = n39_O_8_2; // @[Top.scala 401:11]
  assign n48_I_9_0 = n39_O_9_0; // @[Top.scala 401:11]
  assign n48_I_9_1 = n39_O_9_1; // @[Top.scala 401:11]
  assign n48_I_9_2 = n39_O_9_2; // @[Top.scala 401:11]
  assign n48_I_10_0 = n39_O_10_0; // @[Top.scala 401:11]
  assign n48_I_10_1 = n39_O_10_1; // @[Top.scala 401:11]
  assign n48_I_10_2 = n39_O_10_2; // @[Top.scala 401:11]
  assign n48_I_11_0 = n39_O_11_0; // @[Top.scala 401:11]
  assign n48_I_11_1 = n39_O_11_1; // @[Top.scala 401:11]
  assign n48_I_11_2 = n39_O_11_2; // @[Top.scala 401:11]
  assign n48_I_12_0 = n39_O_12_0; // @[Top.scala 401:11]
  assign n48_I_12_1 = n39_O_12_1; // @[Top.scala 401:11]
  assign n48_I_12_2 = n39_O_12_2; // @[Top.scala 401:11]
  assign n48_I_13_0 = n39_O_13_0; // @[Top.scala 401:11]
  assign n48_I_13_1 = n39_O_13_1; // @[Top.scala 401:11]
  assign n48_I_13_2 = n39_O_13_2; // @[Top.scala 401:11]
  assign n48_I_14_0 = n39_O_14_0; // @[Top.scala 401:11]
  assign n48_I_14_1 = n39_O_14_1; // @[Top.scala 401:11]
  assign n48_I_14_2 = n39_O_14_2; // @[Top.scala 401:11]
  assign n48_I_15_0 = n39_O_15_0; // @[Top.scala 401:11]
  assign n48_I_15_1 = n39_O_15_1; // @[Top.scala 401:11]
  assign n48_I_15_2 = n39_O_15_2; // @[Top.scala 401:11]
  assign n55_valid_up = n48_valid_down; // @[Top.scala 405:18]
  assign n55_I_0_0_0 = n48_O_0_0_0; // @[Top.scala 404:11]
  assign n55_I_0_0_1 = n48_O_0_0_1; // @[Top.scala 404:11]
  assign n55_I_0_0_2 = n48_O_0_0_2; // @[Top.scala 404:11]
  assign n55_I_1_0_0 = n48_O_1_0_0; // @[Top.scala 404:11]
  assign n55_I_1_0_1 = n48_O_1_0_1; // @[Top.scala 404:11]
  assign n55_I_1_0_2 = n48_O_1_0_2; // @[Top.scala 404:11]
  assign n55_I_2_0_0 = n48_O_2_0_0; // @[Top.scala 404:11]
  assign n55_I_2_0_1 = n48_O_2_0_1; // @[Top.scala 404:11]
  assign n55_I_2_0_2 = n48_O_2_0_2; // @[Top.scala 404:11]
  assign n55_I_3_0_0 = n48_O_3_0_0; // @[Top.scala 404:11]
  assign n55_I_3_0_1 = n48_O_3_0_1; // @[Top.scala 404:11]
  assign n55_I_3_0_2 = n48_O_3_0_2; // @[Top.scala 404:11]
  assign n55_I_4_0_0 = n48_O_4_0_0; // @[Top.scala 404:11]
  assign n55_I_4_0_1 = n48_O_4_0_1; // @[Top.scala 404:11]
  assign n55_I_4_0_2 = n48_O_4_0_2; // @[Top.scala 404:11]
  assign n55_I_5_0_0 = n48_O_5_0_0; // @[Top.scala 404:11]
  assign n55_I_5_0_1 = n48_O_5_0_1; // @[Top.scala 404:11]
  assign n55_I_5_0_2 = n48_O_5_0_2; // @[Top.scala 404:11]
  assign n55_I_6_0_0 = n48_O_6_0_0; // @[Top.scala 404:11]
  assign n55_I_6_0_1 = n48_O_6_0_1; // @[Top.scala 404:11]
  assign n55_I_6_0_2 = n48_O_6_0_2; // @[Top.scala 404:11]
  assign n55_I_7_0_0 = n48_O_7_0_0; // @[Top.scala 404:11]
  assign n55_I_7_0_1 = n48_O_7_0_1; // @[Top.scala 404:11]
  assign n55_I_7_0_2 = n48_O_7_0_2; // @[Top.scala 404:11]
  assign n55_I_8_0_0 = n48_O_8_0_0; // @[Top.scala 404:11]
  assign n55_I_8_0_1 = n48_O_8_0_1; // @[Top.scala 404:11]
  assign n55_I_8_0_2 = n48_O_8_0_2; // @[Top.scala 404:11]
  assign n55_I_9_0_0 = n48_O_9_0_0; // @[Top.scala 404:11]
  assign n55_I_9_0_1 = n48_O_9_0_1; // @[Top.scala 404:11]
  assign n55_I_9_0_2 = n48_O_9_0_2; // @[Top.scala 404:11]
  assign n55_I_10_0_0 = n48_O_10_0_0; // @[Top.scala 404:11]
  assign n55_I_10_0_1 = n48_O_10_0_1; // @[Top.scala 404:11]
  assign n55_I_10_0_2 = n48_O_10_0_2; // @[Top.scala 404:11]
  assign n55_I_11_0_0 = n48_O_11_0_0; // @[Top.scala 404:11]
  assign n55_I_11_0_1 = n48_O_11_0_1; // @[Top.scala 404:11]
  assign n55_I_11_0_2 = n48_O_11_0_2; // @[Top.scala 404:11]
  assign n55_I_12_0_0 = n48_O_12_0_0; // @[Top.scala 404:11]
  assign n55_I_12_0_1 = n48_O_12_0_1; // @[Top.scala 404:11]
  assign n55_I_12_0_2 = n48_O_12_0_2; // @[Top.scala 404:11]
  assign n55_I_13_0_0 = n48_O_13_0_0; // @[Top.scala 404:11]
  assign n55_I_13_0_1 = n48_O_13_0_1; // @[Top.scala 404:11]
  assign n55_I_13_0_2 = n48_O_13_0_2; // @[Top.scala 404:11]
  assign n55_I_14_0_0 = n48_O_14_0_0; // @[Top.scala 404:11]
  assign n55_I_14_0_1 = n48_O_14_0_1; // @[Top.scala 404:11]
  assign n55_I_14_0_2 = n48_O_14_0_2; // @[Top.scala 404:11]
  assign n55_I_15_0_0 = n48_O_15_0_0; // @[Top.scala 404:11]
  assign n55_I_15_0_1 = n48_O_15_0_1; // @[Top.scala 404:11]
  assign n55_I_15_0_2 = n48_O_15_0_2; // @[Top.scala 404:11]
  assign n56_valid_up = n29_valid_down & n55_valid_down; // @[Top.scala 409:18]
  assign n56_I0_0_0 = n29_O_0_0; // @[Top.scala 407:12]
  assign n56_I0_0_1 = n29_O_0_1; // @[Top.scala 407:12]
  assign n56_I0_0_2 = n29_O_0_2; // @[Top.scala 407:12]
  assign n56_I0_1_0 = n29_O_1_0; // @[Top.scala 407:12]
  assign n56_I0_1_1 = n29_O_1_1; // @[Top.scala 407:12]
  assign n56_I0_1_2 = n29_O_1_2; // @[Top.scala 407:12]
  assign n56_I0_2_0 = n29_O_2_0; // @[Top.scala 407:12]
  assign n56_I0_2_1 = n29_O_2_1; // @[Top.scala 407:12]
  assign n56_I0_2_2 = n29_O_2_2; // @[Top.scala 407:12]
  assign n56_I0_3_0 = n29_O_3_0; // @[Top.scala 407:12]
  assign n56_I0_3_1 = n29_O_3_1; // @[Top.scala 407:12]
  assign n56_I0_3_2 = n29_O_3_2; // @[Top.scala 407:12]
  assign n56_I0_4_0 = n29_O_4_0; // @[Top.scala 407:12]
  assign n56_I0_4_1 = n29_O_4_1; // @[Top.scala 407:12]
  assign n56_I0_4_2 = n29_O_4_2; // @[Top.scala 407:12]
  assign n56_I0_5_0 = n29_O_5_0; // @[Top.scala 407:12]
  assign n56_I0_5_1 = n29_O_5_1; // @[Top.scala 407:12]
  assign n56_I0_5_2 = n29_O_5_2; // @[Top.scala 407:12]
  assign n56_I0_6_0 = n29_O_6_0; // @[Top.scala 407:12]
  assign n56_I0_6_1 = n29_O_6_1; // @[Top.scala 407:12]
  assign n56_I0_6_2 = n29_O_6_2; // @[Top.scala 407:12]
  assign n56_I0_7_0 = n29_O_7_0; // @[Top.scala 407:12]
  assign n56_I0_7_1 = n29_O_7_1; // @[Top.scala 407:12]
  assign n56_I0_7_2 = n29_O_7_2; // @[Top.scala 407:12]
  assign n56_I0_8_0 = n29_O_8_0; // @[Top.scala 407:12]
  assign n56_I0_8_1 = n29_O_8_1; // @[Top.scala 407:12]
  assign n56_I0_8_2 = n29_O_8_2; // @[Top.scala 407:12]
  assign n56_I0_9_0 = n29_O_9_0; // @[Top.scala 407:12]
  assign n56_I0_9_1 = n29_O_9_1; // @[Top.scala 407:12]
  assign n56_I0_9_2 = n29_O_9_2; // @[Top.scala 407:12]
  assign n56_I0_10_0 = n29_O_10_0; // @[Top.scala 407:12]
  assign n56_I0_10_1 = n29_O_10_1; // @[Top.scala 407:12]
  assign n56_I0_10_2 = n29_O_10_2; // @[Top.scala 407:12]
  assign n56_I0_11_0 = n29_O_11_0; // @[Top.scala 407:12]
  assign n56_I0_11_1 = n29_O_11_1; // @[Top.scala 407:12]
  assign n56_I0_11_2 = n29_O_11_2; // @[Top.scala 407:12]
  assign n56_I0_12_0 = n29_O_12_0; // @[Top.scala 407:12]
  assign n56_I0_12_1 = n29_O_12_1; // @[Top.scala 407:12]
  assign n56_I0_12_2 = n29_O_12_2; // @[Top.scala 407:12]
  assign n56_I0_13_0 = n29_O_13_0; // @[Top.scala 407:12]
  assign n56_I0_13_1 = n29_O_13_1; // @[Top.scala 407:12]
  assign n56_I0_13_2 = n29_O_13_2; // @[Top.scala 407:12]
  assign n56_I0_14_0 = n29_O_14_0; // @[Top.scala 407:12]
  assign n56_I0_14_1 = n29_O_14_1; // @[Top.scala 407:12]
  assign n56_I0_14_2 = n29_O_14_2; // @[Top.scala 407:12]
  assign n56_I0_15_0 = n29_O_15_0; // @[Top.scala 407:12]
  assign n56_I0_15_1 = n29_O_15_1; // @[Top.scala 407:12]
  assign n56_I0_15_2 = n29_O_15_2; // @[Top.scala 407:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 408:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 408:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 408:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 408:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 408:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 408:12]
  assign n56_I1_2_0 = n55_O_2_0; // @[Top.scala 408:12]
  assign n56_I1_2_1 = n55_O_2_1; // @[Top.scala 408:12]
  assign n56_I1_2_2 = n55_O_2_2; // @[Top.scala 408:12]
  assign n56_I1_3_0 = n55_O_3_0; // @[Top.scala 408:12]
  assign n56_I1_3_1 = n55_O_3_1; // @[Top.scala 408:12]
  assign n56_I1_3_2 = n55_O_3_2; // @[Top.scala 408:12]
  assign n56_I1_4_0 = n55_O_4_0; // @[Top.scala 408:12]
  assign n56_I1_4_1 = n55_O_4_1; // @[Top.scala 408:12]
  assign n56_I1_4_2 = n55_O_4_2; // @[Top.scala 408:12]
  assign n56_I1_5_0 = n55_O_5_0; // @[Top.scala 408:12]
  assign n56_I1_5_1 = n55_O_5_1; // @[Top.scala 408:12]
  assign n56_I1_5_2 = n55_O_5_2; // @[Top.scala 408:12]
  assign n56_I1_6_0 = n55_O_6_0; // @[Top.scala 408:12]
  assign n56_I1_6_1 = n55_O_6_1; // @[Top.scala 408:12]
  assign n56_I1_6_2 = n55_O_6_2; // @[Top.scala 408:12]
  assign n56_I1_7_0 = n55_O_7_0; // @[Top.scala 408:12]
  assign n56_I1_7_1 = n55_O_7_1; // @[Top.scala 408:12]
  assign n56_I1_7_2 = n55_O_7_2; // @[Top.scala 408:12]
  assign n56_I1_8_0 = n55_O_8_0; // @[Top.scala 408:12]
  assign n56_I1_8_1 = n55_O_8_1; // @[Top.scala 408:12]
  assign n56_I1_8_2 = n55_O_8_2; // @[Top.scala 408:12]
  assign n56_I1_9_0 = n55_O_9_0; // @[Top.scala 408:12]
  assign n56_I1_9_1 = n55_O_9_1; // @[Top.scala 408:12]
  assign n56_I1_9_2 = n55_O_9_2; // @[Top.scala 408:12]
  assign n56_I1_10_0 = n55_O_10_0; // @[Top.scala 408:12]
  assign n56_I1_10_1 = n55_O_10_1; // @[Top.scala 408:12]
  assign n56_I1_10_2 = n55_O_10_2; // @[Top.scala 408:12]
  assign n56_I1_11_0 = n55_O_11_0; // @[Top.scala 408:12]
  assign n56_I1_11_1 = n55_O_11_1; // @[Top.scala 408:12]
  assign n56_I1_11_2 = n55_O_11_2; // @[Top.scala 408:12]
  assign n56_I1_12_0 = n55_O_12_0; // @[Top.scala 408:12]
  assign n56_I1_12_1 = n55_O_12_1; // @[Top.scala 408:12]
  assign n56_I1_12_2 = n55_O_12_2; // @[Top.scala 408:12]
  assign n56_I1_13_0 = n55_O_13_0; // @[Top.scala 408:12]
  assign n56_I1_13_1 = n55_O_13_1; // @[Top.scala 408:12]
  assign n56_I1_13_2 = n55_O_13_2; // @[Top.scala 408:12]
  assign n56_I1_14_0 = n55_O_14_0; // @[Top.scala 408:12]
  assign n56_I1_14_1 = n55_O_14_1; // @[Top.scala 408:12]
  assign n56_I1_14_2 = n55_O_14_2; // @[Top.scala 408:12]
  assign n56_I1_15_0 = n55_O_15_0; // @[Top.scala 408:12]
  assign n56_I1_15_1 = n55_O_15_1; // @[Top.scala 408:12]
  assign n56_I1_15_2 = n55_O_15_2; // @[Top.scala 408:12]
  assign n63_clock = clock;
  assign n63_valid_up = n1_valid_down; // @[Top.scala 412:18]
  assign n63_I_0 = n1_O_0; // @[Top.scala 411:11]
  assign n63_I_1 = n1_O_1; // @[Top.scala 411:11]
  assign n63_I_2 = n1_O_2; // @[Top.scala 411:11]
  assign n63_I_3 = n1_O_3; // @[Top.scala 411:11]
  assign n63_I_4 = n1_O_4; // @[Top.scala 411:11]
  assign n63_I_5 = n1_O_5; // @[Top.scala 411:11]
  assign n63_I_6 = n1_O_6; // @[Top.scala 411:11]
  assign n63_I_7 = n1_O_7; // @[Top.scala 411:11]
  assign n63_I_8 = n1_O_8; // @[Top.scala 411:11]
  assign n63_I_9 = n1_O_9; // @[Top.scala 411:11]
  assign n63_I_10 = n1_O_10; // @[Top.scala 411:11]
  assign n63_I_11 = n1_O_11; // @[Top.scala 411:11]
  assign n63_I_12 = n1_O_12; // @[Top.scala 411:11]
  assign n63_I_13 = n1_O_13; // @[Top.scala 411:11]
  assign n63_I_14 = n1_O_14; // @[Top.scala 411:11]
  assign n63_I_15 = n1_O_15; // @[Top.scala 411:11]
  assign n64_clock = clock;
  assign n64_valid_up = n63_valid_down; // @[Top.scala 415:18]
  assign n64_I_0 = n63_O_0; // @[Top.scala 414:11]
  assign n64_I_1 = n63_O_1; // @[Top.scala 414:11]
  assign n64_I_2 = n63_O_2; // @[Top.scala 414:11]
  assign n64_I_3 = n63_O_3; // @[Top.scala 414:11]
  assign n64_I_4 = n63_O_4; // @[Top.scala 414:11]
  assign n64_I_5 = n63_O_5; // @[Top.scala 414:11]
  assign n64_I_6 = n63_O_6; // @[Top.scala 414:11]
  assign n64_I_7 = n63_O_7; // @[Top.scala 414:11]
  assign n64_I_8 = n63_O_8; // @[Top.scala 414:11]
  assign n64_I_9 = n63_O_9; // @[Top.scala 414:11]
  assign n64_I_10 = n63_O_10; // @[Top.scala 414:11]
  assign n64_I_11 = n63_O_11; // @[Top.scala 414:11]
  assign n64_I_12 = n63_O_12; // @[Top.scala 414:11]
  assign n64_I_13 = n63_O_13; // @[Top.scala 414:11]
  assign n64_I_14 = n63_O_14; // @[Top.scala 414:11]
  assign n64_I_15 = n63_O_15; // @[Top.scala 414:11]
  assign n65_valid_up = n64_valid_down & n63_valid_down; // @[Top.scala 419:18]
  assign n65_I0_0 = n64_O_0; // @[Top.scala 417:12]
  assign n65_I0_1 = n64_O_1; // @[Top.scala 417:12]
  assign n65_I0_2 = n64_O_2; // @[Top.scala 417:12]
  assign n65_I0_3 = n64_O_3; // @[Top.scala 417:12]
  assign n65_I0_4 = n64_O_4; // @[Top.scala 417:12]
  assign n65_I0_5 = n64_O_5; // @[Top.scala 417:12]
  assign n65_I0_6 = n64_O_6; // @[Top.scala 417:12]
  assign n65_I0_7 = n64_O_7; // @[Top.scala 417:12]
  assign n65_I0_8 = n64_O_8; // @[Top.scala 417:12]
  assign n65_I0_9 = n64_O_9; // @[Top.scala 417:12]
  assign n65_I0_10 = n64_O_10; // @[Top.scala 417:12]
  assign n65_I0_11 = n64_O_11; // @[Top.scala 417:12]
  assign n65_I0_12 = n64_O_12; // @[Top.scala 417:12]
  assign n65_I0_13 = n64_O_13; // @[Top.scala 417:12]
  assign n65_I0_14 = n64_O_14; // @[Top.scala 417:12]
  assign n65_I0_15 = n64_O_15; // @[Top.scala 417:12]
  assign n65_I1_0 = n63_O_0; // @[Top.scala 418:12]
  assign n65_I1_1 = n63_O_1; // @[Top.scala 418:12]
  assign n65_I1_2 = n63_O_2; // @[Top.scala 418:12]
  assign n65_I1_3 = n63_O_3; // @[Top.scala 418:12]
  assign n65_I1_4 = n63_O_4; // @[Top.scala 418:12]
  assign n65_I1_5 = n63_O_5; // @[Top.scala 418:12]
  assign n65_I1_6 = n63_O_6; // @[Top.scala 418:12]
  assign n65_I1_7 = n63_O_7; // @[Top.scala 418:12]
  assign n65_I1_8 = n63_O_8; // @[Top.scala 418:12]
  assign n65_I1_9 = n63_O_9; // @[Top.scala 418:12]
  assign n65_I1_10 = n63_O_10; // @[Top.scala 418:12]
  assign n65_I1_11 = n63_O_11; // @[Top.scala 418:12]
  assign n65_I1_12 = n63_O_12; // @[Top.scala 418:12]
  assign n65_I1_13 = n63_O_13; // @[Top.scala 418:12]
  assign n65_I1_14 = n63_O_14; // @[Top.scala 418:12]
  assign n65_I1_15 = n63_O_15; // @[Top.scala 418:12]
  assign n72_valid_up = n65_valid_down & n1_valid_down; // @[Top.scala 423:18]
  assign n72_I0_0_0 = n65_O_0_0; // @[Top.scala 421:12]
  assign n72_I0_0_1 = n65_O_0_1; // @[Top.scala 421:12]
  assign n72_I0_1_0 = n65_O_1_0; // @[Top.scala 421:12]
  assign n72_I0_1_1 = n65_O_1_1; // @[Top.scala 421:12]
  assign n72_I0_2_0 = n65_O_2_0; // @[Top.scala 421:12]
  assign n72_I0_2_1 = n65_O_2_1; // @[Top.scala 421:12]
  assign n72_I0_3_0 = n65_O_3_0; // @[Top.scala 421:12]
  assign n72_I0_3_1 = n65_O_3_1; // @[Top.scala 421:12]
  assign n72_I0_4_0 = n65_O_4_0; // @[Top.scala 421:12]
  assign n72_I0_4_1 = n65_O_4_1; // @[Top.scala 421:12]
  assign n72_I0_5_0 = n65_O_5_0; // @[Top.scala 421:12]
  assign n72_I0_5_1 = n65_O_5_1; // @[Top.scala 421:12]
  assign n72_I0_6_0 = n65_O_6_0; // @[Top.scala 421:12]
  assign n72_I0_6_1 = n65_O_6_1; // @[Top.scala 421:12]
  assign n72_I0_7_0 = n65_O_7_0; // @[Top.scala 421:12]
  assign n72_I0_7_1 = n65_O_7_1; // @[Top.scala 421:12]
  assign n72_I0_8_0 = n65_O_8_0; // @[Top.scala 421:12]
  assign n72_I0_8_1 = n65_O_8_1; // @[Top.scala 421:12]
  assign n72_I0_9_0 = n65_O_9_0; // @[Top.scala 421:12]
  assign n72_I0_9_1 = n65_O_9_1; // @[Top.scala 421:12]
  assign n72_I0_10_0 = n65_O_10_0; // @[Top.scala 421:12]
  assign n72_I0_10_1 = n65_O_10_1; // @[Top.scala 421:12]
  assign n72_I0_11_0 = n65_O_11_0; // @[Top.scala 421:12]
  assign n72_I0_11_1 = n65_O_11_1; // @[Top.scala 421:12]
  assign n72_I0_12_0 = n65_O_12_0; // @[Top.scala 421:12]
  assign n72_I0_12_1 = n65_O_12_1; // @[Top.scala 421:12]
  assign n72_I0_13_0 = n65_O_13_0; // @[Top.scala 421:12]
  assign n72_I0_13_1 = n65_O_13_1; // @[Top.scala 421:12]
  assign n72_I0_14_0 = n65_O_14_0; // @[Top.scala 421:12]
  assign n72_I0_14_1 = n65_O_14_1; // @[Top.scala 421:12]
  assign n72_I0_15_0 = n65_O_15_0; // @[Top.scala 421:12]
  assign n72_I0_15_1 = n65_O_15_1; // @[Top.scala 421:12]
  assign n72_I1_0 = n1_O_0; // @[Top.scala 422:12]
  assign n72_I1_1 = n1_O_1; // @[Top.scala 422:12]
  assign n72_I1_2 = n1_O_2; // @[Top.scala 422:12]
  assign n72_I1_3 = n1_O_3; // @[Top.scala 422:12]
  assign n72_I1_4 = n1_O_4; // @[Top.scala 422:12]
  assign n72_I1_5 = n1_O_5; // @[Top.scala 422:12]
  assign n72_I1_6 = n1_O_6; // @[Top.scala 422:12]
  assign n72_I1_7 = n1_O_7; // @[Top.scala 422:12]
  assign n72_I1_8 = n1_O_8; // @[Top.scala 422:12]
  assign n72_I1_9 = n1_O_9; // @[Top.scala 422:12]
  assign n72_I1_10 = n1_O_10; // @[Top.scala 422:12]
  assign n72_I1_11 = n1_O_11; // @[Top.scala 422:12]
  assign n72_I1_12 = n1_O_12; // @[Top.scala 422:12]
  assign n72_I1_13 = n1_O_13; // @[Top.scala 422:12]
  assign n72_I1_14 = n1_O_14; // @[Top.scala 422:12]
  assign n72_I1_15 = n1_O_15; // @[Top.scala 422:12]
  assign n81_valid_up = n72_valid_down; // @[Top.scala 426:18]
  assign n81_I_0_0 = n72_O_0_0; // @[Top.scala 425:11]
  assign n81_I_0_1 = n72_O_0_1; // @[Top.scala 425:11]
  assign n81_I_0_2 = n72_O_0_2; // @[Top.scala 425:11]
  assign n81_I_1_0 = n72_O_1_0; // @[Top.scala 425:11]
  assign n81_I_1_1 = n72_O_1_1; // @[Top.scala 425:11]
  assign n81_I_1_2 = n72_O_1_2; // @[Top.scala 425:11]
  assign n81_I_2_0 = n72_O_2_0; // @[Top.scala 425:11]
  assign n81_I_2_1 = n72_O_2_1; // @[Top.scala 425:11]
  assign n81_I_2_2 = n72_O_2_2; // @[Top.scala 425:11]
  assign n81_I_3_0 = n72_O_3_0; // @[Top.scala 425:11]
  assign n81_I_3_1 = n72_O_3_1; // @[Top.scala 425:11]
  assign n81_I_3_2 = n72_O_3_2; // @[Top.scala 425:11]
  assign n81_I_4_0 = n72_O_4_0; // @[Top.scala 425:11]
  assign n81_I_4_1 = n72_O_4_1; // @[Top.scala 425:11]
  assign n81_I_4_2 = n72_O_4_2; // @[Top.scala 425:11]
  assign n81_I_5_0 = n72_O_5_0; // @[Top.scala 425:11]
  assign n81_I_5_1 = n72_O_5_1; // @[Top.scala 425:11]
  assign n81_I_5_2 = n72_O_5_2; // @[Top.scala 425:11]
  assign n81_I_6_0 = n72_O_6_0; // @[Top.scala 425:11]
  assign n81_I_6_1 = n72_O_6_1; // @[Top.scala 425:11]
  assign n81_I_6_2 = n72_O_6_2; // @[Top.scala 425:11]
  assign n81_I_7_0 = n72_O_7_0; // @[Top.scala 425:11]
  assign n81_I_7_1 = n72_O_7_1; // @[Top.scala 425:11]
  assign n81_I_7_2 = n72_O_7_2; // @[Top.scala 425:11]
  assign n81_I_8_0 = n72_O_8_0; // @[Top.scala 425:11]
  assign n81_I_8_1 = n72_O_8_1; // @[Top.scala 425:11]
  assign n81_I_8_2 = n72_O_8_2; // @[Top.scala 425:11]
  assign n81_I_9_0 = n72_O_9_0; // @[Top.scala 425:11]
  assign n81_I_9_1 = n72_O_9_1; // @[Top.scala 425:11]
  assign n81_I_9_2 = n72_O_9_2; // @[Top.scala 425:11]
  assign n81_I_10_0 = n72_O_10_0; // @[Top.scala 425:11]
  assign n81_I_10_1 = n72_O_10_1; // @[Top.scala 425:11]
  assign n81_I_10_2 = n72_O_10_2; // @[Top.scala 425:11]
  assign n81_I_11_0 = n72_O_11_0; // @[Top.scala 425:11]
  assign n81_I_11_1 = n72_O_11_1; // @[Top.scala 425:11]
  assign n81_I_11_2 = n72_O_11_2; // @[Top.scala 425:11]
  assign n81_I_12_0 = n72_O_12_0; // @[Top.scala 425:11]
  assign n81_I_12_1 = n72_O_12_1; // @[Top.scala 425:11]
  assign n81_I_12_2 = n72_O_12_2; // @[Top.scala 425:11]
  assign n81_I_13_0 = n72_O_13_0; // @[Top.scala 425:11]
  assign n81_I_13_1 = n72_O_13_1; // @[Top.scala 425:11]
  assign n81_I_13_2 = n72_O_13_2; // @[Top.scala 425:11]
  assign n81_I_14_0 = n72_O_14_0; // @[Top.scala 425:11]
  assign n81_I_14_1 = n72_O_14_1; // @[Top.scala 425:11]
  assign n81_I_14_2 = n72_O_14_2; // @[Top.scala 425:11]
  assign n81_I_15_0 = n72_O_15_0; // @[Top.scala 425:11]
  assign n81_I_15_1 = n72_O_15_1; // @[Top.scala 425:11]
  assign n81_I_15_2 = n72_O_15_2; // @[Top.scala 425:11]
  assign n88_valid_up = n81_valid_down; // @[Top.scala 429:18]
  assign n88_I_0_0_0 = n81_O_0_0_0; // @[Top.scala 428:11]
  assign n88_I_0_0_1 = n81_O_0_0_1; // @[Top.scala 428:11]
  assign n88_I_0_0_2 = n81_O_0_0_2; // @[Top.scala 428:11]
  assign n88_I_1_0_0 = n81_O_1_0_0; // @[Top.scala 428:11]
  assign n88_I_1_0_1 = n81_O_1_0_1; // @[Top.scala 428:11]
  assign n88_I_1_0_2 = n81_O_1_0_2; // @[Top.scala 428:11]
  assign n88_I_2_0_0 = n81_O_2_0_0; // @[Top.scala 428:11]
  assign n88_I_2_0_1 = n81_O_2_0_1; // @[Top.scala 428:11]
  assign n88_I_2_0_2 = n81_O_2_0_2; // @[Top.scala 428:11]
  assign n88_I_3_0_0 = n81_O_3_0_0; // @[Top.scala 428:11]
  assign n88_I_3_0_1 = n81_O_3_0_1; // @[Top.scala 428:11]
  assign n88_I_3_0_2 = n81_O_3_0_2; // @[Top.scala 428:11]
  assign n88_I_4_0_0 = n81_O_4_0_0; // @[Top.scala 428:11]
  assign n88_I_4_0_1 = n81_O_4_0_1; // @[Top.scala 428:11]
  assign n88_I_4_0_2 = n81_O_4_0_2; // @[Top.scala 428:11]
  assign n88_I_5_0_0 = n81_O_5_0_0; // @[Top.scala 428:11]
  assign n88_I_5_0_1 = n81_O_5_0_1; // @[Top.scala 428:11]
  assign n88_I_5_0_2 = n81_O_5_0_2; // @[Top.scala 428:11]
  assign n88_I_6_0_0 = n81_O_6_0_0; // @[Top.scala 428:11]
  assign n88_I_6_0_1 = n81_O_6_0_1; // @[Top.scala 428:11]
  assign n88_I_6_0_2 = n81_O_6_0_2; // @[Top.scala 428:11]
  assign n88_I_7_0_0 = n81_O_7_0_0; // @[Top.scala 428:11]
  assign n88_I_7_0_1 = n81_O_7_0_1; // @[Top.scala 428:11]
  assign n88_I_7_0_2 = n81_O_7_0_2; // @[Top.scala 428:11]
  assign n88_I_8_0_0 = n81_O_8_0_0; // @[Top.scala 428:11]
  assign n88_I_8_0_1 = n81_O_8_0_1; // @[Top.scala 428:11]
  assign n88_I_8_0_2 = n81_O_8_0_2; // @[Top.scala 428:11]
  assign n88_I_9_0_0 = n81_O_9_0_0; // @[Top.scala 428:11]
  assign n88_I_9_0_1 = n81_O_9_0_1; // @[Top.scala 428:11]
  assign n88_I_9_0_2 = n81_O_9_0_2; // @[Top.scala 428:11]
  assign n88_I_10_0_0 = n81_O_10_0_0; // @[Top.scala 428:11]
  assign n88_I_10_0_1 = n81_O_10_0_1; // @[Top.scala 428:11]
  assign n88_I_10_0_2 = n81_O_10_0_2; // @[Top.scala 428:11]
  assign n88_I_11_0_0 = n81_O_11_0_0; // @[Top.scala 428:11]
  assign n88_I_11_0_1 = n81_O_11_0_1; // @[Top.scala 428:11]
  assign n88_I_11_0_2 = n81_O_11_0_2; // @[Top.scala 428:11]
  assign n88_I_12_0_0 = n81_O_12_0_0; // @[Top.scala 428:11]
  assign n88_I_12_0_1 = n81_O_12_0_1; // @[Top.scala 428:11]
  assign n88_I_12_0_2 = n81_O_12_0_2; // @[Top.scala 428:11]
  assign n88_I_13_0_0 = n81_O_13_0_0; // @[Top.scala 428:11]
  assign n88_I_13_0_1 = n81_O_13_0_1; // @[Top.scala 428:11]
  assign n88_I_13_0_2 = n81_O_13_0_2; // @[Top.scala 428:11]
  assign n88_I_14_0_0 = n81_O_14_0_0; // @[Top.scala 428:11]
  assign n88_I_14_0_1 = n81_O_14_0_1; // @[Top.scala 428:11]
  assign n88_I_14_0_2 = n81_O_14_0_2; // @[Top.scala 428:11]
  assign n88_I_15_0_0 = n81_O_15_0_0; // @[Top.scala 428:11]
  assign n88_I_15_0_1 = n81_O_15_0_1; // @[Top.scala 428:11]
  assign n88_I_15_0_2 = n81_O_15_0_2; // @[Top.scala 428:11]
  assign n89_valid_up = n56_valid_down & n88_valid_down; // @[Top.scala 433:18]
  assign n89_I0_0_0_0 = n56_O_0_0_0; // @[Top.scala 431:12]
  assign n89_I0_0_0_1 = n56_O_0_0_1; // @[Top.scala 431:12]
  assign n89_I0_0_0_2 = n56_O_0_0_2; // @[Top.scala 431:12]
  assign n89_I0_0_1_0 = n56_O_0_1_0; // @[Top.scala 431:12]
  assign n89_I0_0_1_1 = n56_O_0_1_1; // @[Top.scala 431:12]
  assign n89_I0_0_1_2 = n56_O_0_1_2; // @[Top.scala 431:12]
  assign n89_I0_1_0_0 = n56_O_1_0_0; // @[Top.scala 431:12]
  assign n89_I0_1_0_1 = n56_O_1_0_1; // @[Top.scala 431:12]
  assign n89_I0_1_0_2 = n56_O_1_0_2; // @[Top.scala 431:12]
  assign n89_I0_1_1_0 = n56_O_1_1_0; // @[Top.scala 431:12]
  assign n89_I0_1_1_1 = n56_O_1_1_1; // @[Top.scala 431:12]
  assign n89_I0_1_1_2 = n56_O_1_1_2; // @[Top.scala 431:12]
  assign n89_I0_2_0_0 = n56_O_2_0_0; // @[Top.scala 431:12]
  assign n89_I0_2_0_1 = n56_O_2_0_1; // @[Top.scala 431:12]
  assign n89_I0_2_0_2 = n56_O_2_0_2; // @[Top.scala 431:12]
  assign n89_I0_2_1_0 = n56_O_2_1_0; // @[Top.scala 431:12]
  assign n89_I0_2_1_1 = n56_O_2_1_1; // @[Top.scala 431:12]
  assign n89_I0_2_1_2 = n56_O_2_1_2; // @[Top.scala 431:12]
  assign n89_I0_3_0_0 = n56_O_3_0_0; // @[Top.scala 431:12]
  assign n89_I0_3_0_1 = n56_O_3_0_1; // @[Top.scala 431:12]
  assign n89_I0_3_0_2 = n56_O_3_0_2; // @[Top.scala 431:12]
  assign n89_I0_3_1_0 = n56_O_3_1_0; // @[Top.scala 431:12]
  assign n89_I0_3_1_1 = n56_O_3_1_1; // @[Top.scala 431:12]
  assign n89_I0_3_1_2 = n56_O_3_1_2; // @[Top.scala 431:12]
  assign n89_I0_4_0_0 = n56_O_4_0_0; // @[Top.scala 431:12]
  assign n89_I0_4_0_1 = n56_O_4_0_1; // @[Top.scala 431:12]
  assign n89_I0_4_0_2 = n56_O_4_0_2; // @[Top.scala 431:12]
  assign n89_I0_4_1_0 = n56_O_4_1_0; // @[Top.scala 431:12]
  assign n89_I0_4_1_1 = n56_O_4_1_1; // @[Top.scala 431:12]
  assign n89_I0_4_1_2 = n56_O_4_1_2; // @[Top.scala 431:12]
  assign n89_I0_5_0_0 = n56_O_5_0_0; // @[Top.scala 431:12]
  assign n89_I0_5_0_1 = n56_O_5_0_1; // @[Top.scala 431:12]
  assign n89_I0_5_0_2 = n56_O_5_0_2; // @[Top.scala 431:12]
  assign n89_I0_5_1_0 = n56_O_5_1_0; // @[Top.scala 431:12]
  assign n89_I0_5_1_1 = n56_O_5_1_1; // @[Top.scala 431:12]
  assign n89_I0_5_1_2 = n56_O_5_1_2; // @[Top.scala 431:12]
  assign n89_I0_6_0_0 = n56_O_6_0_0; // @[Top.scala 431:12]
  assign n89_I0_6_0_1 = n56_O_6_0_1; // @[Top.scala 431:12]
  assign n89_I0_6_0_2 = n56_O_6_0_2; // @[Top.scala 431:12]
  assign n89_I0_6_1_0 = n56_O_6_1_0; // @[Top.scala 431:12]
  assign n89_I0_6_1_1 = n56_O_6_1_1; // @[Top.scala 431:12]
  assign n89_I0_6_1_2 = n56_O_6_1_2; // @[Top.scala 431:12]
  assign n89_I0_7_0_0 = n56_O_7_0_0; // @[Top.scala 431:12]
  assign n89_I0_7_0_1 = n56_O_7_0_1; // @[Top.scala 431:12]
  assign n89_I0_7_0_2 = n56_O_7_0_2; // @[Top.scala 431:12]
  assign n89_I0_7_1_0 = n56_O_7_1_0; // @[Top.scala 431:12]
  assign n89_I0_7_1_1 = n56_O_7_1_1; // @[Top.scala 431:12]
  assign n89_I0_7_1_2 = n56_O_7_1_2; // @[Top.scala 431:12]
  assign n89_I0_8_0_0 = n56_O_8_0_0; // @[Top.scala 431:12]
  assign n89_I0_8_0_1 = n56_O_8_0_1; // @[Top.scala 431:12]
  assign n89_I0_8_0_2 = n56_O_8_0_2; // @[Top.scala 431:12]
  assign n89_I0_8_1_0 = n56_O_8_1_0; // @[Top.scala 431:12]
  assign n89_I0_8_1_1 = n56_O_8_1_1; // @[Top.scala 431:12]
  assign n89_I0_8_1_2 = n56_O_8_1_2; // @[Top.scala 431:12]
  assign n89_I0_9_0_0 = n56_O_9_0_0; // @[Top.scala 431:12]
  assign n89_I0_9_0_1 = n56_O_9_0_1; // @[Top.scala 431:12]
  assign n89_I0_9_0_2 = n56_O_9_0_2; // @[Top.scala 431:12]
  assign n89_I0_9_1_0 = n56_O_9_1_0; // @[Top.scala 431:12]
  assign n89_I0_9_1_1 = n56_O_9_1_1; // @[Top.scala 431:12]
  assign n89_I0_9_1_2 = n56_O_9_1_2; // @[Top.scala 431:12]
  assign n89_I0_10_0_0 = n56_O_10_0_0; // @[Top.scala 431:12]
  assign n89_I0_10_0_1 = n56_O_10_0_1; // @[Top.scala 431:12]
  assign n89_I0_10_0_2 = n56_O_10_0_2; // @[Top.scala 431:12]
  assign n89_I0_10_1_0 = n56_O_10_1_0; // @[Top.scala 431:12]
  assign n89_I0_10_1_1 = n56_O_10_1_1; // @[Top.scala 431:12]
  assign n89_I0_10_1_2 = n56_O_10_1_2; // @[Top.scala 431:12]
  assign n89_I0_11_0_0 = n56_O_11_0_0; // @[Top.scala 431:12]
  assign n89_I0_11_0_1 = n56_O_11_0_1; // @[Top.scala 431:12]
  assign n89_I0_11_0_2 = n56_O_11_0_2; // @[Top.scala 431:12]
  assign n89_I0_11_1_0 = n56_O_11_1_0; // @[Top.scala 431:12]
  assign n89_I0_11_1_1 = n56_O_11_1_1; // @[Top.scala 431:12]
  assign n89_I0_11_1_2 = n56_O_11_1_2; // @[Top.scala 431:12]
  assign n89_I0_12_0_0 = n56_O_12_0_0; // @[Top.scala 431:12]
  assign n89_I0_12_0_1 = n56_O_12_0_1; // @[Top.scala 431:12]
  assign n89_I0_12_0_2 = n56_O_12_0_2; // @[Top.scala 431:12]
  assign n89_I0_12_1_0 = n56_O_12_1_0; // @[Top.scala 431:12]
  assign n89_I0_12_1_1 = n56_O_12_1_1; // @[Top.scala 431:12]
  assign n89_I0_12_1_2 = n56_O_12_1_2; // @[Top.scala 431:12]
  assign n89_I0_13_0_0 = n56_O_13_0_0; // @[Top.scala 431:12]
  assign n89_I0_13_0_1 = n56_O_13_0_1; // @[Top.scala 431:12]
  assign n89_I0_13_0_2 = n56_O_13_0_2; // @[Top.scala 431:12]
  assign n89_I0_13_1_0 = n56_O_13_1_0; // @[Top.scala 431:12]
  assign n89_I0_13_1_1 = n56_O_13_1_1; // @[Top.scala 431:12]
  assign n89_I0_13_1_2 = n56_O_13_1_2; // @[Top.scala 431:12]
  assign n89_I0_14_0_0 = n56_O_14_0_0; // @[Top.scala 431:12]
  assign n89_I0_14_0_1 = n56_O_14_0_1; // @[Top.scala 431:12]
  assign n89_I0_14_0_2 = n56_O_14_0_2; // @[Top.scala 431:12]
  assign n89_I0_14_1_0 = n56_O_14_1_0; // @[Top.scala 431:12]
  assign n89_I0_14_1_1 = n56_O_14_1_1; // @[Top.scala 431:12]
  assign n89_I0_14_1_2 = n56_O_14_1_2; // @[Top.scala 431:12]
  assign n89_I0_15_0_0 = n56_O_15_0_0; // @[Top.scala 431:12]
  assign n89_I0_15_0_1 = n56_O_15_0_1; // @[Top.scala 431:12]
  assign n89_I0_15_0_2 = n56_O_15_0_2; // @[Top.scala 431:12]
  assign n89_I0_15_1_0 = n56_O_15_1_0; // @[Top.scala 431:12]
  assign n89_I0_15_1_1 = n56_O_15_1_1; // @[Top.scala 431:12]
  assign n89_I0_15_1_2 = n56_O_15_1_2; // @[Top.scala 431:12]
  assign n89_I1_0_0 = n88_O_0_0; // @[Top.scala 432:12]
  assign n89_I1_0_1 = n88_O_0_1; // @[Top.scala 432:12]
  assign n89_I1_0_2 = n88_O_0_2; // @[Top.scala 432:12]
  assign n89_I1_1_0 = n88_O_1_0; // @[Top.scala 432:12]
  assign n89_I1_1_1 = n88_O_1_1; // @[Top.scala 432:12]
  assign n89_I1_1_2 = n88_O_1_2; // @[Top.scala 432:12]
  assign n89_I1_2_0 = n88_O_2_0; // @[Top.scala 432:12]
  assign n89_I1_2_1 = n88_O_2_1; // @[Top.scala 432:12]
  assign n89_I1_2_2 = n88_O_2_2; // @[Top.scala 432:12]
  assign n89_I1_3_0 = n88_O_3_0; // @[Top.scala 432:12]
  assign n89_I1_3_1 = n88_O_3_1; // @[Top.scala 432:12]
  assign n89_I1_3_2 = n88_O_3_2; // @[Top.scala 432:12]
  assign n89_I1_4_0 = n88_O_4_0; // @[Top.scala 432:12]
  assign n89_I1_4_1 = n88_O_4_1; // @[Top.scala 432:12]
  assign n89_I1_4_2 = n88_O_4_2; // @[Top.scala 432:12]
  assign n89_I1_5_0 = n88_O_5_0; // @[Top.scala 432:12]
  assign n89_I1_5_1 = n88_O_5_1; // @[Top.scala 432:12]
  assign n89_I1_5_2 = n88_O_5_2; // @[Top.scala 432:12]
  assign n89_I1_6_0 = n88_O_6_0; // @[Top.scala 432:12]
  assign n89_I1_6_1 = n88_O_6_1; // @[Top.scala 432:12]
  assign n89_I1_6_2 = n88_O_6_2; // @[Top.scala 432:12]
  assign n89_I1_7_0 = n88_O_7_0; // @[Top.scala 432:12]
  assign n89_I1_7_1 = n88_O_7_1; // @[Top.scala 432:12]
  assign n89_I1_7_2 = n88_O_7_2; // @[Top.scala 432:12]
  assign n89_I1_8_0 = n88_O_8_0; // @[Top.scala 432:12]
  assign n89_I1_8_1 = n88_O_8_1; // @[Top.scala 432:12]
  assign n89_I1_8_2 = n88_O_8_2; // @[Top.scala 432:12]
  assign n89_I1_9_0 = n88_O_9_0; // @[Top.scala 432:12]
  assign n89_I1_9_1 = n88_O_9_1; // @[Top.scala 432:12]
  assign n89_I1_9_2 = n88_O_9_2; // @[Top.scala 432:12]
  assign n89_I1_10_0 = n88_O_10_0; // @[Top.scala 432:12]
  assign n89_I1_10_1 = n88_O_10_1; // @[Top.scala 432:12]
  assign n89_I1_10_2 = n88_O_10_2; // @[Top.scala 432:12]
  assign n89_I1_11_0 = n88_O_11_0; // @[Top.scala 432:12]
  assign n89_I1_11_1 = n88_O_11_1; // @[Top.scala 432:12]
  assign n89_I1_11_2 = n88_O_11_2; // @[Top.scala 432:12]
  assign n89_I1_12_0 = n88_O_12_0; // @[Top.scala 432:12]
  assign n89_I1_12_1 = n88_O_12_1; // @[Top.scala 432:12]
  assign n89_I1_12_2 = n88_O_12_2; // @[Top.scala 432:12]
  assign n89_I1_13_0 = n88_O_13_0; // @[Top.scala 432:12]
  assign n89_I1_13_1 = n88_O_13_1; // @[Top.scala 432:12]
  assign n89_I1_13_2 = n88_O_13_2; // @[Top.scala 432:12]
  assign n89_I1_14_0 = n88_O_14_0; // @[Top.scala 432:12]
  assign n89_I1_14_1 = n88_O_14_1; // @[Top.scala 432:12]
  assign n89_I1_14_2 = n88_O_14_2; // @[Top.scala 432:12]
  assign n89_I1_15_0 = n88_O_15_0; // @[Top.scala 432:12]
  assign n89_I1_15_1 = n88_O_15_1; // @[Top.scala 432:12]
  assign n89_I1_15_2 = n88_O_15_2; // @[Top.scala 432:12]
  assign n98_valid_up = n89_valid_down; // @[Top.scala 436:18]
  assign n98_I_0_0_0 = n89_O_0_0_0; // @[Top.scala 435:11]
  assign n98_I_0_0_1 = n89_O_0_0_1; // @[Top.scala 435:11]
  assign n98_I_0_0_2 = n89_O_0_0_2; // @[Top.scala 435:11]
  assign n98_I_0_1_0 = n89_O_0_1_0; // @[Top.scala 435:11]
  assign n98_I_0_1_1 = n89_O_0_1_1; // @[Top.scala 435:11]
  assign n98_I_0_1_2 = n89_O_0_1_2; // @[Top.scala 435:11]
  assign n98_I_0_2_0 = n89_O_0_2_0; // @[Top.scala 435:11]
  assign n98_I_0_2_1 = n89_O_0_2_1; // @[Top.scala 435:11]
  assign n98_I_0_2_2 = n89_O_0_2_2; // @[Top.scala 435:11]
  assign n98_I_1_0_0 = n89_O_1_0_0; // @[Top.scala 435:11]
  assign n98_I_1_0_1 = n89_O_1_0_1; // @[Top.scala 435:11]
  assign n98_I_1_0_2 = n89_O_1_0_2; // @[Top.scala 435:11]
  assign n98_I_1_1_0 = n89_O_1_1_0; // @[Top.scala 435:11]
  assign n98_I_1_1_1 = n89_O_1_1_1; // @[Top.scala 435:11]
  assign n98_I_1_1_2 = n89_O_1_1_2; // @[Top.scala 435:11]
  assign n98_I_1_2_0 = n89_O_1_2_0; // @[Top.scala 435:11]
  assign n98_I_1_2_1 = n89_O_1_2_1; // @[Top.scala 435:11]
  assign n98_I_1_2_2 = n89_O_1_2_2; // @[Top.scala 435:11]
  assign n98_I_2_0_0 = n89_O_2_0_0; // @[Top.scala 435:11]
  assign n98_I_2_0_1 = n89_O_2_0_1; // @[Top.scala 435:11]
  assign n98_I_2_0_2 = n89_O_2_0_2; // @[Top.scala 435:11]
  assign n98_I_2_1_0 = n89_O_2_1_0; // @[Top.scala 435:11]
  assign n98_I_2_1_1 = n89_O_2_1_1; // @[Top.scala 435:11]
  assign n98_I_2_1_2 = n89_O_2_1_2; // @[Top.scala 435:11]
  assign n98_I_2_2_0 = n89_O_2_2_0; // @[Top.scala 435:11]
  assign n98_I_2_2_1 = n89_O_2_2_1; // @[Top.scala 435:11]
  assign n98_I_2_2_2 = n89_O_2_2_2; // @[Top.scala 435:11]
  assign n98_I_3_0_0 = n89_O_3_0_0; // @[Top.scala 435:11]
  assign n98_I_3_0_1 = n89_O_3_0_1; // @[Top.scala 435:11]
  assign n98_I_3_0_2 = n89_O_3_0_2; // @[Top.scala 435:11]
  assign n98_I_3_1_0 = n89_O_3_1_0; // @[Top.scala 435:11]
  assign n98_I_3_1_1 = n89_O_3_1_1; // @[Top.scala 435:11]
  assign n98_I_3_1_2 = n89_O_3_1_2; // @[Top.scala 435:11]
  assign n98_I_3_2_0 = n89_O_3_2_0; // @[Top.scala 435:11]
  assign n98_I_3_2_1 = n89_O_3_2_1; // @[Top.scala 435:11]
  assign n98_I_3_2_2 = n89_O_3_2_2; // @[Top.scala 435:11]
  assign n98_I_4_0_0 = n89_O_4_0_0; // @[Top.scala 435:11]
  assign n98_I_4_0_1 = n89_O_4_0_1; // @[Top.scala 435:11]
  assign n98_I_4_0_2 = n89_O_4_0_2; // @[Top.scala 435:11]
  assign n98_I_4_1_0 = n89_O_4_1_0; // @[Top.scala 435:11]
  assign n98_I_4_1_1 = n89_O_4_1_1; // @[Top.scala 435:11]
  assign n98_I_4_1_2 = n89_O_4_1_2; // @[Top.scala 435:11]
  assign n98_I_4_2_0 = n89_O_4_2_0; // @[Top.scala 435:11]
  assign n98_I_4_2_1 = n89_O_4_2_1; // @[Top.scala 435:11]
  assign n98_I_4_2_2 = n89_O_4_2_2; // @[Top.scala 435:11]
  assign n98_I_5_0_0 = n89_O_5_0_0; // @[Top.scala 435:11]
  assign n98_I_5_0_1 = n89_O_5_0_1; // @[Top.scala 435:11]
  assign n98_I_5_0_2 = n89_O_5_0_2; // @[Top.scala 435:11]
  assign n98_I_5_1_0 = n89_O_5_1_0; // @[Top.scala 435:11]
  assign n98_I_5_1_1 = n89_O_5_1_1; // @[Top.scala 435:11]
  assign n98_I_5_1_2 = n89_O_5_1_2; // @[Top.scala 435:11]
  assign n98_I_5_2_0 = n89_O_5_2_0; // @[Top.scala 435:11]
  assign n98_I_5_2_1 = n89_O_5_2_1; // @[Top.scala 435:11]
  assign n98_I_5_2_2 = n89_O_5_2_2; // @[Top.scala 435:11]
  assign n98_I_6_0_0 = n89_O_6_0_0; // @[Top.scala 435:11]
  assign n98_I_6_0_1 = n89_O_6_0_1; // @[Top.scala 435:11]
  assign n98_I_6_0_2 = n89_O_6_0_2; // @[Top.scala 435:11]
  assign n98_I_6_1_0 = n89_O_6_1_0; // @[Top.scala 435:11]
  assign n98_I_6_1_1 = n89_O_6_1_1; // @[Top.scala 435:11]
  assign n98_I_6_1_2 = n89_O_6_1_2; // @[Top.scala 435:11]
  assign n98_I_6_2_0 = n89_O_6_2_0; // @[Top.scala 435:11]
  assign n98_I_6_2_1 = n89_O_6_2_1; // @[Top.scala 435:11]
  assign n98_I_6_2_2 = n89_O_6_2_2; // @[Top.scala 435:11]
  assign n98_I_7_0_0 = n89_O_7_0_0; // @[Top.scala 435:11]
  assign n98_I_7_0_1 = n89_O_7_0_1; // @[Top.scala 435:11]
  assign n98_I_7_0_2 = n89_O_7_0_2; // @[Top.scala 435:11]
  assign n98_I_7_1_0 = n89_O_7_1_0; // @[Top.scala 435:11]
  assign n98_I_7_1_1 = n89_O_7_1_1; // @[Top.scala 435:11]
  assign n98_I_7_1_2 = n89_O_7_1_2; // @[Top.scala 435:11]
  assign n98_I_7_2_0 = n89_O_7_2_0; // @[Top.scala 435:11]
  assign n98_I_7_2_1 = n89_O_7_2_1; // @[Top.scala 435:11]
  assign n98_I_7_2_2 = n89_O_7_2_2; // @[Top.scala 435:11]
  assign n98_I_8_0_0 = n89_O_8_0_0; // @[Top.scala 435:11]
  assign n98_I_8_0_1 = n89_O_8_0_1; // @[Top.scala 435:11]
  assign n98_I_8_0_2 = n89_O_8_0_2; // @[Top.scala 435:11]
  assign n98_I_8_1_0 = n89_O_8_1_0; // @[Top.scala 435:11]
  assign n98_I_8_1_1 = n89_O_8_1_1; // @[Top.scala 435:11]
  assign n98_I_8_1_2 = n89_O_8_1_2; // @[Top.scala 435:11]
  assign n98_I_8_2_0 = n89_O_8_2_0; // @[Top.scala 435:11]
  assign n98_I_8_2_1 = n89_O_8_2_1; // @[Top.scala 435:11]
  assign n98_I_8_2_2 = n89_O_8_2_2; // @[Top.scala 435:11]
  assign n98_I_9_0_0 = n89_O_9_0_0; // @[Top.scala 435:11]
  assign n98_I_9_0_1 = n89_O_9_0_1; // @[Top.scala 435:11]
  assign n98_I_9_0_2 = n89_O_9_0_2; // @[Top.scala 435:11]
  assign n98_I_9_1_0 = n89_O_9_1_0; // @[Top.scala 435:11]
  assign n98_I_9_1_1 = n89_O_9_1_1; // @[Top.scala 435:11]
  assign n98_I_9_1_2 = n89_O_9_1_2; // @[Top.scala 435:11]
  assign n98_I_9_2_0 = n89_O_9_2_0; // @[Top.scala 435:11]
  assign n98_I_9_2_1 = n89_O_9_2_1; // @[Top.scala 435:11]
  assign n98_I_9_2_2 = n89_O_9_2_2; // @[Top.scala 435:11]
  assign n98_I_10_0_0 = n89_O_10_0_0; // @[Top.scala 435:11]
  assign n98_I_10_0_1 = n89_O_10_0_1; // @[Top.scala 435:11]
  assign n98_I_10_0_2 = n89_O_10_0_2; // @[Top.scala 435:11]
  assign n98_I_10_1_0 = n89_O_10_1_0; // @[Top.scala 435:11]
  assign n98_I_10_1_1 = n89_O_10_1_1; // @[Top.scala 435:11]
  assign n98_I_10_1_2 = n89_O_10_1_2; // @[Top.scala 435:11]
  assign n98_I_10_2_0 = n89_O_10_2_0; // @[Top.scala 435:11]
  assign n98_I_10_2_1 = n89_O_10_2_1; // @[Top.scala 435:11]
  assign n98_I_10_2_2 = n89_O_10_2_2; // @[Top.scala 435:11]
  assign n98_I_11_0_0 = n89_O_11_0_0; // @[Top.scala 435:11]
  assign n98_I_11_0_1 = n89_O_11_0_1; // @[Top.scala 435:11]
  assign n98_I_11_0_2 = n89_O_11_0_2; // @[Top.scala 435:11]
  assign n98_I_11_1_0 = n89_O_11_1_0; // @[Top.scala 435:11]
  assign n98_I_11_1_1 = n89_O_11_1_1; // @[Top.scala 435:11]
  assign n98_I_11_1_2 = n89_O_11_1_2; // @[Top.scala 435:11]
  assign n98_I_11_2_0 = n89_O_11_2_0; // @[Top.scala 435:11]
  assign n98_I_11_2_1 = n89_O_11_2_1; // @[Top.scala 435:11]
  assign n98_I_11_2_2 = n89_O_11_2_2; // @[Top.scala 435:11]
  assign n98_I_12_0_0 = n89_O_12_0_0; // @[Top.scala 435:11]
  assign n98_I_12_0_1 = n89_O_12_0_1; // @[Top.scala 435:11]
  assign n98_I_12_0_2 = n89_O_12_0_2; // @[Top.scala 435:11]
  assign n98_I_12_1_0 = n89_O_12_1_0; // @[Top.scala 435:11]
  assign n98_I_12_1_1 = n89_O_12_1_1; // @[Top.scala 435:11]
  assign n98_I_12_1_2 = n89_O_12_1_2; // @[Top.scala 435:11]
  assign n98_I_12_2_0 = n89_O_12_2_0; // @[Top.scala 435:11]
  assign n98_I_12_2_1 = n89_O_12_2_1; // @[Top.scala 435:11]
  assign n98_I_12_2_2 = n89_O_12_2_2; // @[Top.scala 435:11]
  assign n98_I_13_0_0 = n89_O_13_0_0; // @[Top.scala 435:11]
  assign n98_I_13_0_1 = n89_O_13_0_1; // @[Top.scala 435:11]
  assign n98_I_13_0_2 = n89_O_13_0_2; // @[Top.scala 435:11]
  assign n98_I_13_1_0 = n89_O_13_1_0; // @[Top.scala 435:11]
  assign n98_I_13_1_1 = n89_O_13_1_1; // @[Top.scala 435:11]
  assign n98_I_13_1_2 = n89_O_13_1_2; // @[Top.scala 435:11]
  assign n98_I_13_2_0 = n89_O_13_2_0; // @[Top.scala 435:11]
  assign n98_I_13_2_1 = n89_O_13_2_1; // @[Top.scala 435:11]
  assign n98_I_13_2_2 = n89_O_13_2_2; // @[Top.scala 435:11]
  assign n98_I_14_0_0 = n89_O_14_0_0; // @[Top.scala 435:11]
  assign n98_I_14_0_1 = n89_O_14_0_1; // @[Top.scala 435:11]
  assign n98_I_14_0_2 = n89_O_14_0_2; // @[Top.scala 435:11]
  assign n98_I_14_1_0 = n89_O_14_1_0; // @[Top.scala 435:11]
  assign n98_I_14_1_1 = n89_O_14_1_1; // @[Top.scala 435:11]
  assign n98_I_14_1_2 = n89_O_14_1_2; // @[Top.scala 435:11]
  assign n98_I_14_2_0 = n89_O_14_2_0; // @[Top.scala 435:11]
  assign n98_I_14_2_1 = n89_O_14_2_1; // @[Top.scala 435:11]
  assign n98_I_14_2_2 = n89_O_14_2_2; // @[Top.scala 435:11]
  assign n98_I_15_0_0 = n89_O_15_0_0; // @[Top.scala 435:11]
  assign n98_I_15_0_1 = n89_O_15_0_1; // @[Top.scala 435:11]
  assign n98_I_15_0_2 = n89_O_15_0_2; // @[Top.scala 435:11]
  assign n98_I_15_1_0 = n89_O_15_1_0; // @[Top.scala 435:11]
  assign n98_I_15_1_1 = n89_O_15_1_1; // @[Top.scala 435:11]
  assign n98_I_15_1_2 = n89_O_15_1_2; // @[Top.scala 435:11]
  assign n98_I_15_2_0 = n89_O_15_2_0; // @[Top.scala 435:11]
  assign n98_I_15_2_1 = n89_O_15_2_1; // @[Top.scala 435:11]
  assign n98_I_15_2_2 = n89_O_15_2_2; // @[Top.scala 435:11]
  assign n105_valid_up = n98_valid_down; // @[Top.scala 439:19]
  assign n105_I_0_0_0_0 = n98_O_0_0_0_0; // @[Top.scala 438:12]
  assign n105_I_0_0_0_1 = n98_O_0_0_0_1; // @[Top.scala 438:12]
  assign n105_I_0_0_0_2 = n98_O_0_0_0_2; // @[Top.scala 438:12]
  assign n105_I_0_0_1_0 = n98_O_0_0_1_0; // @[Top.scala 438:12]
  assign n105_I_0_0_1_1 = n98_O_0_0_1_1; // @[Top.scala 438:12]
  assign n105_I_0_0_1_2 = n98_O_0_0_1_2; // @[Top.scala 438:12]
  assign n105_I_0_0_2_0 = n98_O_0_0_2_0; // @[Top.scala 438:12]
  assign n105_I_0_0_2_1 = n98_O_0_0_2_1; // @[Top.scala 438:12]
  assign n105_I_0_0_2_2 = n98_O_0_0_2_2; // @[Top.scala 438:12]
  assign n105_I_1_0_0_0 = n98_O_1_0_0_0; // @[Top.scala 438:12]
  assign n105_I_1_0_0_1 = n98_O_1_0_0_1; // @[Top.scala 438:12]
  assign n105_I_1_0_0_2 = n98_O_1_0_0_2; // @[Top.scala 438:12]
  assign n105_I_1_0_1_0 = n98_O_1_0_1_0; // @[Top.scala 438:12]
  assign n105_I_1_0_1_1 = n98_O_1_0_1_1; // @[Top.scala 438:12]
  assign n105_I_1_0_1_2 = n98_O_1_0_1_2; // @[Top.scala 438:12]
  assign n105_I_1_0_2_0 = n98_O_1_0_2_0; // @[Top.scala 438:12]
  assign n105_I_1_0_2_1 = n98_O_1_0_2_1; // @[Top.scala 438:12]
  assign n105_I_1_0_2_2 = n98_O_1_0_2_2; // @[Top.scala 438:12]
  assign n105_I_2_0_0_0 = n98_O_2_0_0_0; // @[Top.scala 438:12]
  assign n105_I_2_0_0_1 = n98_O_2_0_0_1; // @[Top.scala 438:12]
  assign n105_I_2_0_0_2 = n98_O_2_0_0_2; // @[Top.scala 438:12]
  assign n105_I_2_0_1_0 = n98_O_2_0_1_0; // @[Top.scala 438:12]
  assign n105_I_2_0_1_1 = n98_O_2_0_1_1; // @[Top.scala 438:12]
  assign n105_I_2_0_1_2 = n98_O_2_0_1_2; // @[Top.scala 438:12]
  assign n105_I_2_0_2_0 = n98_O_2_0_2_0; // @[Top.scala 438:12]
  assign n105_I_2_0_2_1 = n98_O_2_0_2_1; // @[Top.scala 438:12]
  assign n105_I_2_0_2_2 = n98_O_2_0_2_2; // @[Top.scala 438:12]
  assign n105_I_3_0_0_0 = n98_O_3_0_0_0; // @[Top.scala 438:12]
  assign n105_I_3_0_0_1 = n98_O_3_0_0_1; // @[Top.scala 438:12]
  assign n105_I_3_0_0_2 = n98_O_3_0_0_2; // @[Top.scala 438:12]
  assign n105_I_3_0_1_0 = n98_O_3_0_1_0; // @[Top.scala 438:12]
  assign n105_I_3_0_1_1 = n98_O_3_0_1_1; // @[Top.scala 438:12]
  assign n105_I_3_0_1_2 = n98_O_3_0_1_2; // @[Top.scala 438:12]
  assign n105_I_3_0_2_0 = n98_O_3_0_2_0; // @[Top.scala 438:12]
  assign n105_I_3_0_2_1 = n98_O_3_0_2_1; // @[Top.scala 438:12]
  assign n105_I_3_0_2_2 = n98_O_3_0_2_2; // @[Top.scala 438:12]
  assign n105_I_4_0_0_0 = n98_O_4_0_0_0; // @[Top.scala 438:12]
  assign n105_I_4_0_0_1 = n98_O_4_0_0_1; // @[Top.scala 438:12]
  assign n105_I_4_0_0_2 = n98_O_4_0_0_2; // @[Top.scala 438:12]
  assign n105_I_4_0_1_0 = n98_O_4_0_1_0; // @[Top.scala 438:12]
  assign n105_I_4_0_1_1 = n98_O_4_0_1_1; // @[Top.scala 438:12]
  assign n105_I_4_0_1_2 = n98_O_4_0_1_2; // @[Top.scala 438:12]
  assign n105_I_4_0_2_0 = n98_O_4_0_2_0; // @[Top.scala 438:12]
  assign n105_I_4_0_2_1 = n98_O_4_0_2_1; // @[Top.scala 438:12]
  assign n105_I_4_0_2_2 = n98_O_4_0_2_2; // @[Top.scala 438:12]
  assign n105_I_5_0_0_0 = n98_O_5_0_0_0; // @[Top.scala 438:12]
  assign n105_I_5_0_0_1 = n98_O_5_0_0_1; // @[Top.scala 438:12]
  assign n105_I_5_0_0_2 = n98_O_5_0_0_2; // @[Top.scala 438:12]
  assign n105_I_5_0_1_0 = n98_O_5_0_1_0; // @[Top.scala 438:12]
  assign n105_I_5_0_1_1 = n98_O_5_0_1_1; // @[Top.scala 438:12]
  assign n105_I_5_0_1_2 = n98_O_5_0_1_2; // @[Top.scala 438:12]
  assign n105_I_5_0_2_0 = n98_O_5_0_2_0; // @[Top.scala 438:12]
  assign n105_I_5_0_2_1 = n98_O_5_0_2_1; // @[Top.scala 438:12]
  assign n105_I_5_0_2_2 = n98_O_5_0_2_2; // @[Top.scala 438:12]
  assign n105_I_6_0_0_0 = n98_O_6_0_0_0; // @[Top.scala 438:12]
  assign n105_I_6_0_0_1 = n98_O_6_0_0_1; // @[Top.scala 438:12]
  assign n105_I_6_0_0_2 = n98_O_6_0_0_2; // @[Top.scala 438:12]
  assign n105_I_6_0_1_0 = n98_O_6_0_1_0; // @[Top.scala 438:12]
  assign n105_I_6_0_1_1 = n98_O_6_0_1_1; // @[Top.scala 438:12]
  assign n105_I_6_0_1_2 = n98_O_6_0_1_2; // @[Top.scala 438:12]
  assign n105_I_6_0_2_0 = n98_O_6_0_2_0; // @[Top.scala 438:12]
  assign n105_I_6_0_2_1 = n98_O_6_0_2_1; // @[Top.scala 438:12]
  assign n105_I_6_0_2_2 = n98_O_6_0_2_2; // @[Top.scala 438:12]
  assign n105_I_7_0_0_0 = n98_O_7_0_0_0; // @[Top.scala 438:12]
  assign n105_I_7_0_0_1 = n98_O_7_0_0_1; // @[Top.scala 438:12]
  assign n105_I_7_0_0_2 = n98_O_7_0_0_2; // @[Top.scala 438:12]
  assign n105_I_7_0_1_0 = n98_O_7_0_1_0; // @[Top.scala 438:12]
  assign n105_I_7_0_1_1 = n98_O_7_0_1_1; // @[Top.scala 438:12]
  assign n105_I_7_0_1_2 = n98_O_7_0_1_2; // @[Top.scala 438:12]
  assign n105_I_7_0_2_0 = n98_O_7_0_2_0; // @[Top.scala 438:12]
  assign n105_I_7_0_2_1 = n98_O_7_0_2_1; // @[Top.scala 438:12]
  assign n105_I_7_0_2_2 = n98_O_7_0_2_2; // @[Top.scala 438:12]
  assign n105_I_8_0_0_0 = n98_O_8_0_0_0; // @[Top.scala 438:12]
  assign n105_I_8_0_0_1 = n98_O_8_0_0_1; // @[Top.scala 438:12]
  assign n105_I_8_0_0_2 = n98_O_8_0_0_2; // @[Top.scala 438:12]
  assign n105_I_8_0_1_0 = n98_O_8_0_1_0; // @[Top.scala 438:12]
  assign n105_I_8_0_1_1 = n98_O_8_0_1_1; // @[Top.scala 438:12]
  assign n105_I_8_0_1_2 = n98_O_8_0_1_2; // @[Top.scala 438:12]
  assign n105_I_8_0_2_0 = n98_O_8_0_2_0; // @[Top.scala 438:12]
  assign n105_I_8_0_2_1 = n98_O_8_0_2_1; // @[Top.scala 438:12]
  assign n105_I_8_0_2_2 = n98_O_8_0_2_2; // @[Top.scala 438:12]
  assign n105_I_9_0_0_0 = n98_O_9_0_0_0; // @[Top.scala 438:12]
  assign n105_I_9_0_0_1 = n98_O_9_0_0_1; // @[Top.scala 438:12]
  assign n105_I_9_0_0_2 = n98_O_9_0_0_2; // @[Top.scala 438:12]
  assign n105_I_9_0_1_0 = n98_O_9_0_1_0; // @[Top.scala 438:12]
  assign n105_I_9_0_1_1 = n98_O_9_0_1_1; // @[Top.scala 438:12]
  assign n105_I_9_0_1_2 = n98_O_9_0_1_2; // @[Top.scala 438:12]
  assign n105_I_9_0_2_0 = n98_O_9_0_2_0; // @[Top.scala 438:12]
  assign n105_I_9_0_2_1 = n98_O_9_0_2_1; // @[Top.scala 438:12]
  assign n105_I_9_0_2_2 = n98_O_9_0_2_2; // @[Top.scala 438:12]
  assign n105_I_10_0_0_0 = n98_O_10_0_0_0; // @[Top.scala 438:12]
  assign n105_I_10_0_0_1 = n98_O_10_0_0_1; // @[Top.scala 438:12]
  assign n105_I_10_0_0_2 = n98_O_10_0_0_2; // @[Top.scala 438:12]
  assign n105_I_10_0_1_0 = n98_O_10_0_1_0; // @[Top.scala 438:12]
  assign n105_I_10_0_1_1 = n98_O_10_0_1_1; // @[Top.scala 438:12]
  assign n105_I_10_0_1_2 = n98_O_10_0_1_2; // @[Top.scala 438:12]
  assign n105_I_10_0_2_0 = n98_O_10_0_2_0; // @[Top.scala 438:12]
  assign n105_I_10_0_2_1 = n98_O_10_0_2_1; // @[Top.scala 438:12]
  assign n105_I_10_0_2_2 = n98_O_10_0_2_2; // @[Top.scala 438:12]
  assign n105_I_11_0_0_0 = n98_O_11_0_0_0; // @[Top.scala 438:12]
  assign n105_I_11_0_0_1 = n98_O_11_0_0_1; // @[Top.scala 438:12]
  assign n105_I_11_0_0_2 = n98_O_11_0_0_2; // @[Top.scala 438:12]
  assign n105_I_11_0_1_0 = n98_O_11_0_1_0; // @[Top.scala 438:12]
  assign n105_I_11_0_1_1 = n98_O_11_0_1_1; // @[Top.scala 438:12]
  assign n105_I_11_0_1_2 = n98_O_11_0_1_2; // @[Top.scala 438:12]
  assign n105_I_11_0_2_0 = n98_O_11_0_2_0; // @[Top.scala 438:12]
  assign n105_I_11_0_2_1 = n98_O_11_0_2_1; // @[Top.scala 438:12]
  assign n105_I_11_0_2_2 = n98_O_11_0_2_2; // @[Top.scala 438:12]
  assign n105_I_12_0_0_0 = n98_O_12_0_0_0; // @[Top.scala 438:12]
  assign n105_I_12_0_0_1 = n98_O_12_0_0_1; // @[Top.scala 438:12]
  assign n105_I_12_0_0_2 = n98_O_12_0_0_2; // @[Top.scala 438:12]
  assign n105_I_12_0_1_0 = n98_O_12_0_1_0; // @[Top.scala 438:12]
  assign n105_I_12_0_1_1 = n98_O_12_0_1_1; // @[Top.scala 438:12]
  assign n105_I_12_0_1_2 = n98_O_12_0_1_2; // @[Top.scala 438:12]
  assign n105_I_12_0_2_0 = n98_O_12_0_2_0; // @[Top.scala 438:12]
  assign n105_I_12_0_2_1 = n98_O_12_0_2_1; // @[Top.scala 438:12]
  assign n105_I_12_0_2_2 = n98_O_12_0_2_2; // @[Top.scala 438:12]
  assign n105_I_13_0_0_0 = n98_O_13_0_0_0; // @[Top.scala 438:12]
  assign n105_I_13_0_0_1 = n98_O_13_0_0_1; // @[Top.scala 438:12]
  assign n105_I_13_0_0_2 = n98_O_13_0_0_2; // @[Top.scala 438:12]
  assign n105_I_13_0_1_0 = n98_O_13_0_1_0; // @[Top.scala 438:12]
  assign n105_I_13_0_1_1 = n98_O_13_0_1_1; // @[Top.scala 438:12]
  assign n105_I_13_0_1_2 = n98_O_13_0_1_2; // @[Top.scala 438:12]
  assign n105_I_13_0_2_0 = n98_O_13_0_2_0; // @[Top.scala 438:12]
  assign n105_I_13_0_2_1 = n98_O_13_0_2_1; // @[Top.scala 438:12]
  assign n105_I_13_0_2_2 = n98_O_13_0_2_2; // @[Top.scala 438:12]
  assign n105_I_14_0_0_0 = n98_O_14_0_0_0; // @[Top.scala 438:12]
  assign n105_I_14_0_0_1 = n98_O_14_0_0_1; // @[Top.scala 438:12]
  assign n105_I_14_0_0_2 = n98_O_14_0_0_2; // @[Top.scala 438:12]
  assign n105_I_14_0_1_0 = n98_O_14_0_1_0; // @[Top.scala 438:12]
  assign n105_I_14_0_1_1 = n98_O_14_0_1_1; // @[Top.scala 438:12]
  assign n105_I_14_0_1_2 = n98_O_14_0_1_2; // @[Top.scala 438:12]
  assign n105_I_14_0_2_0 = n98_O_14_0_2_0; // @[Top.scala 438:12]
  assign n105_I_14_0_2_1 = n98_O_14_0_2_1; // @[Top.scala 438:12]
  assign n105_I_14_0_2_2 = n98_O_14_0_2_2; // @[Top.scala 438:12]
  assign n105_I_15_0_0_0 = n98_O_15_0_0_0; // @[Top.scala 438:12]
  assign n105_I_15_0_0_1 = n98_O_15_0_0_1; // @[Top.scala 438:12]
  assign n105_I_15_0_0_2 = n98_O_15_0_0_2; // @[Top.scala 438:12]
  assign n105_I_15_0_1_0 = n98_O_15_0_1_0; // @[Top.scala 438:12]
  assign n105_I_15_0_1_1 = n98_O_15_0_1_1; // @[Top.scala 438:12]
  assign n105_I_15_0_1_2 = n98_O_15_0_1_2; // @[Top.scala 438:12]
  assign n105_I_15_0_2_0 = n98_O_15_0_2_0; // @[Top.scala 438:12]
  assign n105_I_15_0_2_1 = n98_O_15_0_2_1; // @[Top.scala 438:12]
  assign n105_I_15_0_2_2 = n98_O_15_0_2_2; // @[Top.scala 438:12]
  assign n106_valid_up = n105_valid_down; // @[Top.scala 442:19]
  assign n106_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 441:12]
  assign n106_I_0_0_1 = n105_O_0_0_1; // @[Top.scala 441:12]
  assign n106_I_0_0_2 = n105_O_0_0_2; // @[Top.scala 441:12]
  assign n106_I_0_1_0 = n105_O_0_1_0; // @[Top.scala 441:12]
  assign n106_I_0_1_1 = n105_O_0_1_1; // @[Top.scala 441:12]
  assign n106_I_0_1_2 = n105_O_0_1_2; // @[Top.scala 441:12]
  assign n106_I_0_2_0 = n105_O_0_2_0; // @[Top.scala 441:12]
  assign n106_I_0_2_1 = n105_O_0_2_1; // @[Top.scala 441:12]
  assign n106_I_0_2_2 = n105_O_0_2_2; // @[Top.scala 441:12]
  assign n106_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 441:12]
  assign n106_I_1_0_1 = n105_O_1_0_1; // @[Top.scala 441:12]
  assign n106_I_1_0_2 = n105_O_1_0_2; // @[Top.scala 441:12]
  assign n106_I_1_1_0 = n105_O_1_1_0; // @[Top.scala 441:12]
  assign n106_I_1_1_1 = n105_O_1_1_1; // @[Top.scala 441:12]
  assign n106_I_1_1_2 = n105_O_1_1_2; // @[Top.scala 441:12]
  assign n106_I_1_2_0 = n105_O_1_2_0; // @[Top.scala 441:12]
  assign n106_I_1_2_1 = n105_O_1_2_1; // @[Top.scala 441:12]
  assign n106_I_1_2_2 = n105_O_1_2_2; // @[Top.scala 441:12]
  assign n106_I_2_0_0 = n105_O_2_0_0; // @[Top.scala 441:12]
  assign n106_I_2_0_1 = n105_O_2_0_1; // @[Top.scala 441:12]
  assign n106_I_2_0_2 = n105_O_2_0_2; // @[Top.scala 441:12]
  assign n106_I_2_1_0 = n105_O_2_1_0; // @[Top.scala 441:12]
  assign n106_I_2_1_1 = n105_O_2_1_1; // @[Top.scala 441:12]
  assign n106_I_2_1_2 = n105_O_2_1_2; // @[Top.scala 441:12]
  assign n106_I_2_2_0 = n105_O_2_2_0; // @[Top.scala 441:12]
  assign n106_I_2_2_1 = n105_O_2_2_1; // @[Top.scala 441:12]
  assign n106_I_2_2_2 = n105_O_2_2_2; // @[Top.scala 441:12]
  assign n106_I_3_0_0 = n105_O_3_0_0; // @[Top.scala 441:12]
  assign n106_I_3_0_1 = n105_O_3_0_1; // @[Top.scala 441:12]
  assign n106_I_3_0_2 = n105_O_3_0_2; // @[Top.scala 441:12]
  assign n106_I_3_1_0 = n105_O_3_1_0; // @[Top.scala 441:12]
  assign n106_I_3_1_1 = n105_O_3_1_1; // @[Top.scala 441:12]
  assign n106_I_3_1_2 = n105_O_3_1_2; // @[Top.scala 441:12]
  assign n106_I_3_2_0 = n105_O_3_2_0; // @[Top.scala 441:12]
  assign n106_I_3_2_1 = n105_O_3_2_1; // @[Top.scala 441:12]
  assign n106_I_3_2_2 = n105_O_3_2_2; // @[Top.scala 441:12]
  assign n106_I_4_0_0 = n105_O_4_0_0; // @[Top.scala 441:12]
  assign n106_I_4_0_1 = n105_O_4_0_1; // @[Top.scala 441:12]
  assign n106_I_4_0_2 = n105_O_4_0_2; // @[Top.scala 441:12]
  assign n106_I_4_1_0 = n105_O_4_1_0; // @[Top.scala 441:12]
  assign n106_I_4_1_1 = n105_O_4_1_1; // @[Top.scala 441:12]
  assign n106_I_4_1_2 = n105_O_4_1_2; // @[Top.scala 441:12]
  assign n106_I_4_2_0 = n105_O_4_2_0; // @[Top.scala 441:12]
  assign n106_I_4_2_1 = n105_O_4_2_1; // @[Top.scala 441:12]
  assign n106_I_4_2_2 = n105_O_4_2_2; // @[Top.scala 441:12]
  assign n106_I_5_0_0 = n105_O_5_0_0; // @[Top.scala 441:12]
  assign n106_I_5_0_1 = n105_O_5_0_1; // @[Top.scala 441:12]
  assign n106_I_5_0_2 = n105_O_5_0_2; // @[Top.scala 441:12]
  assign n106_I_5_1_0 = n105_O_5_1_0; // @[Top.scala 441:12]
  assign n106_I_5_1_1 = n105_O_5_1_1; // @[Top.scala 441:12]
  assign n106_I_5_1_2 = n105_O_5_1_2; // @[Top.scala 441:12]
  assign n106_I_5_2_0 = n105_O_5_2_0; // @[Top.scala 441:12]
  assign n106_I_5_2_1 = n105_O_5_2_1; // @[Top.scala 441:12]
  assign n106_I_5_2_2 = n105_O_5_2_2; // @[Top.scala 441:12]
  assign n106_I_6_0_0 = n105_O_6_0_0; // @[Top.scala 441:12]
  assign n106_I_6_0_1 = n105_O_6_0_1; // @[Top.scala 441:12]
  assign n106_I_6_0_2 = n105_O_6_0_2; // @[Top.scala 441:12]
  assign n106_I_6_1_0 = n105_O_6_1_0; // @[Top.scala 441:12]
  assign n106_I_6_1_1 = n105_O_6_1_1; // @[Top.scala 441:12]
  assign n106_I_6_1_2 = n105_O_6_1_2; // @[Top.scala 441:12]
  assign n106_I_6_2_0 = n105_O_6_2_0; // @[Top.scala 441:12]
  assign n106_I_6_2_1 = n105_O_6_2_1; // @[Top.scala 441:12]
  assign n106_I_6_2_2 = n105_O_6_2_2; // @[Top.scala 441:12]
  assign n106_I_7_0_0 = n105_O_7_0_0; // @[Top.scala 441:12]
  assign n106_I_7_0_1 = n105_O_7_0_1; // @[Top.scala 441:12]
  assign n106_I_7_0_2 = n105_O_7_0_2; // @[Top.scala 441:12]
  assign n106_I_7_1_0 = n105_O_7_1_0; // @[Top.scala 441:12]
  assign n106_I_7_1_1 = n105_O_7_1_1; // @[Top.scala 441:12]
  assign n106_I_7_1_2 = n105_O_7_1_2; // @[Top.scala 441:12]
  assign n106_I_7_2_0 = n105_O_7_2_0; // @[Top.scala 441:12]
  assign n106_I_7_2_1 = n105_O_7_2_1; // @[Top.scala 441:12]
  assign n106_I_7_2_2 = n105_O_7_2_2; // @[Top.scala 441:12]
  assign n106_I_8_0_0 = n105_O_8_0_0; // @[Top.scala 441:12]
  assign n106_I_8_0_1 = n105_O_8_0_1; // @[Top.scala 441:12]
  assign n106_I_8_0_2 = n105_O_8_0_2; // @[Top.scala 441:12]
  assign n106_I_8_1_0 = n105_O_8_1_0; // @[Top.scala 441:12]
  assign n106_I_8_1_1 = n105_O_8_1_1; // @[Top.scala 441:12]
  assign n106_I_8_1_2 = n105_O_8_1_2; // @[Top.scala 441:12]
  assign n106_I_8_2_0 = n105_O_8_2_0; // @[Top.scala 441:12]
  assign n106_I_8_2_1 = n105_O_8_2_1; // @[Top.scala 441:12]
  assign n106_I_8_2_2 = n105_O_8_2_2; // @[Top.scala 441:12]
  assign n106_I_9_0_0 = n105_O_9_0_0; // @[Top.scala 441:12]
  assign n106_I_9_0_1 = n105_O_9_0_1; // @[Top.scala 441:12]
  assign n106_I_9_0_2 = n105_O_9_0_2; // @[Top.scala 441:12]
  assign n106_I_9_1_0 = n105_O_9_1_0; // @[Top.scala 441:12]
  assign n106_I_9_1_1 = n105_O_9_1_1; // @[Top.scala 441:12]
  assign n106_I_9_1_2 = n105_O_9_1_2; // @[Top.scala 441:12]
  assign n106_I_9_2_0 = n105_O_9_2_0; // @[Top.scala 441:12]
  assign n106_I_9_2_1 = n105_O_9_2_1; // @[Top.scala 441:12]
  assign n106_I_9_2_2 = n105_O_9_2_2; // @[Top.scala 441:12]
  assign n106_I_10_0_0 = n105_O_10_0_0; // @[Top.scala 441:12]
  assign n106_I_10_0_1 = n105_O_10_0_1; // @[Top.scala 441:12]
  assign n106_I_10_0_2 = n105_O_10_0_2; // @[Top.scala 441:12]
  assign n106_I_10_1_0 = n105_O_10_1_0; // @[Top.scala 441:12]
  assign n106_I_10_1_1 = n105_O_10_1_1; // @[Top.scala 441:12]
  assign n106_I_10_1_2 = n105_O_10_1_2; // @[Top.scala 441:12]
  assign n106_I_10_2_0 = n105_O_10_2_0; // @[Top.scala 441:12]
  assign n106_I_10_2_1 = n105_O_10_2_1; // @[Top.scala 441:12]
  assign n106_I_10_2_2 = n105_O_10_2_2; // @[Top.scala 441:12]
  assign n106_I_11_0_0 = n105_O_11_0_0; // @[Top.scala 441:12]
  assign n106_I_11_0_1 = n105_O_11_0_1; // @[Top.scala 441:12]
  assign n106_I_11_0_2 = n105_O_11_0_2; // @[Top.scala 441:12]
  assign n106_I_11_1_0 = n105_O_11_1_0; // @[Top.scala 441:12]
  assign n106_I_11_1_1 = n105_O_11_1_1; // @[Top.scala 441:12]
  assign n106_I_11_1_2 = n105_O_11_1_2; // @[Top.scala 441:12]
  assign n106_I_11_2_0 = n105_O_11_2_0; // @[Top.scala 441:12]
  assign n106_I_11_2_1 = n105_O_11_2_1; // @[Top.scala 441:12]
  assign n106_I_11_2_2 = n105_O_11_2_2; // @[Top.scala 441:12]
  assign n106_I_12_0_0 = n105_O_12_0_0; // @[Top.scala 441:12]
  assign n106_I_12_0_1 = n105_O_12_0_1; // @[Top.scala 441:12]
  assign n106_I_12_0_2 = n105_O_12_0_2; // @[Top.scala 441:12]
  assign n106_I_12_1_0 = n105_O_12_1_0; // @[Top.scala 441:12]
  assign n106_I_12_1_1 = n105_O_12_1_1; // @[Top.scala 441:12]
  assign n106_I_12_1_2 = n105_O_12_1_2; // @[Top.scala 441:12]
  assign n106_I_12_2_0 = n105_O_12_2_0; // @[Top.scala 441:12]
  assign n106_I_12_2_1 = n105_O_12_2_1; // @[Top.scala 441:12]
  assign n106_I_12_2_2 = n105_O_12_2_2; // @[Top.scala 441:12]
  assign n106_I_13_0_0 = n105_O_13_0_0; // @[Top.scala 441:12]
  assign n106_I_13_0_1 = n105_O_13_0_1; // @[Top.scala 441:12]
  assign n106_I_13_0_2 = n105_O_13_0_2; // @[Top.scala 441:12]
  assign n106_I_13_1_0 = n105_O_13_1_0; // @[Top.scala 441:12]
  assign n106_I_13_1_1 = n105_O_13_1_1; // @[Top.scala 441:12]
  assign n106_I_13_1_2 = n105_O_13_1_2; // @[Top.scala 441:12]
  assign n106_I_13_2_0 = n105_O_13_2_0; // @[Top.scala 441:12]
  assign n106_I_13_2_1 = n105_O_13_2_1; // @[Top.scala 441:12]
  assign n106_I_13_2_2 = n105_O_13_2_2; // @[Top.scala 441:12]
  assign n106_I_14_0_0 = n105_O_14_0_0; // @[Top.scala 441:12]
  assign n106_I_14_0_1 = n105_O_14_0_1; // @[Top.scala 441:12]
  assign n106_I_14_0_2 = n105_O_14_0_2; // @[Top.scala 441:12]
  assign n106_I_14_1_0 = n105_O_14_1_0; // @[Top.scala 441:12]
  assign n106_I_14_1_1 = n105_O_14_1_1; // @[Top.scala 441:12]
  assign n106_I_14_1_2 = n105_O_14_1_2; // @[Top.scala 441:12]
  assign n106_I_14_2_0 = n105_O_14_2_0; // @[Top.scala 441:12]
  assign n106_I_14_2_1 = n105_O_14_2_1; // @[Top.scala 441:12]
  assign n106_I_14_2_2 = n105_O_14_2_2; // @[Top.scala 441:12]
  assign n106_I_15_0_0 = n105_O_15_0_0; // @[Top.scala 441:12]
  assign n106_I_15_0_1 = n105_O_15_0_1; // @[Top.scala 441:12]
  assign n106_I_15_0_2 = n105_O_15_0_2; // @[Top.scala 441:12]
  assign n106_I_15_1_0 = n105_O_15_1_0; // @[Top.scala 441:12]
  assign n106_I_15_1_1 = n105_O_15_1_1; // @[Top.scala 441:12]
  assign n106_I_15_1_2 = n105_O_15_1_2; // @[Top.scala 441:12]
  assign n106_I_15_2_0 = n105_O_15_2_0; // @[Top.scala 441:12]
  assign n106_I_15_2_1 = n105_O_15_2_1; // @[Top.scala 441:12]
  assign n106_I_15_2_2 = n105_O_15_2_2; // @[Top.scala 441:12]
  assign n443_clock = clock;
  assign n443_reset = reset;
  assign n443_valid_up = n106_valid_down; // @[Top.scala 445:19]
  assign n443_I_0_0_0 = n106_O_0_0_0; // @[Top.scala 444:12]
  assign n443_I_0_0_1 = n106_O_0_0_1; // @[Top.scala 444:12]
  assign n443_I_0_0_2 = n106_O_0_0_2; // @[Top.scala 444:12]
  assign n443_I_0_1_0 = n106_O_0_1_0; // @[Top.scala 444:12]
  assign n443_I_0_1_1 = n106_O_0_1_1; // @[Top.scala 444:12]
  assign n443_I_0_1_2 = n106_O_0_1_2; // @[Top.scala 444:12]
  assign n443_I_0_2_0 = n106_O_0_2_0; // @[Top.scala 444:12]
  assign n443_I_0_2_1 = n106_O_0_2_1; // @[Top.scala 444:12]
  assign n443_I_0_2_2 = n106_O_0_2_2; // @[Top.scala 444:12]
  assign n443_I_1_0_0 = n106_O_1_0_0; // @[Top.scala 444:12]
  assign n443_I_1_0_1 = n106_O_1_0_1; // @[Top.scala 444:12]
  assign n443_I_1_0_2 = n106_O_1_0_2; // @[Top.scala 444:12]
  assign n443_I_1_1_0 = n106_O_1_1_0; // @[Top.scala 444:12]
  assign n443_I_1_1_1 = n106_O_1_1_1; // @[Top.scala 444:12]
  assign n443_I_1_1_2 = n106_O_1_1_2; // @[Top.scala 444:12]
  assign n443_I_1_2_0 = n106_O_1_2_0; // @[Top.scala 444:12]
  assign n443_I_1_2_1 = n106_O_1_2_1; // @[Top.scala 444:12]
  assign n443_I_1_2_2 = n106_O_1_2_2; // @[Top.scala 444:12]
  assign n443_I_2_0_0 = n106_O_2_0_0; // @[Top.scala 444:12]
  assign n443_I_2_0_1 = n106_O_2_0_1; // @[Top.scala 444:12]
  assign n443_I_2_0_2 = n106_O_2_0_2; // @[Top.scala 444:12]
  assign n443_I_2_1_0 = n106_O_2_1_0; // @[Top.scala 444:12]
  assign n443_I_2_1_1 = n106_O_2_1_1; // @[Top.scala 444:12]
  assign n443_I_2_1_2 = n106_O_2_1_2; // @[Top.scala 444:12]
  assign n443_I_2_2_0 = n106_O_2_2_0; // @[Top.scala 444:12]
  assign n443_I_2_2_1 = n106_O_2_2_1; // @[Top.scala 444:12]
  assign n443_I_2_2_2 = n106_O_2_2_2; // @[Top.scala 444:12]
  assign n443_I_3_0_0 = n106_O_3_0_0; // @[Top.scala 444:12]
  assign n443_I_3_0_1 = n106_O_3_0_1; // @[Top.scala 444:12]
  assign n443_I_3_0_2 = n106_O_3_0_2; // @[Top.scala 444:12]
  assign n443_I_3_1_0 = n106_O_3_1_0; // @[Top.scala 444:12]
  assign n443_I_3_1_1 = n106_O_3_1_1; // @[Top.scala 444:12]
  assign n443_I_3_1_2 = n106_O_3_1_2; // @[Top.scala 444:12]
  assign n443_I_3_2_0 = n106_O_3_2_0; // @[Top.scala 444:12]
  assign n443_I_3_2_1 = n106_O_3_2_1; // @[Top.scala 444:12]
  assign n443_I_3_2_2 = n106_O_3_2_2; // @[Top.scala 444:12]
  assign n443_I_4_0_0 = n106_O_4_0_0; // @[Top.scala 444:12]
  assign n443_I_4_0_1 = n106_O_4_0_1; // @[Top.scala 444:12]
  assign n443_I_4_0_2 = n106_O_4_0_2; // @[Top.scala 444:12]
  assign n443_I_4_1_0 = n106_O_4_1_0; // @[Top.scala 444:12]
  assign n443_I_4_1_1 = n106_O_4_1_1; // @[Top.scala 444:12]
  assign n443_I_4_1_2 = n106_O_4_1_2; // @[Top.scala 444:12]
  assign n443_I_4_2_0 = n106_O_4_2_0; // @[Top.scala 444:12]
  assign n443_I_4_2_1 = n106_O_4_2_1; // @[Top.scala 444:12]
  assign n443_I_4_2_2 = n106_O_4_2_2; // @[Top.scala 444:12]
  assign n443_I_5_0_0 = n106_O_5_0_0; // @[Top.scala 444:12]
  assign n443_I_5_0_1 = n106_O_5_0_1; // @[Top.scala 444:12]
  assign n443_I_5_0_2 = n106_O_5_0_2; // @[Top.scala 444:12]
  assign n443_I_5_1_0 = n106_O_5_1_0; // @[Top.scala 444:12]
  assign n443_I_5_1_1 = n106_O_5_1_1; // @[Top.scala 444:12]
  assign n443_I_5_1_2 = n106_O_5_1_2; // @[Top.scala 444:12]
  assign n443_I_5_2_0 = n106_O_5_2_0; // @[Top.scala 444:12]
  assign n443_I_5_2_1 = n106_O_5_2_1; // @[Top.scala 444:12]
  assign n443_I_5_2_2 = n106_O_5_2_2; // @[Top.scala 444:12]
  assign n443_I_6_0_0 = n106_O_6_0_0; // @[Top.scala 444:12]
  assign n443_I_6_0_1 = n106_O_6_0_1; // @[Top.scala 444:12]
  assign n443_I_6_0_2 = n106_O_6_0_2; // @[Top.scala 444:12]
  assign n443_I_6_1_0 = n106_O_6_1_0; // @[Top.scala 444:12]
  assign n443_I_6_1_1 = n106_O_6_1_1; // @[Top.scala 444:12]
  assign n443_I_6_1_2 = n106_O_6_1_2; // @[Top.scala 444:12]
  assign n443_I_6_2_0 = n106_O_6_2_0; // @[Top.scala 444:12]
  assign n443_I_6_2_1 = n106_O_6_2_1; // @[Top.scala 444:12]
  assign n443_I_6_2_2 = n106_O_6_2_2; // @[Top.scala 444:12]
  assign n443_I_7_0_0 = n106_O_7_0_0; // @[Top.scala 444:12]
  assign n443_I_7_0_1 = n106_O_7_0_1; // @[Top.scala 444:12]
  assign n443_I_7_0_2 = n106_O_7_0_2; // @[Top.scala 444:12]
  assign n443_I_7_1_0 = n106_O_7_1_0; // @[Top.scala 444:12]
  assign n443_I_7_1_1 = n106_O_7_1_1; // @[Top.scala 444:12]
  assign n443_I_7_1_2 = n106_O_7_1_2; // @[Top.scala 444:12]
  assign n443_I_7_2_0 = n106_O_7_2_0; // @[Top.scala 444:12]
  assign n443_I_7_2_1 = n106_O_7_2_1; // @[Top.scala 444:12]
  assign n443_I_7_2_2 = n106_O_7_2_2; // @[Top.scala 444:12]
  assign n443_I_8_0_0 = n106_O_8_0_0; // @[Top.scala 444:12]
  assign n443_I_8_0_1 = n106_O_8_0_1; // @[Top.scala 444:12]
  assign n443_I_8_0_2 = n106_O_8_0_2; // @[Top.scala 444:12]
  assign n443_I_8_1_0 = n106_O_8_1_0; // @[Top.scala 444:12]
  assign n443_I_8_1_1 = n106_O_8_1_1; // @[Top.scala 444:12]
  assign n443_I_8_1_2 = n106_O_8_1_2; // @[Top.scala 444:12]
  assign n443_I_8_2_0 = n106_O_8_2_0; // @[Top.scala 444:12]
  assign n443_I_8_2_1 = n106_O_8_2_1; // @[Top.scala 444:12]
  assign n443_I_8_2_2 = n106_O_8_2_2; // @[Top.scala 444:12]
  assign n443_I_9_0_0 = n106_O_9_0_0; // @[Top.scala 444:12]
  assign n443_I_9_0_1 = n106_O_9_0_1; // @[Top.scala 444:12]
  assign n443_I_9_0_2 = n106_O_9_0_2; // @[Top.scala 444:12]
  assign n443_I_9_1_0 = n106_O_9_1_0; // @[Top.scala 444:12]
  assign n443_I_9_1_1 = n106_O_9_1_1; // @[Top.scala 444:12]
  assign n443_I_9_1_2 = n106_O_9_1_2; // @[Top.scala 444:12]
  assign n443_I_9_2_0 = n106_O_9_2_0; // @[Top.scala 444:12]
  assign n443_I_9_2_1 = n106_O_9_2_1; // @[Top.scala 444:12]
  assign n443_I_9_2_2 = n106_O_9_2_2; // @[Top.scala 444:12]
  assign n443_I_10_0_0 = n106_O_10_0_0; // @[Top.scala 444:12]
  assign n443_I_10_0_1 = n106_O_10_0_1; // @[Top.scala 444:12]
  assign n443_I_10_0_2 = n106_O_10_0_2; // @[Top.scala 444:12]
  assign n443_I_10_1_0 = n106_O_10_1_0; // @[Top.scala 444:12]
  assign n443_I_10_1_1 = n106_O_10_1_1; // @[Top.scala 444:12]
  assign n443_I_10_1_2 = n106_O_10_1_2; // @[Top.scala 444:12]
  assign n443_I_10_2_0 = n106_O_10_2_0; // @[Top.scala 444:12]
  assign n443_I_10_2_1 = n106_O_10_2_1; // @[Top.scala 444:12]
  assign n443_I_10_2_2 = n106_O_10_2_2; // @[Top.scala 444:12]
  assign n443_I_11_0_0 = n106_O_11_0_0; // @[Top.scala 444:12]
  assign n443_I_11_0_1 = n106_O_11_0_1; // @[Top.scala 444:12]
  assign n443_I_11_0_2 = n106_O_11_0_2; // @[Top.scala 444:12]
  assign n443_I_11_1_0 = n106_O_11_1_0; // @[Top.scala 444:12]
  assign n443_I_11_1_1 = n106_O_11_1_1; // @[Top.scala 444:12]
  assign n443_I_11_1_2 = n106_O_11_1_2; // @[Top.scala 444:12]
  assign n443_I_11_2_0 = n106_O_11_2_0; // @[Top.scala 444:12]
  assign n443_I_11_2_1 = n106_O_11_2_1; // @[Top.scala 444:12]
  assign n443_I_11_2_2 = n106_O_11_2_2; // @[Top.scala 444:12]
  assign n443_I_12_0_0 = n106_O_12_0_0; // @[Top.scala 444:12]
  assign n443_I_12_0_1 = n106_O_12_0_1; // @[Top.scala 444:12]
  assign n443_I_12_0_2 = n106_O_12_0_2; // @[Top.scala 444:12]
  assign n443_I_12_1_0 = n106_O_12_1_0; // @[Top.scala 444:12]
  assign n443_I_12_1_1 = n106_O_12_1_1; // @[Top.scala 444:12]
  assign n443_I_12_1_2 = n106_O_12_1_2; // @[Top.scala 444:12]
  assign n443_I_12_2_0 = n106_O_12_2_0; // @[Top.scala 444:12]
  assign n443_I_12_2_1 = n106_O_12_2_1; // @[Top.scala 444:12]
  assign n443_I_12_2_2 = n106_O_12_2_2; // @[Top.scala 444:12]
  assign n443_I_13_0_0 = n106_O_13_0_0; // @[Top.scala 444:12]
  assign n443_I_13_0_1 = n106_O_13_0_1; // @[Top.scala 444:12]
  assign n443_I_13_0_2 = n106_O_13_0_2; // @[Top.scala 444:12]
  assign n443_I_13_1_0 = n106_O_13_1_0; // @[Top.scala 444:12]
  assign n443_I_13_1_1 = n106_O_13_1_1; // @[Top.scala 444:12]
  assign n443_I_13_1_2 = n106_O_13_1_2; // @[Top.scala 444:12]
  assign n443_I_13_2_0 = n106_O_13_2_0; // @[Top.scala 444:12]
  assign n443_I_13_2_1 = n106_O_13_2_1; // @[Top.scala 444:12]
  assign n443_I_13_2_2 = n106_O_13_2_2; // @[Top.scala 444:12]
  assign n443_I_14_0_0 = n106_O_14_0_0; // @[Top.scala 444:12]
  assign n443_I_14_0_1 = n106_O_14_0_1; // @[Top.scala 444:12]
  assign n443_I_14_0_2 = n106_O_14_0_2; // @[Top.scala 444:12]
  assign n443_I_14_1_0 = n106_O_14_1_0; // @[Top.scala 444:12]
  assign n443_I_14_1_1 = n106_O_14_1_1; // @[Top.scala 444:12]
  assign n443_I_14_1_2 = n106_O_14_1_2; // @[Top.scala 444:12]
  assign n443_I_14_2_0 = n106_O_14_2_0; // @[Top.scala 444:12]
  assign n443_I_14_2_1 = n106_O_14_2_1; // @[Top.scala 444:12]
  assign n443_I_14_2_2 = n106_O_14_2_2; // @[Top.scala 444:12]
  assign n443_I_15_0_0 = n106_O_15_0_0; // @[Top.scala 444:12]
  assign n443_I_15_0_1 = n106_O_15_0_1; // @[Top.scala 444:12]
  assign n443_I_15_0_2 = n106_O_15_0_2; // @[Top.scala 444:12]
  assign n443_I_15_1_0 = n106_O_15_1_0; // @[Top.scala 444:12]
  assign n443_I_15_1_1 = n106_O_15_1_1; // @[Top.scala 444:12]
  assign n443_I_15_1_2 = n106_O_15_1_2; // @[Top.scala 444:12]
  assign n443_I_15_2_0 = n106_O_15_2_0; // @[Top.scala 444:12]
  assign n443_I_15_2_1 = n106_O_15_2_1; // @[Top.scala 444:12]
  assign n443_I_15_2_2 = n106_O_15_2_2; // @[Top.scala 444:12]
  assign n444_valid_up = n443_valid_down; // @[Top.scala 448:19]
  assign n444_I_0_0_0_t0b = n443_O_0_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_0_0_0_t1b_t0b = n443_O_0_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_0_0_0_t1b_t1b = n443_O_0_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_1_0_0_t0b = n443_O_1_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_1_0_0_t1b_t0b = n443_O_1_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_1_0_0_t1b_t1b = n443_O_1_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_2_0_0_t0b = n443_O_2_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_2_0_0_t1b_t0b = n443_O_2_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_2_0_0_t1b_t1b = n443_O_2_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_3_0_0_t0b = n443_O_3_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_3_0_0_t1b_t0b = n443_O_3_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_3_0_0_t1b_t1b = n443_O_3_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_4_0_0_t0b = n443_O_4_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_4_0_0_t1b_t0b = n443_O_4_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_4_0_0_t1b_t1b = n443_O_4_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_5_0_0_t0b = n443_O_5_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_5_0_0_t1b_t0b = n443_O_5_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_5_0_0_t1b_t1b = n443_O_5_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_6_0_0_t0b = n443_O_6_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_6_0_0_t1b_t0b = n443_O_6_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_6_0_0_t1b_t1b = n443_O_6_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_7_0_0_t0b = n443_O_7_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_7_0_0_t1b_t0b = n443_O_7_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_7_0_0_t1b_t1b = n443_O_7_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_8_0_0_t0b = n443_O_8_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_8_0_0_t1b_t0b = n443_O_8_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_8_0_0_t1b_t1b = n443_O_8_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_9_0_0_t0b = n443_O_9_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_9_0_0_t1b_t0b = n443_O_9_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_9_0_0_t1b_t1b = n443_O_9_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_10_0_0_t0b = n443_O_10_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_10_0_0_t1b_t0b = n443_O_10_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_10_0_0_t1b_t1b = n443_O_10_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_11_0_0_t0b = n443_O_11_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_11_0_0_t1b_t0b = n443_O_11_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_11_0_0_t1b_t1b = n443_O_11_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_12_0_0_t0b = n443_O_12_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_12_0_0_t1b_t0b = n443_O_12_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_12_0_0_t1b_t1b = n443_O_12_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_13_0_0_t0b = n443_O_13_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_13_0_0_t1b_t0b = n443_O_13_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_13_0_0_t1b_t1b = n443_O_13_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_14_0_0_t0b = n443_O_14_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_14_0_0_t1b_t0b = n443_O_14_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_14_0_0_t1b_t1b = n443_O_14_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n444_I_15_0_0_t0b = n443_O_15_0_0_t0b; // @[Top.scala 447:12]
  assign n444_I_15_0_0_t1b_t0b = n443_O_15_0_0_t1b_t0b; // @[Top.scala 447:12]
  assign n444_I_15_0_0_t1b_t1b = n443_O_15_0_0_t1b_t1b; // @[Top.scala 447:12]
  assign n445_valid_up = n444_valid_down; // @[Top.scala 451:19]
  assign n445_I_0_0_0_t0b = n444_O_0_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_0_0_0_t1b_t0b = n444_O_0_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_0_0_0_t1b_t1b = n444_O_0_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_1_0_0_t0b = n444_O_1_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_1_0_0_t1b_t0b = n444_O_1_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_1_0_0_t1b_t1b = n444_O_1_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_2_0_0_t0b = n444_O_2_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_2_0_0_t1b_t0b = n444_O_2_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_2_0_0_t1b_t1b = n444_O_2_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_3_0_0_t0b = n444_O_3_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_3_0_0_t1b_t0b = n444_O_3_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_3_0_0_t1b_t1b = n444_O_3_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_4_0_0_t0b = n444_O_4_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_4_0_0_t1b_t0b = n444_O_4_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_4_0_0_t1b_t1b = n444_O_4_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_5_0_0_t0b = n444_O_5_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_5_0_0_t1b_t0b = n444_O_5_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_5_0_0_t1b_t1b = n444_O_5_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_6_0_0_t0b = n444_O_6_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_6_0_0_t1b_t0b = n444_O_6_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_6_0_0_t1b_t1b = n444_O_6_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_7_0_0_t0b = n444_O_7_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_7_0_0_t1b_t0b = n444_O_7_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_7_0_0_t1b_t1b = n444_O_7_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_8_0_0_t0b = n444_O_8_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_8_0_0_t1b_t0b = n444_O_8_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_8_0_0_t1b_t1b = n444_O_8_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_9_0_0_t0b = n444_O_9_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_9_0_0_t1b_t0b = n444_O_9_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_9_0_0_t1b_t1b = n444_O_9_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_10_0_0_t0b = n444_O_10_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_10_0_0_t1b_t0b = n444_O_10_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_10_0_0_t1b_t1b = n444_O_10_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_11_0_0_t0b = n444_O_11_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_11_0_0_t1b_t0b = n444_O_11_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_11_0_0_t1b_t1b = n444_O_11_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_12_0_0_t0b = n444_O_12_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_12_0_0_t1b_t0b = n444_O_12_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_12_0_0_t1b_t1b = n444_O_12_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_13_0_0_t0b = n444_O_13_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_13_0_0_t1b_t0b = n444_O_13_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_13_0_0_t1b_t1b = n444_O_13_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_14_0_0_t0b = n444_O_14_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_14_0_0_t1b_t0b = n444_O_14_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_14_0_0_t1b_t1b = n444_O_14_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n445_I_15_0_0_t0b = n444_O_15_0_0_t0b; // @[Top.scala 450:12]
  assign n445_I_15_0_0_t1b_t0b = n444_O_15_0_0_t1b_t0b; // @[Top.scala 450:12]
  assign n445_I_15_0_0_t1b_t1b = n444_O_15_0_0_t1b_t1b; // @[Top.scala 450:12]
  assign n446_valid_up = n445_valid_down; // @[Top.scala 454:19]
  assign n446_I_0_0_t0b = n445_O_0_0_t0b; // @[Top.scala 453:12]
  assign n446_I_0_0_t1b_t0b = n445_O_0_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_0_0_t1b_t1b = n445_O_0_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_1_0_t0b = n445_O_1_0_t0b; // @[Top.scala 453:12]
  assign n446_I_1_0_t1b_t0b = n445_O_1_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_1_0_t1b_t1b = n445_O_1_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_2_0_t0b = n445_O_2_0_t0b; // @[Top.scala 453:12]
  assign n446_I_2_0_t1b_t0b = n445_O_2_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_2_0_t1b_t1b = n445_O_2_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_3_0_t0b = n445_O_3_0_t0b; // @[Top.scala 453:12]
  assign n446_I_3_0_t1b_t0b = n445_O_3_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_3_0_t1b_t1b = n445_O_3_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_4_0_t0b = n445_O_4_0_t0b; // @[Top.scala 453:12]
  assign n446_I_4_0_t1b_t0b = n445_O_4_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_4_0_t1b_t1b = n445_O_4_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_5_0_t0b = n445_O_5_0_t0b; // @[Top.scala 453:12]
  assign n446_I_5_0_t1b_t0b = n445_O_5_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_5_0_t1b_t1b = n445_O_5_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_6_0_t0b = n445_O_6_0_t0b; // @[Top.scala 453:12]
  assign n446_I_6_0_t1b_t0b = n445_O_6_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_6_0_t1b_t1b = n445_O_6_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_7_0_t0b = n445_O_7_0_t0b; // @[Top.scala 453:12]
  assign n446_I_7_0_t1b_t0b = n445_O_7_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_7_0_t1b_t1b = n445_O_7_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_8_0_t0b = n445_O_8_0_t0b; // @[Top.scala 453:12]
  assign n446_I_8_0_t1b_t0b = n445_O_8_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_8_0_t1b_t1b = n445_O_8_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_9_0_t0b = n445_O_9_0_t0b; // @[Top.scala 453:12]
  assign n446_I_9_0_t1b_t0b = n445_O_9_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_9_0_t1b_t1b = n445_O_9_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_10_0_t0b = n445_O_10_0_t0b; // @[Top.scala 453:12]
  assign n446_I_10_0_t1b_t0b = n445_O_10_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_10_0_t1b_t1b = n445_O_10_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_11_0_t0b = n445_O_11_0_t0b; // @[Top.scala 453:12]
  assign n446_I_11_0_t1b_t0b = n445_O_11_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_11_0_t1b_t1b = n445_O_11_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_12_0_t0b = n445_O_12_0_t0b; // @[Top.scala 453:12]
  assign n446_I_12_0_t1b_t0b = n445_O_12_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_12_0_t1b_t1b = n445_O_12_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_13_0_t0b = n445_O_13_0_t0b; // @[Top.scala 453:12]
  assign n446_I_13_0_t1b_t0b = n445_O_13_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_13_0_t1b_t1b = n445_O_13_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_14_0_t0b = n445_O_14_0_t0b; // @[Top.scala 453:12]
  assign n446_I_14_0_t1b_t0b = n445_O_14_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_14_0_t1b_t1b = n445_O_14_0_t1b_t1b; // @[Top.scala 453:12]
  assign n446_I_15_0_t0b = n445_O_15_0_t0b; // @[Top.scala 453:12]
  assign n446_I_15_0_t1b_t0b = n445_O_15_0_t1b_t0b; // @[Top.scala 453:12]
  assign n446_I_15_0_t1b_t1b = n445_O_15_0_t1b_t1b; // @[Top.scala 453:12]
  assign n447_clock = clock;
  assign n447_reset = reset;
  assign n447_valid_up = n446_valid_down; // @[Top.scala 457:19]
  assign n447_I_0_t0b = n446_O_0_t0b; // @[Top.scala 456:12]
  assign n447_I_0_t1b_t0b = n446_O_0_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_0_t1b_t1b = n446_O_0_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_1_t0b = n446_O_1_t0b; // @[Top.scala 456:12]
  assign n447_I_1_t1b_t0b = n446_O_1_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_1_t1b_t1b = n446_O_1_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_2_t0b = n446_O_2_t0b; // @[Top.scala 456:12]
  assign n447_I_2_t1b_t0b = n446_O_2_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_2_t1b_t1b = n446_O_2_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_3_t0b = n446_O_3_t0b; // @[Top.scala 456:12]
  assign n447_I_3_t1b_t0b = n446_O_3_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_3_t1b_t1b = n446_O_3_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_4_t0b = n446_O_4_t0b; // @[Top.scala 456:12]
  assign n447_I_4_t1b_t0b = n446_O_4_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_4_t1b_t1b = n446_O_4_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_5_t0b = n446_O_5_t0b; // @[Top.scala 456:12]
  assign n447_I_5_t1b_t0b = n446_O_5_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_5_t1b_t1b = n446_O_5_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_6_t0b = n446_O_6_t0b; // @[Top.scala 456:12]
  assign n447_I_6_t1b_t0b = n446_O_6_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_6_t1b_t1b = n446_O_6_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_7_t0b = n446_O_7_t0b; // @[Top.scala 456:12]
  assign n447_I_7_t1b_t0b = n446_O_7_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_7_t1b_t1b = n446_O_7_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_8_t0b = n446_O_8_t0b; // @[Top.scala 456:12]
  assign n447_I_8_t1b_t0b = n446_O_8_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_8_t1b_t1b = n446_O_8_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_9_t0b = n446_O_9_t0b; // @[Top.scala 456:12]
  assign n447_I_9_t1b_t0b = n446_O_9_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_9_t1b_t1b = n446_O_9_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_10_t0b = n446_O_10_t0b; // @[Top.scala 456:12]
  assign n447_I_10_t1b_t0b = n446_O_10_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_10_t1b_t1b = n446_O_10_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_11_t0b = n446_O_11_t0b; // @[Top.scala 456:12]
  assign n447_I_11_t1b_t0b = n446_O_11_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_11_t1b_t1b = n446_O_11_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_12_t0b = n446_O_12_t0b; // @[Top.scala 456:12]
  assign n447_I_12_t1b_t0b = n446_O_12_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_12_t1b_t1b = n446_O_12_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_13_t0b = n446_O_13_t0b; // @[Top.scala 456:12]
  assign n447_I_13_t1b_t0b = n446_O_13_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_13_t1b_t1b = n446_O_13_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_14_t0b = n446_O_14_t0b; // @[Top.scala 456:12]
  assign n447_I_14_t1b_t0b = n446_O_14_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_14_t1b_t1b = n446_O_14_t1b_t1b; // @[Top.scala 456:12]
  assign n447_I_15_t0b = n446_O_15_t0b; // @[Top.scala 456:12]
  assign n447_I_15_t1b_t0b = n446_O_15_t1b_t0b; // @[Top.scala 456:12]
  assign n447_I_15_t1b_t1b = n446_O_15_t1b_t1b; // @[Top.scala 456:12]
  assign n448_clock = clock;
  assign n448_reset = reset;
  assign n448_valid_up = n447_valid_down; // @[Top.scala 460:19]
  assign n448_I_0_t0b = n447_O_0_t0b; // @[Top.scala 459:12]
  assign n448_I_0_t1b_t0b = n447_O_0_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_0_t1b_t1b = n447_O_0_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_1_t0b = n447_O_1_t0b; // @[Top.scala 459:12]
  assign n448_I_1_t1b_t0b = n447_O_1_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_1_t1b_t1b = n447_O_1_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_2_t0b = n447_O_2_t0b; // @[Top.scala 459:12]
  assign n448_I_2_t1b_t0b = n447_O_2_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_2_t1b_t1b = n447_O_2_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_3_t0b = n447_O_3_t0b; // @[Top.scala 459:12]
  assign n448_I_3_t1b_t0b = n447_O_3_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_3_t1b_t1b = n447_O_3_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_4_t0b = n447_O_4_t0b; // @[Top.scala 459:12]
  assign n448_I_4_t1b_t0b = n447_O_4_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_4_t1b_t1b = n447_O_4_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_5_t0b = n447_O_5_t0b; // @[Top.scala 459:12]
  assign n448_I_5_t1b_t0b = n447_O_5_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_5_t1b_t1b = n447_O_5_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_6_t0b = n447_O_6_t0b; // @[Top.scala 459:12]
  assign n448_I_6_t1b_t0b = n447_O_6_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_6_t1b_t1b = n447_O_6_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_7_t0b = n447_O_7_t0b; // @[Top.scala 459:12]
  assign n448_I_7_t1b_t0b = n447_O_7_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_7_t1b_t1b = n447_O_7_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_8_t0b = n447_O_8_t0b; // @[Top.scala 459:12]
  assign n448_I_8_t1b_t0b = n447_O_8_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_8_t1b_t1b = n447_O_8_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_9_t0b = n447_O_9_t0b; // @[Top.scala 459:12]
  assign n448_I_9_t1b_t0b = n447_O_9_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_9_t1b_t1b = n447_O_9_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_10_t0b = n447_O_10_t0b; // @[Top.scala 459:12]
  assign n448_I_10_t1b_t0b = n447_O_10_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_10_t1b_t1b = n447_O_10_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_11_t0b = n447_O_11_t0b; // @[Top.scala 459:12]
  assign n448_I_11_t1b_t0b = n447_O_11_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_11_t1b_t1b = n447_O_11_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_12_t0b = n447_O_12_t0b; // @[Top.scala 459:12]
  assign n448_I_12_t1b_t0b = n447_O_12_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_12_t1b_t1b = n447_O_12_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_13_t0b = n447_O_13_t0b; // @[Top.scala 459:12]
  assign n448_I_13_t1b_t0b = n447_O_13_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_13_t1b_t1b = n447_O_13_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_14_t0b = n447_O_14_t0b; // @[Top.scala 459:12]
  assign n448_I_14_t1b_t0b = n447_O_14_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_14_t1b_t1b = n447_O_14_t1b_t1b; // @[Top.scala 459:12]
  assign n448_I_15_t0b = n447_O_15_t0b; // @[Top.scala 459:12]
  assign n448_I_15_t1b_t0b = n447_O_15_t1b_t0b; // @[Top.scala 459:12]
  assign n448_I_15_t1b_t1b = n447_O_15_t1b_t1b; // @[Top.scala 459:12]
  assign n449_clock = clock;
  assign n449_reset = reset;
  assign n449_valid_up = n448_valid_down; // @[Top.scala 463:19]
  assign n449_I_0_t0b = n448_O_0_t0b; // @[Top.scala 462:12]
  assign n449_I_0_t1b_t0b = n448_O_0_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_0_t1b_t1b = n448_O_0_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_1_t0b = n448_O_1_t0b; // @[Top.scala 462:12]
  assign n449_I_1_t1b_t0b = n448_O_1_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_1_t1b_t1b = n448_O_1_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_2_t0b = n448_O_2_t0b; // @[Top.scala 462:12]
  assign n449_I_2_t1b_t0b = n448_O_2_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_2_t1b_t1b = n448_O_2_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_3_t0b = n448_O_3_t0b; // @[Top.scala 462:12]
  assign n449_I_3_t1b_t0b = n448_O_3_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_3_t1b_t1b = n448_O_3_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_4_t0b = n448_O_4_t0b; // @[Top.scala 462:12]
  assign n449_I_4_t1b_t0b = n448_O_4_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_4_t1b_t1b = n448_O_4_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_5_t0b = n448_O_5_t0b; // @[Top.scala 462:12]
  assign n449_I_5_t1b_t0b = n448_O_5_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_5_t1b_t1b = n448_O_5_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_6_t0b = n448_O_6_t0b; // @[Top.scala 462:12]
  assign n449_I_6_t1b_t0b = n448_O_6_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_6_t1b_t1b = n448_O_6_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_7_t0b = n448_O_7_t0b; // @[Top.scala 462:12]
  assign n449_I_7_t1b_t0b = n448_O_7_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_7_t1b_t1b = n448_O_7_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_8_t0b = n448_O_8_t0b; // @[Top.scala 462:12]
  assign n449_I_8_t1b_t0b = n448_O_8_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_8_t1b_t1b = n448_O_8_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_9_t0b = n448_O_9_t0b; // @[Top.scala 462:12]
  assign n449_I_9_t1b_t0b = n448_O_9_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_9_t1b_t1b = n448_O_9_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_10_t0b = n448_O_10_t0b; // @[Top.scala 462:12]
  assign n449_I_10_t1b_t0b = n448_O_10_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_10_t1b_t1b = n448_O_10_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_11_t0b = n448_O_11_t0b; // @[Top.scala 462:12]
  assign n449_I_11_t1b_t0b = n448_O_11_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_11_t1b_t1b = n448_O_11_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_12_t0b = n448_O_12_t0b; // @[Top.scala 462:12]
  assign n449_I_12_t1b_t0b = n448_O_12_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_12_t1b_t1b = n448_O_12_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_13_t0b = n448_O_13_t0b; // @[Top.scala 462:12]
  assign n449_I_13_t1b_t0b = n448_O_13_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_13_t1b_t1b = n448_O_13_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_14_t0b = n448_O_14_t0b; // @[Top.scala 462:12]
  assign n449_I_14_t1b_t0b = n448_O_14_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_14_t1b_t1b = n448_O_14_t1b_t1b; // @[Top.scala 462:12]
  assign n449_I_15_t0b = n448_O_15_t0b; // @[Top.scala 462:12]
  assign n449_I_15_t1b_t0b = n448_O_15_t1b_t0b; // @[Top.scala 462:12]
  assign n449_I_15_t1b_t1b = n448_O_15_t1b_t1b; // @[Top.scala 462:12]
endmodule
