module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  output [31:0] O_0,
  output [31:0] O_1
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x266_TREADY(dontcare), // @[:@1298.4]
    .io_in_x266_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x266_TID(8'h0),
    .io_in_x266_TDEST(8'h0),
    .io_in_x267_TVALID(valid_down), // @[:@1298.4]
    .io_in_x267_TDATA({O_0,O_1}), // @[:@1298.4]
    .io_in_x267_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x274_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule

module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh25); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh25); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x268_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x542_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x471_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x269_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x270_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x274_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x290_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x520_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x280_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x290_inr_Foreach_kernelx290_inr_Foreach_concrete1( // @[:@4748.2]
  input         clock, // @[:@4749.4]
  input         reset, // @[:@4750.4]
  output        io_in_x270_fifoinpacked_0_wPort_0_en_0, // @[:@4751.4]
  input         io_in_x270_fifoinpacked_0_full, // @[:@4751.4]
  output        io_in_x270_fifoinpacked_0_active_0_in, // @[:@4751.4]
  input         io_in_x270_fifoinpacked_0_active_0_out, // @[:@4751.4]
  input         io_sigsIn_backpressure, // @[:@4751.4]
  input         io_sigsIn_datapathEn, // @[:@4751.4]
  input         io_sigsIn_break, // @[:@4751.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4751.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4751.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4751.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4751.4]
  input         io_rr // @[:@4751.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4785.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4785.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4797.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@4797.4]
  wire  x520_sub_1_clock; // @[Math.scala 191:24:@4824.4]
  wire  x520_sub_1_reset; // @[Math.scala 191:24:@4824.4]
  wire [31:0] x520_sub_1_io_a; // @[Math.scala 191:24:@4824.4]
  wire [31:0] x520_sub_1_io_b; // @[Math.scala 191:24:@4824.4]
  wire  x520_sub_1_io_flow; // @[Math.scala 191:24:@4824.4]
  wire [31:0] x520_sub_1_io_result; // @[Math.scala 191:24:@4824.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4834.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4834.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4834.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4834.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4834.4]
  wire  x280_sum_1_clock; // @[Math.scala 150:24:@4843.4]
  wire  x280_sum_1_reset; // @[Math.scala 150:24:@4843.4]
  wire [31:0] x280_sum_1_io_a; // @[Math.scala 150:24:@4843.4]
  wire [31:0] x280_sum_1_io_b; // @[Math.scala 150:24:@4843.4]
  wire  x280_sum_1_io_flow; // @[Math.scala 150:24:@4843.4]
  wire [31:0] x280_sum_1_io_result; // @[Math.scala 150:24:@4843.4]
  wire  x281_sum_1_clock; // @[Math.scala 150:24:@4855.4]
  wire  x281_sum_1_reset; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x281_sum_1_io_a; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x281_sum_1_io_b; // @[Math.scala 150:24:@4855.4]
  wire  x281_sum_1_io_flow; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x281_sum_1_io_result; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x283_1_io_b; // @[Math.scala 720:24:@4876.4]
  wire [31:0] x283_1_io_result; // @[Math.scala 720:24:@4876.4]
  wire  x284_sum_1_clock; // @[Math.scala 150:24:@4887.4]
  wire  x284_sum_1_reset; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x284_sum_1_io_a; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x284_sum_1_io_b; // @[Math.scala 150:24:@4887.4]
  wire  x284_sum_1_io_flow; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x284_sum_1_io_result; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x286_1_io_b; // @[Math.scala 720:24:@4908.4]
  wire [31:0] x286_1_io_result; // @[Math.scala 720:24:@4908.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4943.4]
  wire  _T_327; // @[sm_x290_inr_Foreach.scala 62:18:@4810.4]
  wire  _T_328; // @[sm_x290_inr_Foreach.scala 62:55:@4811.4]
  wire [31:0] b275_number; // @[Math.scala 723:22:@4790.4 Math.scala 724:14:@4791.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@4815.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@4815.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@4820.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@4820.4]
  wire [31:0] x281_sum_number; // @[Math.scala 154:22:@4861.4 Math.scala 155:14:@4862.4]
  wire [31:0] _T_358; // @[Math.scala 406:49:@4868.4]
  wire [31:0] _T_360; // @[Math.scala 406:56:@4870.4]
  wire [31:0] _T_361; // @[Math.scala 406:56:@4871.4]
  wire [31:0] x284_sum_number; // @[Math.scala 154:22:@4893.4 Math.scala 155:14:@4894.4]
  wire [31:0] _T_380; // @[Math.scala 406:49:@4900.4]
  wire [31:0] _T_382; // @[Math.scala 406:56:@4902.4]
  wire [31:0] _T_383; // @[Math.scala 406:56:@4903.4]
  wire  _T_403; // @[sm_x290_inr_Foreach.scala 95:131:@4940.4]
  wire  _T_407; // @[package.scala 96:25:@4948.4 package.scala 96:25:@4949.4]
  wire  _T_409; // @[implicits.scala 55:10:@4950.4]
  wire  _T_410; // @[sm_x290_inr_Foreach.scala 95:148:@4951.4]
  wire  _T_412; // @[sm_x290_inr_Foreach.scala 95:236:@4953.4]
  wire  _T_413; // @[sm_x290_inr_Foreach.scala 95:255:@4954.4]
  wire  x545_b277_D3; // @[package.scala 96:25:@4928.4 package.scala 96:25:@4929.4]
  wire  _T_416; // @[sm_x290_inr_Foreach.scala 95:291:@4956.4]
  wire  x546_b278_D3; // @[package.scala 96:25:@4937.4 package.scala 96:25:@4938.4]
  _ _ ( // @[Math.scala 720:24:@4785.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@4797.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x520_sub x520_sub_1 ( // @[Math.scala 191:24:@4824.4]
    .clock(x520_sub_1_clock),
    .reset(x520_sub_1_reset),
    .io_a(x520_sub_1_io_a),
    .io_b(x520_sub_1_io_b),
    .io_flow(x520_sub_1_io_flow),
    .io_result(x520_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4834.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x280_sum x280_sum_1 ( // @[Math.scala 150:24:@4843.4]
    .clock(x280_sum_1_clock),
    .reset(x280_sum_1_reset),
    .io_a(x280_sum_1_io_a),
    .io_b(x280_sum_1_io_b),
    .io_flow(x280_sum_1_io_flow),
    .io_result(x280_sum_1_io_result)
  );
  x280_sum x281_sum_1 ( // @[Math.scala 150:24:@4855.4]
    .clock(x281_sum_1_clock),
    .reset(x281_sum_1_reset),
    .io_a(x281_sum_1_io_a),
    .io_b(x281_sum_1_io_b),
    .io_flow(x281_sum_1_io_flow),
    .io_result(x281_sum_1_io_result)
  );
  _ x283_1 ( // @[Math.scala 720:24:@4876.4]
    .io_b(x283_1_io_b),
    .io_result(x283_1_io_result)
  );
  x280_sum x284_sum_1 ( // @[Math.scala 150:24:@4887.4]
    .clock(x284_sum_1_clock),
    .reset(x284_sum_1_reset),
    .io_a(x284_sum_1_io_a),
    .io_b(x284_sum_1_io_b),
    .io_flow(x284_sum_1_io_flow),
    .io_result(x284_sum_1_io_result)
  );
  _ x286_1 ( // @[Math.scala 720:24:@4908.4]
    .io_b(x286_1_io_b),
    .io_result(x286_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4923.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4932.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4943.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x270_fifoinpacked_0_full; // @[sm_x290_inr_Foreach.scala 62:18:@4810.4]
  assign _T_328 = ~ io_in_x270_fifoinpacked_0_active_0_out; // @[sm_x290_inr_Foreach.scala 62:55:@4811.4]
  assign b275_number = __io_result; // @[Math.scala 723:22:@4790.4 Math.scala 724:14:@4791.4]
  assign _GEN_0 = {{11'd0}, b275_number}; // @[Math.scala 461:32:@4815.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@4815.4]
  assign _GEN_1 = {{7'd0}, b275_number}; // @[Math.scala 461:32:@4820.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@4820.4]
  assign x281_sum_number = x281_sum_1_io_result; // @[Math.scala 154:22:@4861.4 Math.scala 155:14:@4862.4]
  assign _T_358 = $signed(x281_sum_number); // @[Math.scala 406:49:@4868.4]
  assign _T_360 = $signed(_T_358) & $signed(32'shff); // @[Math.scala 406:56:@4870.4]
  assign _T_361 = $signed(_T_360); // @[Math.scala 406:56:@4871.4]
  assign x284_sum_number = x284_sum_1_io_result; // @[Math.scala 154:22:@4893.4 Math.scala 155:14:@4894.4]
  assign _T_380 = $signed(x284_sum_number); // @[Math.scala 406:49:@4900.4]
  assign _T_382 = $signed(_T_380) & $signed(32'shff); // @[Math.scala 406:56:@4902.4]
  assign _T_383 = $signed(_T_382); // @[Math.scala 406:56:@4903.4]
  assign _T_403 = ~ io_sigsIn_break; // @[sm_x290_inr_Foreach.scala 95:131:@4940.4]
  assign _T_407 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4948.4 package.scala 96:25:@4949.4]
  assign _T_409 = io_rr ? _T_407 : 1'h0; // @[implicits.scala 55:10:@4950.4]
  assign _T_410 = _T_403 & _T_409; // @[sm_x290_inr_Foreach.scala 95:148:@4951.4]
  assign _T_412 = _T_410 & _T_403; // @[sm_x290_inr_Foreach.scala 95:236:@4953.4]
  assign _T_413 = _T_412 & io_sigsIn_backpressure; // @[sm_x290_inr_Foreach.scala 95:255:@4954.4]
  assign x545_b277_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4928.4 package.scala 96:25:@4929.4]
  assign _T_416 = _T_413 & x545_b277_D3; // @[sm_x290_inr_Foreach.scala 95:291:@4956.4]
  assign x546_b278_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4937.4 package.scala 96:25:@4938.4]
  assign io_in_x270_fifoinpacked_0_wPort_0_en_0 = _T_416 & x546_b278_D3; // @[MemInterfaceType.scala 93:57:@4960.4]
  assign io_in_x270_fifoinpacked_0_active_0_in = x545_b277_D3 & x546_b278_D3; // @[MemInterfaceType.scala 147:18:@4963.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4788.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@4800.4]
  assign x520_sub_1_clock = clock; // @[:@4825.4]
  assign x520_sub_1_reset = reset; // @[:@4826.4]
  assign x520_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@4827.4]
  assign x520_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@4828.4]
  assign x520_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4829.4]
  assign RetimeWrapper_clock = clock; // @[:@4835.4]
  assign RetimeWrapper_reset = reset; // @[:@4836.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4838.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4837.4]
  assign x280_sum_1_clock = clock; // @[:@4844.4]
  assign x280_sum_1_reset = reset; // @[:@4845.4]
  assign x280_sum_1_io_a = x520_sub_1_io_result; // @[Math.scala 151:17:@4846.4]
  assign x280_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4847.4]
  assign x280_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4848.4]
  assign x281_sum_1_clock = clock; // @[:@4856.4]
  assign x281_sum_1_reset = reset; // @[:@4857.4]
  assign x281_sum_1_io_a = x280_sum_1_io_result; // @[Math.scala 151:17:@4858.4]
  assign x281_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4859.4]
  assign x281_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4860.4]
  assign x283_1_io_b = $unsigned(_T_361); // @[Math.scala 721:17:@4879.4]
  assign x284_sum_1_clock = clock; // @[:@4888.4]
  assign x284_sum_1_reset = reset; // @[:@4889.4]
  assign x284_sum_1_io_a = x280_sum_1_io_result; // @[Math.scala 151:17:@4890.4]
  assign x284_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@4891.4]
  assign x284_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4892.4]
  assign x286_1_io_b = $unsigned(_T_383); // @[Math.scala 721:17:@4911.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4924.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4925.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4927.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4926.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4933.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4934.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4936.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4935.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4944.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4945.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4947.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4946.4]
endmodule
module RetimeWrapper_42( // @[:@6081.2]
  input   clock, // @[:@6082.4]
  input   reset, // @[:@6083.4]
  input   io_flow, // @[:@6084.4]
  input   io_in, // @[:@6084.4]
  output  io_out // @[:@6084.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(74)) sr ( // @[RetimeShiftRegister.scala 15:20:@6086.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6099.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6098.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6097.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6096.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6095.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6093.4]
endmodule
module RetimeWrapper_46( // @[:@6209.2]
  input   clock, // @[:@6210.4]
  input   reset, // @[:@6211.4]
  input   io_flow, // @[:@6212.4]
  input   io_in, // @[:@6212.4]
  output  io_out // @[:@6212.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(73)) sr ( // @[RetimeShiftRegister.scala 15:20:@6214.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6227.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6226.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6225.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6224.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6223.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6221.4]
endmodule
module x469_inr_Foreach_SAMPLER_BOX_sm( // @[:@6229.2]
  input   clock, // @[:@6230.4]
  input   reset, // @[:@6231.4]
  input   io_enable, // @[:@6232.4]
  output  io_done, // @[:@6232.4]
  output  io_doneLatch, // @[:@6232.4]
  input   io_ctrDone, // @[:@6232.4]
  output  io_datapathEn, // @[:@6232.4]
  output  io_ctrInc, // @[:@6232.4]
  output  io_ctrRst, // @[:@6232.4]
  input   io_parentAck, // @[:@6232.4]
  input   io_backpressure, // @[:@6232.4]
  input   io_break // @[:@6232.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6234.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6234.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6237.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6237.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6329.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6242.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6243.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6244.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6245.4]
  wire  _T_100; // @[package.scala 100:49:@6262.4]
  reg  _T_103; // @[package.scala 48:56:@6263.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6276.4 package.scala 96:25:@6277.4]
  wire  _T_110; // @[package.scala 100:49:@6278.4]
  reg  _T_113; // @[package.scala 48:56:@6279.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6281.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6286.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6287.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6290.4]
  wire  _T_124; // @[package.scala 96:25:@6298.4 package.scala 96:25:@6299.4]
  wire  _T_126; // @[package.scala 100:49:@6300.4]
  reg  _T_129; // @[package.scala 48:56:@6301.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6323.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6325.4]
  reg  _T_153; // @[package.scala 48:56:@6326.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6334.4 package.scala 96:25:@6335.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6336.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6337.4]
  SRFF active ( // @[Controllers.scala 261:22:@6234.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6237.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_42 RetimeWrapper ( // @[package.scala 93:22:@6271.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_1 ( // @[package.scala 93:22:@6293.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6305.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6313.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_4 ( // @[package.scala 93:22:@6329.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6242.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6243.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6244.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6245.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6262.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6276.4 package.scala 96:25:@6277.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6278.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6281.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6286.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6287.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6290.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6298.4 package.scala 96:25:@6299.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6300.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6325.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6334.4 package.scala 96:25:@6335.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6336.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6337.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6304.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6339.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6289.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6292.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6284.4]
  assign active_clock = clock; // @[:@6235.4]
  assign active_reset = reset; // @[:@6236.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6247.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6251.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6252.4]
  assign done_clock = clock; // @[:@6238.4]
  assign done_reset = reset; // @[:@6239.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6267.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6260.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6261.4]
  assign RetimeWrapper_clock = clock; // @[:@6272.4]
  assign RetimeWrapper_reset = reset; // @[:@6273.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6275.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6274.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6294.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6295.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6297.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6296.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6306.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6307.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6309.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6308.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6314.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6315.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6317.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6316.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6330.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6331.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6333.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6332.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_50( // @[:@6530.2]
  input         clock, // @[:@6531.4]
  input         reset, // @[:@6532.4]
  input         io_flow, // @[:@6533.4]
  input  [63:0] io_in, // @[:@6533.4]
  output [63:0] io_out // @[:@6533.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6535.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6548.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6547.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@6546.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6545.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6544.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6542.4]
endmodule
module SRAM_1( // @[:@6566.2]
  input         clock, // @[:@6567.4]
  input         reset, // @[:@6568.4]
  input  [8:0]  io_raddr, // @[:@6569.4]
  input         io_wen, // @[:@6569.4]
  input  [8:0]  io_waddr, // @[:@6569.4]
  input  [31:0] io_wdata, // @[:@6569.4]
  output [31:0] io_rdata, // @[:@6569.4]
  input         io_backpressure // @[:@6569.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6571.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6571.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6571.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6571.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6589.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6590.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6591.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6593.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(480), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6571.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6589.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6590.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6598.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6585.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6586.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6583.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6588.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6587.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6584.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6582.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6581.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_51( // @[:@6612.2]
  input        clock, // @[:@6613.4]
  input        reset, // @[:@6614.4]
  input        io_flow, // @[:@6615.4]
  input  [8:0] io_in, // @[:@6615.4]
  output [8:0] io_out // @[:@6615.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6617.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6630.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6629.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@6628.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6627.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6626.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6624.4]
endmodule
module Mem1D_5( // @[:@6632.2]
  input         clock, // @[:@6633.4]
  input         reset, // @[:@6634.4]
  input  [8:0]  io_r_ofs_0, // @[:@6635.4]
  input         io_r_backpressure, // @[:@6635.4]
  input  [8:0]  io_w_ofs_0, // @[:@6635.4]
  input  [31:0] io_w_data_0, // @[:@6635.4]
  input         io_w_en_0, // @[:@6635.4]
  output [31:0] io_output // @[:@6635.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6642.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6642.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6642.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6642.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6642.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@6637.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@6639.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_51 RetimeWrapper ( // @[package.scala 93:22:@6642.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h1e0; // @[MemPrimitives.scala 702:32:@6637.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@6655.4]
  assign SRAM_clock = clock; // @[:@6640.4]
  assign SRAM_reset = reset; // @[:@6641.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@6649.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@6652.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@6650.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@6653.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@6654.4]
  assign RetimeWrapper_clock = clock; // @[:@6643.4]
  assign RetimeWrapper_reset = reset; // @[:@6644.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6646.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6645.4]
endmodule
module StickySelects_1( // @[:@8262.2]
  input   clock, // @[:@8263.4]
  input   reset, // @[:@8264.4]
  input   io_ins_0, // @[:@8265.4]
  input   io_ins_1, // @[:@8265.4]
  input   io_ins_2, // @[:@8265.4]
  input   io_ins_3, // @[:@8265.4]
  input   io_ins_4, // @[:@8265.4]
  input   io_ins_5, // @[:@8265.4]
  output  io_outs_0, // @[:@8265.4]
  output  io_outs_1, // @[:@8265.4]
  output  io_outs_2, // @[:@8265.4]
  output  io_outs_3, // @[:@8265.4]
  output  io_outs_4, // @[:@8265.4]
  output  io_outs_5 // @[:@8265.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@8267.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@8268.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@8269.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@8270.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@8271.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@8272.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@8273.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@8274.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@8275.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@8276.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@8277.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@8278.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@8280.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@8281.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@8282.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@8283.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@8284.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@8285.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@8287.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@8288.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@8289.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@8290.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@8291.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@8292.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@8295.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@8296.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@8297.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@8298.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@8299.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@8303.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@8304.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@8305.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@8306.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@8311.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@8312.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@8313.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@8273.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@8274.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@8275.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@8276.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@8277.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@8278.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@8280.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@8281.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@8282.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@8283.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@8284.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@8285.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@8287.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@8288.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@8289.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@8290.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@8291.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@8292.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@8295.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@8296.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@8297.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@8298.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@8299.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@8303.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@8304.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@8305.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@8306.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@8311.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@8312.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@8313.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@8315.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@8316.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@8317.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@8318.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@8319.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@8320.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x301_lb_0( // @[:@12294.2]
  input         clock, // @[:@12295.4]
  input         reset, // @[:@12296.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@12297.4]
  input         io_rPort_11_en_0, // @[:@12297.4]
  input         io_rPort_11_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_11_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@12297.4]
  input         io_rPort_10_en_0, // @[:@12297.4]
  input         io_rPort_10_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_10_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@12297.4]
  input         io_rPort_9_en_0, // @[:@12297.4]
  input         io_rPort_9_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_9_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@12297.4]
  input         io_rPort_8_en_0, // @[:@12297.4]
  input         io_rPort_8_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_8_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@12297.4]
  input         io_rPort_7_en_0, // @[:@12297.4]
  input         io_rPort_7_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_7_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@12297.4]
  input         io_rPort_6_en_0, // @[:@12297.4]
  input         io_rPort_6_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_6_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@12297.4]
  input         io_rPort_5_en_0, // @[:@12297.4]
  input         io_rPort_5_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_5_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@12297.4]
  input         io_rPort_4_en_0, // @[:@12297.4]
  input         io_rPort_4_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_4_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@12297.4]
  input         io_rPort_3_en_0, // @[:@12297.4]
  input         io_rPort_3_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_3_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@12297.4]
  input         io_rPort_2_en_0, // @[:@12297.4]
  input         io_rPort_2_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_2_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@12297.4]
  input         io_rPort_1_en_0, // @[:@12297.4]
  input         io_rPort_1_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_1_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@12297.4]
  input         io_rPort_0_en_0, // @[:@12297.4]
  input         io_rPort_0_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_0_output_0, // @[:@12297.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@12297.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@12297.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@12297.4]
  input  [31:0] io_wPort_1_data_0, // @[:@12297.4]
  input         io_wPort_1_en_0, // @[:@12297.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@12297.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12297.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@12297.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12297.4]
  input         io_wPort_0_en_0 // @[:@12297.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@14965.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@12644.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@12645.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@12646.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@12647.4]
  wire [41:0] _T_450; // @[Cat.scala 30:58:@12649.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@12656.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@12657.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@12658.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@12659.4]
  wire [41:0] _T_461; // @[Cat.scala 30:58:@12661.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@12669.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@12670.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@12671.4]
  wire [41:0] _T_472; // @[Cat.scala 30:58:@12673.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@12681.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@12682.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@12683.4]
  wire [41:0] _T_483; // @[Cat.scala 30:58:@12685.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@12692.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@12694.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@12695.4]
  wire [41:0] _T_494; // @[Cat.scala 30:58:@12697.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@12704.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@12706.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@12707.4]
  wire [41:0] _T_505; // @[Cat.scala 30:58:@12709.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@12718.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@12719.4]
  wire [41:0] _T_516; // @[Cat.scala 30:58:@12721.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@12730.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@12731.4]
  wire [41:0] _T_527; // @[Cat.scala 30:58:@12733.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@12740.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@12742.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@12743.4]
  wire [41:0] _T_538; // @[Cat.scala 30:58:@12745.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@12752.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@12754.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@12755.4]
  wire [41:0] _T_549; // @[Cat.scala 30:58:@12757.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@12766.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@12767.4]
  wire [41:0] _T_560; // @[Cat.scala 30:58:@12769.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@12778.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@12779.4]
  wire [41:0] _T_571; // @[Cat.scala 30:58:@12781.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@12788.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@12790.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@12791.4]
  wire [41:0] _T_582; // @[Cat.scala 30:58:@12793.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@12800.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@12802.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@12803.4]
  wire [41:0] _T_593; // @[Cat.scala 30:58:@12805.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@12814.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@12815.4]
  wire [41:0] _T_604; // @[Cat.scala 30:58:@12817.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@12826.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@12827.4]
  wire [41:0] _T_615; // @[Cat.scala 30:58:@12829.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@12836.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@12837.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@12838.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@12840.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@12841.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@12842.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@12844.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@12845.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@12846.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@12848.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@12849.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@12850.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@12852.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@12853.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@12854.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@12856.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@12857.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@12858.4]
  wire  _T_655; // @[MemPrimitives.scala 126:35:@12869.4]
  wire  _T_656; // @[MemPrimitives.scala 126:35:@12870.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@12871.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@12872.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@12873.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@12874.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@12876.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@12878.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@12880.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@12882.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@12884.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@12886.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@12887.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@12888.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@12889.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@12890.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@12891.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@12898.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@12899.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@12900.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@12902.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@12903.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@12904.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@12906.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@12907.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@12908.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@12910.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@12911.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@12912.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@12914.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@12915.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@12916.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@12918.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@12919.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@12920.4]
  wire  _T_717; // @[MemPrimitives.scala 126:35:@12931.4]
  wire  _T_718; // @[MemPrimitives.scala 126:35:@12932.4]
  wire  _T_719; // @[MemPrimitives.scala 126:35:@12933.4]
  wire  _T_720; // @[MemPrimitives.scala 126:35:@12934.4]
  wire  _T_721; // @[MemPrimitives.scala 126:35:@12935.4]
  wire  _T_722; // @[MemPrimitives.scala 126:35:@12936.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@12938.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@12940.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@12942.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@12944.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@12946.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@12948.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@12949.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@12950.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@12951.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@12952.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@12953.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@12961.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@12962.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@12965.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@12966.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@12969.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@12970.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@12973.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@12974.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@12977.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@12978.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@12981.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@12982.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@12993.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@12994.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@12995.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@12996.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@12997.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@12998.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@13000.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@13002.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@13004.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@13006.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@13008.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@13010.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@13011.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@13012.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@13013.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@13014.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@13015.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@13023.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@13024.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@13027.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@13028.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@13031.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@13032.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@13035.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@13036.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@13039.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@13040.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@13043.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@13044.4]
  wire  _T_841; // @[MemPrimitives.scala 126:35:@13055.4]
  wire  _T_842; // @[MemPrimitives.scala 126:35:@13056.4]
  wire  _T_843; // @[MemPrimitives.scala 126:35:@13057.4]
  wire  _T_844; // @[MemPrimitives.scala 126:35:@13058.4]
  wire  _T_845; // @[MemPrimitives.scala 126:35:@13059.4]
  wire  _T_846; // @[MemPrimitives.scala 126:35:@13060.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@13062.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@13064.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@13066.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@13068.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@13070.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@13072.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@13073.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@13074.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@13075.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@13076.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@13077.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@13084.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@13086.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@13088.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@13090.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@13092.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@13094.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@13096.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@13098.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@13100.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@13102.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@13104.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@13106.4]
  wire  _T_903; // @[MemPrimitives.scala 126:35:@13117.4]
  wire  _T_904; // @[MemPrimitives.scala 126:35:@13118.4]
  wire  _T_905; // @[MemPrimitives.scala 126:35:@13119.4]
  wire  _T_906; // @[MemPrimitives.scala 126:35:@13120.4]
  wire  _T_907; // @[MemPrimitives.scala 126:35:@13121.4]
  wire  _T_908; // @[MemPrimitives.scala 126:35:@13122.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@13124.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@13126.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@13128.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@13130.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@13132.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@13134.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@13135.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@13136.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@13137.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@13138.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@13139.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@13146.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@13148.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@13150.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@13152.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@13154.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@13156.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@13158.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@13160.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@13162.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@13164.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@13166.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@13168.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13179.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13180.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13181.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13182.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13183.4]
  wire  _T_970; // @[MemPrimitives.scala 126:35:@13184.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@13186.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@13188.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@13190.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@13192.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@13194.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@13196.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@13197.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@13198.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@13199.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@13200.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@13201.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@13210.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@13214.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@13218.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@13222.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@13226.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@13230.4]
  wire  _T_1027; // @[MemPrimitives.scala 126:35:@13241.4]
  wire  _T_1028; // @[MemPrimitives.scala 126:35:@13242.4]
  wire  _T_1029; // @[MemPrimitives.scala 126:35:@13243.4]
  wire  _T_1030; // @[MemPrimitives.scala 126:35:@13244.4]
  wire  _T_1031; // @[MemPrimitives.scala 126:35:@13245.4]
  wire  _T_1032; // @[MemPrimitives.scala 126:35:@13246.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@13248.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@13250.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@13252.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@13254.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@13256.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@13258.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@13259.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@13260.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@13261.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@13262.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@13263.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@13272.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@13276.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@13280.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@13284.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_1089; // @[MemPrimitives.scala 126:35:@13303.4]
  wire  _T_1090; // @[MemPrimitives.scala 126:35:@13304.4]
  wire  _T_1091; // @[MemPrimitives.scala 126:35:@13305.4]
  wire  _T_1092; // @[MemPrimitives.scala 126:35:@13306.4]
  wire  _T_1093; // @[MemPrimitives.scala 126:35:@13307.4]
  wire  _T_1094; // @[MemPrimitives.scala 126:35:@13308.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@13310.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@13312.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@13314.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@13316.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@13318.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@13320.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@13321.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@13322.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@13323.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@13324.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@13325.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@13332.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13334.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@13336.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13338.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@13340.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13342.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@13344.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13346.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@13348.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13350.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@13352.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@13354.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13365.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13366.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13367.4]
  wire  _T_1154; // @[MemPrimitives.scala 126:35:@13368.4]
  wire  _T_1155; // @[MemPrimitives.scala 126:35:@13369.4]
  wire  _T_1156; // @[MemPrimitives.scala 126:35:@13370.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@13372.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@13374.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@13376.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@13378.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@13380.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@13382.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@13383.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@13384.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@13385.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@13386.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@13387.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@13394.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@13396.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@13398.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13400.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@13402.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13404.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@13406.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13408.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@13410.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13412.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@13414.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13416.4]
  wire  _T_1213; // @[MemPrimitives.scala 126:35:@13427.4]
  wire  _T_1214; // @[MemPrimitives.scala 126:35:@13428.4]
  wire  _T_1215; // @[MemPrimitives.scala 126:35:@13429.4]
  wire  _T_1216; // @[MemPrimitives.scala 126:35:@13430.4]
  wire  _T_1217; // @[MemPrimitives.scala 126:35:@13431.4]
  wire  _T_1218; // @[MemPrimitives.scala 126:35:@13432.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@13434.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@13436.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@13438.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@13440.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@13442.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@13444.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@13445.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@13446.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@13447.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@13448.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@13449.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@13458.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@13462.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@13466.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@13470.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_1275; // @[MemPrimitives.scala 126:35:@13489.4]
  wire  _T_1276; // @[MemPrimitives.scala 126:35:@13490.4]
  wire  _T_1277; // @[MemPrimitives.scala 126:35:@13491.4]
  wire  _T_1278; // @[MemPrimitives.scala 126:35:@13492.4]
  wire  _T_1279; // @[MemPrimitives.scala 126:35:@13493.4]
  wire  _T_1280; // @[MemPrimitives.scala 126:35:@13494.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@13496.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@13498.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@13500.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@13502.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@13504.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@13506.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@13507.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@13508.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@13509.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@13510.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@13511.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@13520.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@13524.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@13528.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@13532.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@13536.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@13540.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13551.4]
  wire  _T_1338; // @[MemPrimitives.scala 126:35:@13552.4]
  wire  _T_1339; // @[MemPrimitives.scala 126:35:@13553.4]
  wire  _T_1340; // @[MemPrimitives.scala 126:35:@13554.4]
  wire  _T_1341; // @[MemPrimitives.scala 126:35:@13555.4]
  wire  _T_1342; // @[MemPrimitives.scala 126:35:@13556.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@13558.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@13560.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@13562.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@13564.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@13566.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@13568.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@13569.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@13570.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@13571.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@13572.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@13573.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@13580.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@13582.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@13584.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@13586.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@13588.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@13590.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@13592.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@13594.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@13596.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@13598.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@13600.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@13602.4]
  wire  _T_1399; // @[MemPrimitives.scala 126:35:@13613.4]
  wire  _T_1400; // @[MemPrimitives.scala 126:35:@13614.4]
  wire  _T_1401; // @[MemPrimitives.scala 126:35:@13615.4]
  wire  _T_1402; // @[MemPrimitives.scala 126:35:@13616.4]
  wire  _T_1403; // @[MemPrimitives.scala 126:35:@13617.4]
  wire  _T_1404; // @[MemPrimitives.scala 126:35:@13618.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@13620.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@13622.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@13624.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@13626.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@13628.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@13630.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@13631.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@13632.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@13633.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@13634.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@13635.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@13642.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@13644.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@13646.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@13648.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@13650.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@13652.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@13654.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@13656.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@13658.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@13662.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1461; // @[MemPrimitives.scala 126:35:@13675.4]
  wire  _T_1462; // @[MemPrimitives.scala 126:35:@13676.4]
  wire  _T_1463; // @[MemPrimitives.scala 126:35:@13677.4]
  wire  _T_1464; // @[MemPrimitives.scala 126:35:@13678.4]
  wire  _T_1465; // @[MemPrimitives.scala 126:35:@13679.4]
  wire  _T_1466; // @[MemPrimitives.scala 126:35:@13680.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@13682.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@13684.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@13686.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@13688.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@13690.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@13692.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@13693.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@13694.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@13695.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@13696.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@13697.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@13706.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@13710.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@13714.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@13718.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@13722.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@13726.4]
  wire  _T_1523; // @[MemPrimitives.scala 126:35:@13737.4]
  wire  _T_1524; // @[MemPrimitives.scala 126:35:@13738.4]
  wire  _T_1525; // @[MemPrimitives.scala 126:35:@13739.4]
  wire  _T_1526; // @[MemPrimitives.scala 126:35:@13740.4]
  wire  _T_1527; // @[MemPrimitives.scala 126:35:@13741.4]
  wire  _T_1528; // @[MemPrimitives.scala 126:35:@13742.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@13744.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@13746.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@13748.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@13750.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@13752.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@13754.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@13755.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@13756.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@13757.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@13758.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@13759.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@13768.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@13772.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@13776.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@13780.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@13784.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@13788.4]
  wire  _T_1585; // @[MemPrimitives.scala 126:35:@13799.4]
  wire  _T_1586; // @[MemPrimitives.scala 126:35:@13800.4]
  wire  _T_1587; // @[MemPrimitives.scala 126:35:@13801.4]
  wire  _T_1588; // @[MemPrimitives.scala 126:35:@13802.4]
  wire  _T_1589; // @[MemPrimitives.scala 126:35:@13803.4]
  wire  _T_1590; // @[MemPrimitives.scala 126:35:@13804.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@13806.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@13808.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@13810.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@13812.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@13814.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@13816.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@13817.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@13818.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@13819.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@13820.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@13821.4]
  wire  _T_1671; // @[package.scala 96:25:@13906.4 package.scala 96:25:@13907.4]
  wire [31:0] _T_1675; // @[Mux.scala 31:69:@13916.4]
  wire  _T_1668; // @[package.scala 96:25:@13898.4 package.scala 96:25:@13899.4]
  wire [31:0] _T_1676; // @[Mux.scala 31:69:@13917.4]
  wire  _T_1665; // @[package.scala 96:25:@13890.4 package.scala 96:25:@13891.4]
  wire [31:0] _T_1677; // @[Mux.scala 31:69:@13918.4]
  wire  _T_1662; // @[package.scala 96:25:@13882.4 package.scala 96:25:@13883.4]
  wire [31:0] _T_1678; // @[Mux.scala 31:69:@13919.4]
  wire  _T_1659; // @[package.scala 96:25:@13874.4 package.scala 96:25:@13875.4]
  wire [31:0] _T_1679; // @[Mux.scala 31:69:@13920.4]
  wire  _T_1656; // @[package.scala 96:25:@13866.4 package.scala 96:25:@13867.4]
  wire [31:0] _T_1680; // @[Mux.scala 31:69:@13921.4]
  wire  _T_1653; // @[package.scala 96:25:@13858.4 package.scala 96:25:@13859.4]
  wire  _T_1742; // @[package.scala 96:25:@14002.4 package.scala 96:25:@14003.4]
  wire [31:0] _T_1746; // @[Mux.scala 31:69:@14012.4]
  wire  _T_1739; // @[package.scala 96:25:@13994.4 package.scala 96:25:@13995.4]
  wire [31:0] _T_1747; // @[Mux.scala 31:69:@14013.4]
  wire  _T_1736; // @[package.scala 96:25:@13986.4 package.scala 96:25:@13987.4]
  wire [31:0] _T_1748; // @[Mux.scala 31:69:@14014.4]
  wire  _T_1733; // @[package.scala 96:25:@13978.4 package.scala 96:25:@13979.4]
  wire [31:0] _T_1749; // @[Mux.scala 31:69:@14015.4]
  wire  _T_1730; // @[package.scala 96:25:@13970.4 package.scala 96:25:@13971.4]
  wire [31:0] _T_1750; // @[Mux.scala 31:69:@14016.4]
  wire  _T_1727; // @[package.scala 96:25:@13962.4 package.scala 96:25:@13963.4]
  wire [31:0] _T_1751; // @[Mux.scala 31:69:@14017.4]
  wire  _T_1724; // @[package.scala 96:25:@13954.4 package.scala 96:25:@13955.4]
  wire  _T_1813; // @[package.scala 96:25:@14098.4 package.scala 96:25:@14099.4]
  wire [31:0] _T_1817; // @[Mux.scala 31:69:@14108.4]
  wire  _T_1810; // @[package.scala 96:25:@14090.4 package.scala 96:25:@14091.4]
  wire [31:0] _T_1818; // @[Mux.scala 31:69:@14109.4]
  wire  _T_1807; // @[package.scala 96:25:@14082.4 package.scala 96:25:@14083.4]
  wire [31:0] _T_1819; // @[Mux.scala 31:69:@14110.4]
  wire  _T_1804; // @[package.scala 96:25:@14074.4 package.scala 96:25:@14075.4]
  wire [31:0] _T_1820; // @[Mux.scala 31:69:@14111.4]
  wire  _T_1801; // @[package.scala 96:25:@14066.4 package.scala 96:25:@14067.4]
  wire [31:0] _T_1821; // @[Mux.scala 31:69:@14112.4]
  wire  _T_1798; // @[package.scala 96:25:@14058.4 package.scala 96:25:@14059.4]
  wire [31:0] _T_1822; // @[Mux.scala 31:69:@14113.4]
  wire  _T_1795; // @[package.scala 96:25:@14050.4 package.scala 96:25:@14051.4]
  wire  _T_1884; // @[package.scala 96:25:@14194.4 package.scala 96:25:@14195.4]
  wire [31:0] _T_1888; // @[Mux.scala 31:69:@14204.4]
  wire  _T_1881; // @[package.scala 96:25:@14186.4 package.scala 96:25:@14187.4]
  wire [31:0] _T_1889; // @[Mux.scala 31:69:@14205.4]
  wire  _T_1878; // @[package.scala 96:25:@14178.4 package.scala 96:25:@14179.4]
  wire [31:0] _T_1890; // @[Mux.scala 31:69:@14206.4]
  wire  _T_1875; // @[package.scala 96:25:@14170.4 package.scala 96:25:@14171.4]
  wire [31:0] _T_1891; // @[Mux.scala 31:69:@14207.4]
  wire  _T_1872; // @[package.scala 96:25:@14162.4 package.scala 96:25:@14163.4]
  wire [31:0] _T_1892; // @[Mux.scala 31:69:@14208.4]
  wire  _T_1869; // @[package.scala 96:25:@14154.4 package.scala 96:25:@14155.4]
  wire [31:0] _T_1893; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1866; // @[package.scala 96:25:@14146.4 package.scala 96:25:@14147.4]
  wire  _T_1955; // @[package.scala 96:25:@14290.4 package.scala 96:25:@14291.4]
  wire [31:0] _T_1959; // @[Mux.scala 31:69:@14300.4]
  wire  _T_1952; // @[package.scala 96:25:@14282.4 package.scala 96:25:@14283.4]
  wire [31:0] _T_1960; // @[Mux.scala 31:69:@14301.4]
  wire  _T_1949; // @[package.scala 96:25:@14274.4 package.scala 96:25:@14275.4]
  wire [31:0] _T_1961; // @[Mux.scala 31:69:@14302.4]
  wire  _T_1946; // @[package.scala 96:25:@14266.4 package.scala 96:25:@14267.4]
  wire [31:0] _T_1962; // @[Mux.scala 31:69:@14303.4]
  wire  _T_1943; // @[package.scala 96:25:@14258.4 package.scala 96:25:@14259.4]
  wire [31:0] _T_1963; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1940; // @[package.scala 96:25:@14250.4 package.scala 96:25:@14251.4]
  wire [31:0] _T_1964; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1937; // @[package.scala 96:25:@14242.4 package.scala 96:25:@14243.4]
  wire  _T_2026; // @[package.scala 96:25:@14386.4 package.scala 96:25:@14387.4]
  wire [31:0] _T_2030; // @[Mux.scala 31:69:@14396.4]
  wire  _T_2023; // @[package.scala 96:25:@14378.4 package.scala 96:25:@14379.4]
  wire [31:0] _T_2031; // @[Mux.scala 31:69:@14397.4]
  wire  _T_2020; // @[package.scala 96:25:@14370.4 package.scala 96:25:@14371.4]
  wire [31:0] _T_2032; // @[Mux.scala 31:69:@14398.4]
  wire  _T_2017; // @[package.scala 96:25:@14362.4 package.scala 96:25:@14363.4]
  wire [31:0] _T_2033; // @[Mux.scala 31:69:@14399.4]
  wire  _T_2014; // @[package.scala 96:25:@14354.4 package.scala 96:25:@14355.4]
  wire [31:0] _T_2034; // @[Mux.scala 31:69:@14400.4]
  wire  _T_2011; // @[package.scala 96:25:@14346.4 package.scala 96:25:@14347.4]
  wire [31:0] _T_2035; // @[Mux.scala 31:69:@14401.4]
  wire  _T_2008; // @[package.scala 96:25:@14338.4 package.scala 96:25:@14339.4]
  wire  _T_2097; // @[package.scala 96:25:@14482.4 package.scala 96:25:@14483.4]
  wire [31:0] _T_2101; // @[Mux.scala 31:69:@14492.4]
  wire  _T_2094; // @[package.scala 96:25:@14474.4 package.scala 96:25:@14475.4]
  wire [31:0] _T_2102; // @[Mux.scala 31:69:@14493.4]
  wire  _T_2091; // @[package.scala 96:25:@14466.4 package.scala 96:25:@14467.4]
  wire [31:0] _T_2103; // @[Mux.scala 31:69:@14494.4]
  wire  _T_2088; // @[package.scala 96:25:@14458.4 package.scala 96:25:@14459.4]
  wire [31:0] _T_2104; // @[Mux.scala 31:69:@14495.4]
  wire  _T_2085; // @[package.scala 96:25:@14450.4 package.scala 96:25:@14451.4]
  wire [31:0] _T_2105; // @[Mux.scala 31:69:@14496.4]
  wire  _T_2082; // @[package.scala 96:25:@14442.4 package.scala 96:25:@14443.4]
  wire [31:0] _T_2106; // @[Mux.scala 31:69:@14497.4]
  wire  _T_2079; // @[package.scala 96:25:@14434.4 package.scala 96:25:@14435.4]
  wire  _T_2168; // @[package.scala 96:25:@14578.4 package.scala 96:25:@14579.4]
  wire [31:0] _T_2172; // @[Mux.scala 31:69:@14588.4]
  wire  _T_2165; // @[package.scala 96:25:@14570.4 package.scala 96:25:@14571.4]
  wire [31:0] _T_2173; // @[Mux.scala 31:69:@14589.4]
  wire  _T_2162; // @[package.scala 96:25:@14562.4 package.scala 96:25:@14563.4]
  wire [31:0] _T_2174; // @[Mux.scala 31:69:@14590.4]
  wire  _T_2159; // @[package.scala 96:25:@14554.4 package.scala 96:25:@14555.4]
  wire [31:0] _T_2175; // @[Mux.scala 31:69:@14591.4]
  wire  _T_2156; // @[package.scala 96:25:@14546.4 package.scala 96:25:@14547.4]
  wire [31:0] _T_2176; // @[Mux.scala 31:69:@14592.4]
  wire  _T_2153; // @[package.scala 96:25:@14538.4 package.scala 96:25:@14539.4]
  wire [31:0] _T_2177; // @[Mux.scala 31:69:@14593.4]
  wire  _T_2150; // @[package.scala 96:25:@14530.4 package.scala 96:25:@14531.4]
  wire  _T_2239; // @[package.scala 96:25:@14674.4 package.scala 96:25:@14675.4]
  wire [31:0] _T_2243; // @[Mux.scala 31:69:@14684.4]
  wire  _T_2236; // @[package.scala 96:25:@14666.4 package.scala 96:25:@14667.4]
  wire [31:0] _T_2244; // @[Mux.scala 31:69:@14685.4]
  wire  _T_2233; // @[package.scala 96:25:@14658.4 package.scala 96:25:@14659.4]
  wire [31:0] _T_2245; // @[Mux.scala 31:69:@14686.4]
  wire  _T_2230; // @[package.scala 96:25:@14650.4 package.scala 96:25:@14651.4]
  wire [31:0] _T_2246; // @[Mux.scala 31:69:@14687.4]
  wire  _T_2227; // @[package.scala 96:25:@14642.4 package.scala 96:25:@14643.4]
  wire [31:0] _T_2247; // @[Mux.scala 31:69:@14688.4]
  wire  _T_2224; // @[package.scala 96:25:@14634.4 package.scala 96:25:@14635.4]
  wire [31:0] _T_2248; // @[Mux.scala 31:69:@14689.4]
  wire  _T_2221; // @[package.scala 96:25:@14626.4 package.scala 96:25:@14627.4]
  wire  _T_2310; // @[package.scala 96:25:@14770.4 package.scala 96:25:@14771.4]
  wire [31:0] _T_2314; // @[Mux.scala 31:69:@14780.4]
  wire  _T_2307; // @[package.scala 96:25:@14762.4 package.scala 96:25:@14763.4]
  wire [31:0] _T_2315; // @[Mux.scala 31:69:@14781.4]
  wire  _T_2304; // @[package.scala 96:25:@14754.4 package.scala 96:25:@14755.4]
  wire [31:0] _T_2316; // @[Mux.scala 31:69:@14782.4]
  wire  _T_2301; // @[package.scala 96:25:@14746.4 package.scala 96:25:@14747.4]
  wire [31:0] _T_2317; // @[Mux.scala 31:69:@14783.4]
  wire  _T_2298; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  wire [31:0] _T_2318; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2295; // @[package.scala 96:25:@14730.4 package.scala 96:25:@14731.4]
  wire [31:0] _T_2319; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2292; // @[package.scala 96:25:@14722.4 package.scala 96:25:@14723.4]
  wire  _T_2381; // @[package.scala 96:25:@14866.4 package.scala 96:25:@14867.4]
  wire [31:0] _T_2385; // @[Mux.scala 31:69:@14876.4]
  wire  _T_2378; // @[package.scala 96:25:@14858.4 package.scala 96:25:@14859.4]
  wire [31:0] _T_2386; // @[Mux.scala 31:69:@14877.4]
  wire  _T_2375; // @[package.scala 96:25:@14850.4 package.scala 96:25:@14851.4]
  wire [31:0] _T_2387; // @[Mux.scala 31:69:@14878.4]
  wire  _T_2372; // @[package.scala 96:25:@14842.4 package.scala 96:25:@14843.4]
  wire [31:0] _T_2388; // @[Mux.scala 31:69:@14879.4]
  wire  _T_2369; // @[package.scala 96:25:@14834.4 package.scala 96:25:@14835.4]
  wire [31:0] _T_2389; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2366; // @[package.scala 96:25:@14826.4 package.scala 96:25:@14827.4]
  wire [31:0] _T_2390; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2363; // @[package.scala 96:25:@14818.4 package.scala 96:25:@14819.4]
  wire  _T_2452; // @[package.scala 96:25:@14962.4 package.scala 96:25:@14963.4]
  wire [31:0] _T_2456; // @[Mux.scala 31:69:@14972.4]
  wire  _T_2449; // @[package.scala 96:25:@14954.4 package.scala 96:25:@14955.4]
  wire [31:0] _T_2457; // @[Mux.scala 31:69:@14973.4]
  wire  _T_2446; // @[package.scala 96:25:@14946.4 package.scala 96:25:@14947.4]
  wire [31:0] _T_2458; // @[Mux.scala 31:69:@14974.4]
  wire  _T_2443; // @[package.scala 96:25:@14938.4 package.scala 96:25:@14939.4]
  wire [31:0] _T_2459; // @[Mux.scala 31:69:@14975.4]
  wire  _T_2440; // @[package.scala 96:25:@14930.4 package.scala 96:25:@14931.4]
  wire [31:0] _T_2460; // @[Mux.scala 31:69:@14976.4]
  wire  _T_2437; // @[package.scala 96:25:@14922.4 package.scala 96:25:@14923.4]
  wire [31:0] _T_2461; // @[Mux.scala 31:69:@14977.4]
  wire  _T_2434; // @[package.scala 96:25:@14914.4 package.scala 96:25:@14915.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12388.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12404.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12420.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12436.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12452.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12468.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12484.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12500.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12516.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12532.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12548.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12564.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@12580.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@12596.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@12612.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@12628.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@12860.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@12922.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@12984.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13046.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13108.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13170.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13232.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13294.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13356.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13418.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13480.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13542.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@13604.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@13666.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@13728.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@13790.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@13853.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@13861.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@13869.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@13877.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@13885.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@13893.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@13901.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@13909.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@13949.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@13957.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@13965.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@13973.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@13981.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@13989.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@13997.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14005.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14045.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14053.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14061.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14069.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14077.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14085.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14093.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14101.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14141.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14149.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14157.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14165.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14173.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14181.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14189.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14197.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14237.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14245.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14253.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14261.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14269.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14277.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14285.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14293.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14333.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14341.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14349.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14357.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14365.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14373.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14381.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14389.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14429.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14437.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14445.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14453.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14461.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14469.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14477.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14485.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14525.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14533.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14541.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14549.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14557.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14565.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14573.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14581.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14621.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14629.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14637.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14645.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14653.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14661.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14669.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14677.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14717.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14725.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14733.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@14741.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@14749.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@14757.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@14765.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@14773.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@14813.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@14821.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@14829.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@14837.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@14845.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@14853.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@14861.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@14869.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@14909.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@14917.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@14925.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@14933.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@14941.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@14949.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@14957.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@14965.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12644.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@12645.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@12646.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@12647.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12649.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12656.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@12657.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@12658.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@12659.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12661.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@12669.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@12670.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@12671.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12673.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@12681.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@12682.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@12683.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12685.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12692.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@12694.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@12695.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12697.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12704.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@12706.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@12707.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12709.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@12718.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@12719.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12721.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@12730.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@12731.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12733.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12740.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@12742.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@12743.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12745.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12752.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@12754.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@12755.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12757.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@12766.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@12767.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12769.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@12778.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@12779.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12781.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12788.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@12790.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@12791.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12793.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12800.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@12802.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@12803.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12805.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@12814.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@12815.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12817.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@12826.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@12827.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12829.4]
  assign _T_620 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12836.4]
  assign _T_622 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12837.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@12838.4]
  assign _T_626 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12840.4]
  assign _T_628 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12841.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@12842.4]
  assign _T_632 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12844.4]
  assign _T_634 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12845.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@12846.4]
  assign _T_638 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12848.4]
  assign _T_640 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12849.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@12850.4]
  assign _T_644 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12852.4]
  assign _T_646 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12853.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@12854.4]
  assign _T_650 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12856.4]
  assign _T_652 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12857.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@12858.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@12869.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@12870.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@12871.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@12872.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@12873.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@12874.4]
  assign _T_662 = {_T_655,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12876.4]
  assign _T_664 = {_T_656,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12878.4]
  assign _T_666 = {_T_657,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12880.4]
  assign _T_668 = {_T_658,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12882.4]
  assign _T_670 = {_T_659,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12884.4]
  assign _T_672 = {_T_660,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@12886.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@12887.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@12888.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@12889.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@12890.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@12891.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12898.4]
  assign _T_684 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12899.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@12900.4]
  assign _T_688 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12902.4]
  assign _T_690 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12903.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@12904.4]
  assign _T_694 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12906.4]
  assign _T_696 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12907.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@12908.4]
  assign _T_700 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12910.4]
  assign _T_702 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12911.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@12912.4]
  assign _T_706 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12914.4]
  assign _T_708 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12915.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@12916.4]
  assign _T_712 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12918.4]
  assign _T_714 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12919.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@12920.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@12931.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@12932.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@12933.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@12934.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@12935.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@12936.4]
  assign _T_724 = {_T_717,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12938.4]
  assign _T_726 = {_T_718,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12940.4]
  assign _T_728 = {_T_719,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12942.4]
  assign _T_730 = {_T_720,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12944.4]
  assign _T_732 = {_T_721,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@12946.4]
  assign _T_734 = {_T_722,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@12948.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@12949.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@12950.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@12951.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@12952.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@12953.4]
  assign _T_746 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12961.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@12962.4]
  assign _T_752 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12965.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@12966.4]
  assign _T_758 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12969.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@12970.4]
  assign _T_764 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12973.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@12974.4]
  assign _T_770 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12977.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@12978.4]
  assign _T_776 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12981.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@12982.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@12993.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@12994.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@12995.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@12996.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@12997.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@12998.4]
  assign _T_786 = {_T_779,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13000.4]
  assign _T_788 = {_T_780,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13002.4]
  assign _T_790 = {_T_781,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13004.4]
  assign _T_792 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13006.4]
  assign _T_794 = {_T_783,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13008.4]
  assign _T_796 = {_T_784,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13010.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@13011.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@13012.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@13013.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@13014.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@13015.4]
  assign _T_808 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13023.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@13024.4]
  assign _T_814 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13027.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@13028.4]
  assign _T_820 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13031.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@13032.4]
  assign _T_826 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13035.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@13036.4]
  assign _T_832 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13039.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@13040.4]
  assign _T_838 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13043.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@13044.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13055.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13056.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13057.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13058.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13059.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13060.4]
  assign _T_848 = {_T_841,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13062.4]
  assign _T_850 = {_T_842,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13064.4]
  assign _T_852 = {_T_843,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13066.4]
  assign _T_854 = {_T_844,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13068.4]
  assign _T_856 = {_T_845,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13070.4]
  assign _T_858 = {_T_846,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13072.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@13073.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@13074.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@13075.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@13076.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@13077.4]
  assign _T_868 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13084.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@13086.4]
  assign _T_874 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13088.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@13090.4]
  assign _T_880 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13092.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@13094.4]
  assign _T_886 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13096.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@13098.4]
  assign _T_892 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13100.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@13102.4]
  assign _T_898 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13104.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@13106.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13117.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13118.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13119.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13120.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13121.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13122.4]
  assign _T_910 = {_T_903,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13124.4]
  assign _T_912 = {_T_904,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13126.4]
  assign _T_914 = {_T_905,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13128.4]
  assign _T_916 = {_T_906,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13130.4]
  assign _T_918 = {_T_907,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13132.4]
  assign _T_920 = {_T_908,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13134.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@13135.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@13136.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@13137.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@13138.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@13139.4]
  assign _T_930 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13146.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@13148.4]
  assign _T_936 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13150.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@13152.4]
  assign _T_942 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13154.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@13156.4]
  assign _T_948 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13158.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@13160.4]
  assign _T_954 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13162.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@13164.4]
  assign _T_960 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13166.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@13168.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13179.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13180.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13181.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13182.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13183.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13184.4]
  assign _T_972 = {_T_965,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13186.4]
  assign _T_974 = {_T_966,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13188.4]
  assign _T_976 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13190.4]
  assign _T_978 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13192.4]
  assign _T_980 = {_T_969,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13194.4]
  assign _T_982 = {_T_970,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13196.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@13197.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@13198.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@13199.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@13200.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@13201.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@13210.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@13214.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@13218.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@13222.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@13226.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@13230.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13241.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13242.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13243.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13244.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13245.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13246.4]
  assign _T_1034 = {_T_1027,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13248.4]
  assign _T_1036 = {_T_1028,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13250.4]
  assign _T_1038 = {_T_1029,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13252.4]
  assign _T_1040 = {_T_1030,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13254.4]
  assign _T_1042 = {_T_1031,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13256.4]
  assign _T_1044 = {_T_1032,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13258.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@13259.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@13260.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@13261.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@13262.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@13263.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@13272.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@13276.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@13280.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@13284.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13303.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13304.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13305.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13306.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13307.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13308.4]
  assign _T_1096 = {_T_1089,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13310.4]
  assign _T_1098 = {_T_1090,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13312.4]
  assign _T_1100 = {_T_1091,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13314.4]
  assign _T_1102 = {_T_1092,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13316.4]
  assign _T_1104 = {_T_1093,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13318.4]
  assign _T_1106 = {_T_1094,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13320.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@13321.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@13322.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@13323.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@13324.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@13325.4]
  assign _T_1116 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13332.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@13334.4]
  assign _T_1122 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13336.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@13338.4]
  assign _T_1128 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13340.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@13342.4]
  assign _T_1134 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13344.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@13346.4]
  assign _T_1140 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13348.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@13350.4]
  assign _T_1146 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13352.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@13354.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13365.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13366.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13367.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13368.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13369.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13370.4]
  assign _T_1158 = {_T_1151,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13372.4]
  assign _T_1160 = {_T_1152,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13374.4]
  assign _T_1162 = {_T_1153,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13376.4]
  assign _T_1164 = {_T_1154,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13378.4]
  assign _T_1166 = {_T_1155,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13380.4]
  assign _T_1168 = {_T_1156,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13382.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@13383.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@13384.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@13385.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@13386.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@13387.4]
  assign _T_1178 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13394.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@13396.4]
  assign _T_1184 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13398.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@13400.4]
  assign _T_1190 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13402.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@13404.4]
  assign _T_1196 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13406.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@13408.4]
  assign _T_1202 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13410.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@13412.4]
  assign _T_1208 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13414.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@13416.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13427.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13428.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13429.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13430.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13431.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13432.4]
  assign _T_1220 = {_T_1213,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13434.4]
  assign _T_1222 = {_T_1214,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13436.4]
  assign _T_1224 = {_T_1215,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13438.4]
  assign _T_1226 = {_T_1216,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13440.4]
  assign _T_1228 = {_T_1217,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13442.4]
  assign _T_1230 = {_T_1218,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13444.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@13445.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@13446.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@13447.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@13448.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@13449.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@13458.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@13462.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@13466.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@13470.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13489.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13490.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13491.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13492.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13493.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13494.4]
  assign _T_1282 = {_T_1275,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13496.4]
  assign _T_1284 = {_T_1276,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13498.4]
  assign _T_1286 = {_T_1277,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13500.4]
  assign _T_1288 = {_T_1278,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13502.4]
  assign _T_1290 = {_T_1279,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13504.4]
  assign _T_1292 = {_T_1280,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13506.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@13507.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@13508.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@13509.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@13510.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@13511.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@13520.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@13524.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@13528.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@13532.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@13536.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@13540.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13551.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13552.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13553.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13554.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13555.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13556.4]
  assign _T_1344 = {_T_1337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13558.4]
  assign _T_1346 = {_T_1338,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13560.4]
  assign _T_1348 = {_T_1339,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13562.4]
  assign _T_1350 = {_T_1340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13564.4]
  assign _T_1352 = {_T_1341,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13566.4]
  assign _T_1354 = {_T_1342,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13568.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@13569.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@13570.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@13571.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@13572.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@13573.4]
  assign _T_1364 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13580.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@13582.4]
  assign _T_1370 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13584.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@13586.4]
  assign _T_1376 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13588.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@13590.4]
  assign _T_1382 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13592.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@13594.4]
  assign _T_1388 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13596.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@13598.4]
  assign _T_1394 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13600.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@13602.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@13613.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@13614.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@13615.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@13616.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@13617.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@13618.4]
  assign _T_1406 = {_T_1399,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13620.4]
  assign _T_1408 = {_T_1400,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13622.4]
  assign _T_1410 = {_T_1401,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13624.4]
  assign _T_1412 = {_T_1402,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13626.4]
  assign _T_1414 = {_T_1403,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13628.4]
  assign _T_1416 = {_T_1404,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13630.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@13631.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@13632.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@13633.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@13634.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@13635.4]
  assign _T_1426 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13642.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@13644.4]
  assign _T_1432 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13646.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@13648.4]
  assign _T_1438 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13650.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@13652.4]
  assign _T_1444 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13654.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@13656.4]
  assign _T_1450 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13658.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1456 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13662.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@13675.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@13676.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@13677.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@13678.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@13679.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@13680.4]
  assign _T_1468 = {_T_1461,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13682.4]
  assign _T_1470 = {_T_1462,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13684.4]
  assign _T_1472 = {_T_1463,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13686.4]
  assign _T_1474 = {_T_1464,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13688.4]
  assign _T_1476 = {_T_1465,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13690.4]
  assign _T_1478 = {_T_1466,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13692.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@13693.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@13694.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@13695.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@13696.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@13697.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@13706.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@13710.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@13714.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@13718.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@13722.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@13726.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@13737.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@13738.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@13739.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@13740.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@13741.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@13742.4]
  assign _T_1530 = {_T_1523,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13744.4]
  assign _T_1532 = {_T_1524,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13746.4]
  assign _T_1534 = {_T_1525,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13748.4]
  assign _T_1536 = {_T_1526,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13750.4]
  assign _T_1538 = {_T_1527,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13752.4]
  assign _T_1540 = {_T_1528,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13754.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@13755.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@13756.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@13757.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@13758.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@13759.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@13768.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@13772.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@13776.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@13780.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@13784.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@13788.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@13799.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@13800.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@13801.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@13802.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@13803.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@13804.4]
  assign _T_1592 = {_T_1585,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13806.4]
  assign _T_1594 = {_T_1586,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13808.4]
  assign _T_1596 = {_T_1587,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13810.4]
  assign _T_1598 = {_T_1588,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13812.4]
  assign _T_1600 = {_T_1589,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13814.4]
  assign _T_1602 = {_T_1590,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13816.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@13817.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@13818.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@13819.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@13820.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@13821.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@13906.4 package.scala 96:25:@13907.4]
  assign _T_1675 = _T_1671 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@13916.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@13898.4 package.scala 96:25:@13899.4]
  assign _T_1676 = _T_1668 ? Mem1D_10_io_output : _T_1675; // @[Mux.scala 31:69:@13917.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@13890.4 package.scala 96:25:@13891.4]
  assign _T_1677 = _T_1665 ? Mem1D_8_io_output : _T_1676; // @[Mux.scala 31:69:@13918.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@13882.4 package.scala 96:25:@13883.4]
  assign _T_1678 = _T_1662 ? Mem1D_6_io_output : _T_1677; // @[Mux.scala 31:69:@13919.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@13874.4 package.scala 96:25:@13875.4]
  assign _T_1679 = _T_1659 ? Mem1D_4_io_output : _T_1678; // @[Mux.scala 31:69:@13920.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@13866.4 package.scala 96:25:@13867.4]
  assign _T_1680 = _T_1656 ? Mem1D_2_io_output : _T_1679; // @[Mux.scala 31:69:@13921.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@13858.4 package.scala 96:25:@13859.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14002.4 package.scala 96:25:@14003.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14012.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@13994.4 package.scala 96:25:@13995.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@14013.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@13986.4 package.scala 96:25:@13987.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@14014.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@13978.4 package.scala 96:25:@13979.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@14015.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@13970.4 package.scala 96:25:@13971.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@14016.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@13962.4 package.scala 96:25:@13963.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@14017.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@13954.4 package.scala 96:25:@13955.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14098.4 package.scala 96:25:@14099.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14108.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14090.4 package.scala 96:25:@14091.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@14109.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14082.4 package.scala 96:25:@14083.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@14110.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14074.4 package.scala 96:25:@14075.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@14111.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14066.4 package.scala 96:25:@14067.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@14112.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14058.4 package.scala 96:25:@14059.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@14113.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14050.4 package.scala 96:25:@14051.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14194.4 package.scala 96:25:@14195.4]
  assign _T_1888 = _T_1884 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14204.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14186.4 package.scala 96:25:@14187.4]
  assign _T_1889 = _T_1881 ? Mem1D_10_io_output : _T_1888; // @[Mux.scala 31:69:@14205.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14178.4 package.scala 96:25:@14179.4]
  assign _T_1890 = _T_1878 ? Mem1D_8_io_output : _T_1889; // @[Mux.scala 31:69:@14206.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14170.4 package.scala 96:25:@14171.4]
  assign _T_1891 = _T_1875 ? Mem1D_6_io_output : _T_1890; // @[Mux.scala 31:69:@14207.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14162.4 package.scala 96:25:@14163.4]
  assign _T_1892 = _T_1872 ? Mem1D_4_io_output : _T_1891; // @[Mux.scala 31:69:@14208.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14154.4 package.scala 96:25:@14155.4]
  assign _T_1893 = _T_1869 ? Mem1D_2_io_output : _T_1892; // @[Mux.scala 31:69:@14209.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14146.4 package.scala 96:25:@14147.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14290.4 package.scala 96:25:@14291.4]
  assign _T_1959 = _T_1955 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14300.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14282.4 package.scala 96:25:@14283.4]
  assign _T_1960 = _T_1952 ? Mem1D_11_io_output : _T_1959; // @[Mux.scala 31:69:@14301.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14274.4 package.scala 96:25:@14275.4]
  assign _T_1961 = _T_1949 ? Mem1D_9_io_output : _T_1960; // @[Mux.scala 31:69:@14302.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@14266.4 package.scala 96:25:@14267.4]
  assign _T_1962 = _T_1946 ? Mem1D_7_io_output : _T_1961; // @[Mux.scala 31:69:@14303.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14258.4 package.scala 96:25:@14259.4]
  assign _T_1963 = _T_1943 ? Mem1D_5_io_output : _T_1962; // @[Mux.scala 31:69:@14304.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14250.4 package.scala 96:25:@14251.4]
  assign _T_1964 = _T_1940 ? Mem1D_3_io_output : _T_1963; // @[Mux.scala 31:69:@14305.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14242.4 package.scala 96:25:@14243.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14386.4 package.scala 96:25:@14387.4]
  assign _T_2030 = _T_2026 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14396.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14378.4 package.scala 96:25:@14379.4]
  assign _T_2031 = _T_2023 ? Mem1D_10_io_output : _T_2030; // @[Mux.scala 31:69:@14397.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14370.4 package.scala 96:25:@14371.4]
  assign _T_2032 = _T_2020 ? Mem1D_8_io_output : _T_2031; // @[Mux.scala 31:69:@14398.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14362.4 package.scala 96:25:@14363.4]
  assign _T_2033 = _T_2017 ? Mem1D_6_io_output : _T_2032; // @[Mux.scala 31:69:@14399.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14354.4 package.scala 96:25:@14355.4]
  assign _T_2034 = _T_2014 ? Mem1D_4_io_output : _T_2033; // @[Mux.scala 31:69:@14400.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14346.4 package.scala 96:25:@14347.4]
  assign _T_2035 = _T_2011 ? Mem1D_2_io_output : _T_2034; // @[Mux.scala 31:69:@14401.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14338.4 package.scala 96:25:@14339.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14482.4 package.scala 96:25:@14483.4]
  assign _T_2101 = _T_2097 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14492.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14474.4 package.scala 96:25:@14475.4]
  assign _T_2102 = _T_2094 ? Mem1D_11_io_output : _T_2101; // @[Mux.scala 31:69:@14493.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14466.4 package.scala 96:25:@14467.4]
  assign _T_2103 = _T_2091 ? Mem1D_9_io_output : _T_2102; // @[Mux.scala 31:69:@14494.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14458.4 package.scala 96:25:@14459.4]
  assign _T_2104 = _T_2088 ? Mem1D_7_io_output : _T_2103; // @[Mux.scala 31:69:@14495.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14450.4 package.scala 96:25:@14451.4]
  assign _T_2105 = _T_2085 ? Mem1D_5_io_output : _T_2104; // @[Mux.scala 31:69:@14496.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14442.4 package.scala 96:25:@14443.4]
  assign _T_2106 = _T_2082 ? Mem1D_3_io_output : _T_2105; // @[Mux.scala 31:69:@14497.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14434.4 package.scala 96:25:@14435.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14578.4 package.scala 96:25:@14579.4]
  assign _T_2172 = _T_2168 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14588.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14570.4 package.scala 96:25:@14571.4]
  assign _T_2173 = _T_2165 ? Mem1D_11_io_output : _T_2172; // @[Mux.scala 31:69:@14589.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14562.4 package.scala 96:25:@14563.4]
  assign _T_2174 = _T_2162 ? Mem1D_9_io_output : _T_2173; // @[Mux.scala 31:69:@14590.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14554.4 package.scala 96:25:@14555.4]
  assign _T_2175 = _T_2159 ? Mem1D_7_io_output : _T_2174; // @[Mux.scala 31:69:@14591.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14546.4 package.scala 96:25:@14547.4]
  assign _T_2176 = _T_2156 ? Mem1D_5_io_output : _T_2175; // @[Mux.scala 31:69:@14592.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14538.4 package.scala 96:25:@14539.4]
  assign _T_2177 = _T_2153 ? Mem1D_3_io_output : _T_2176; // @[Mux.scala 31:69:@14593.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14530.4 package.scala 96:25:@14531.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14674.4 package.scala 96:25:@14675.4]
  assign _T_2243 = _T_2239 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14684.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14666.4 package.scala 96:25:@14667.4]
  assign _T_2244 = _T_2236 ? Mem1D_10_io_output : _T_2243; // @[Mux.scala 31:69:@14685.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14658.4 package.scala 96:25:@14659.4]
  assign _T_2245 = _T_2233 ? Mem1D_8_io_output : _T_2244; // @[Mux.scala 31:69:@14686.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14650.4 package.scala 96:25:@14651.4]
  assign _T_2246 = _T_2230 ? Mem1D_6_io_output : _T_2245; // @[Mux.scala 31:69:@14687.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14642.4 package.scala 96:25:@14643.4]
  assign _T_2247 = _T_2227 ? Mem1D_4_io_output : _T_2246; // @[Mux.scala 31:69:@14688.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14634.4 package.scala 96:25:@14635.4]
  assign _T_2248 = _T_2224 ? Mem1D_2_io_output : _T_2247; // @[Mux.scala 31:69:@14689.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14626.4 package.scala 96:25:@14627.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@14770.4 package.scala 96:25:@14771.4]
  assign _T_2314 = _T_2310 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14780.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@14762.4 package.scala 96:25:@14763.4]
  assign _T_2315 = _T_2307 ? Mem1D_11_io_output : _T_2314; // @[Mux.scala 31:69:@14781.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@14754.4 package.scala 96:25:@14755.4]
  assign _T_2316 = _T_2304 ? Mem1D_9_io_output : _T_2315; // @[Mux.scala 31:69:@14782.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@14746.4 package.scala 96:25:@14747.4]
  assign _T_2317 = _T_2301 ? Mem1D_7_io_output : _T_2316; // @[Mux.scala 31:69:@14783.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  assign _T_2318 = _T_2298 ? Mem1D_5_io_output : _T_2317; // @[Mux.scala 31:69:@14784.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14730.4 package.scala 96:25:@14731.4]
  assign _T_2319 = _T_2295 ? Mem1D_3_io_output : _T_2318; // @[Mux.scala 31:69:@14785.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14722.4 package.scala 96:25:@14723.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@14866.4 package.scala 96:25:@14867.4]
  assign _T_2385 = _T_2381 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14876.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@14858.4 package.scala 96:25:@14859.4]
  assign _T_2386 = _T_2378 ? Mem1D_10_io_output : _T_2385; // @[Mux.scala 31:69:@14877.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@14850.4 package.scala 96:25:@14851.4]
  assign _T_2387 = _T_2375 ? Mem1D_8_io_output : _T_2386; // @[Mux.scala 31:69:@14878.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@14842.4 package.scala 96:25:@14843.4]
  assign _T_2388 = _T_2372 ? Mem1D_6_io_output : _T_2387; // @[Mux.scala 31:69:@14879.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@14834.4 package.scala 96:25:@14835.4]
  assign _T_2389 = _T_2369 ? Mem1D_4_io_output : _T_2388; // @[Mux.scala 31:69:@14880.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@14826.4 package.scala 96:25:@14827.4]
  assign _T_2390 = _T_2366 ? Mem1D_2_io_output : _T_2389; // @[Mux.scala 31:69:@14881.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@14818.4 package.scala 96:25:@14819.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@14962.4 package.scala 96:25:@14963.4]
  assign _T_2456 = _T_2452 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14972.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@14954.4 package.scala 96:25:@14955.4]
  assign _T_2457 = _T_2449 ? Mem1D_11_io_output : _T_2456; // @[Mux.scala 31:69:@14973.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@14946.4 package.scala 96:25:@14947.4]
  assign _T_2458 = _T_2446 ? Mem1D_9_io_output : _T_2457; // @[Mux.scala 31:69:@14974.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@14938.4 package.scala 96:25:@14939.4]
  assign _T_2459 = _T_2443 ? Mem1D_7_io_output : _T_2458; // @[Mux.scala 31:69:@14975.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@14930.4 package.scala 96:25:@14931.4]
  assign _T_2460 = _T_2440 ? Mem1D_5_io_output : _T_2459; // @[Mux.scala 31:69:@14976.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@14922.4 package.scala 96:25:@14923.4]
  assign _T_2461 = _T_2437 ? Mem1D_3_io_output : _T_2460; // @[Mux.scala 31:69:@14977.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@14914.4 package.scala 96:25:@14915.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_1_io_output : _T_2461; // @[MemPrimitives.scala 152:13:@14979.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_io_output : _T_2390; // @[MemPrimitives.scala 152:13:@14883.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_1_io_output : _T_2319; // @[MemPrimitives.scala 152:13:@14787.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_io_output : _T_2248; // @[MemPrimitives.scala 152:13:@14691.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_1_io_output : _T_2177; // @[MemPrimitives.scala 152:13:@14595.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_1_io_output : _T_2106; // @[MemPrimitives.scala 152:13:@14499.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_io_output : _T_2035; // @[MemPrimitives.scala 152:13:@14403.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_1_io_output : _T_1964; // @[MemPrimitives.scala 152:13:@14307.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_io_output : _T_1893; // @[MemPrimitives.scala 152:13:@14211.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 152:13:@14115.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 152:13:@14019.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_io_output : _T_1680; // @[MemPrimitives.scala 152:13:@13923.4]
  assign Mem1D_clock = clock; // @[:@12389.4]
  assign Mem1D_reset = reset; // @[:@12390.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 131:28:@12895.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 132:32:@12896.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@12653.4]
  assign Mem1D_io_w_data_0 = _T_450[40:9]; // @[MemPrimitives.scala 95:29:@12654.4]
  assign Mem1D_io_w_en_0 = _T_450[41]; // @[MemPrimitives.scala 96:27:@12655.4]
  assign Mem1D_1_clock = clock; // @[:@12405.4]
  assign Mem1D_1_reset = reset; // @[:@12406.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 131:28:@12957.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 132:32:@12958.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@12665.4]
  assign Mem1D_1_io_w_data_0 = _T_461[40:9]; // @[MemPrimitives.scala 95:29:@12666.4]
  assign Mem1D_1_io_w_en_0 = _T_461[41]; // @[MemPrimitives.scala 96:27:@12667.4]
  assign Mem1D_2_clock = clock; // @[:@12421.4]
  assign Mem1D_2_reset = reset; // @[:@12422.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 131:28:@13019.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 132:32:@13020.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@12677.4]
  assign Mem1D_2_io_w_data_0 = _T_472[40:9]; // @[MemPrimitives.scala 95:29:@12678.4]
  assign Mem1D_2_io_w_en_0 = _T_472[41]; // @[MemPrimitives.scala 96:27:@12679.4]
  assign Mem1D_3_clock = clock; // @[:@12437.4]
  assign Mem1D_3_reset = reset; // @[:@12438.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 131:28:@13081.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 132:32:@13082.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@12689.4]
  assign Mem1D_3_io_w_data_0 = _T_483[40:9]; // @[MemPrimitives.scala 95:29:@12690.4]
  assign Mem1D_3_io_w_en_0 = _T_483[41]; // @[MemPrimitives.scala 96:27:@12691.4]
  assign Mem1D_4_clock = clock; // @[:@12453.4]
  assign Mem1D_4_reset = reset; // @[:@12454.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 131:28:@13143.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 132:32:@13144.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@12701.4]
  assign Mem1D_4_io_w_data_0 = _T_494[40:9]; // @[MemPrimitives.scala 95:29:@12702.4]
  assign Mem1D_4_io_w_en_0 = _T_494[41]; // @[MemPrimitives.scala 96:27:@12703.4]
  assign Mem1D_5_clock = clock; // @[:@12469.4]
  assign Mem1D_5_reset = reset; // @[:@12470.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 131:28:@13205.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 132:32:@13206.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@12713.4]
  assign Mem1D_5_io_w_data_0 = _T_505[40:9]; // @[MemPrimitives.scala 95:29:@12714.4]
  assign Mem1D_5_io_w_en_0 = _T_505[41]; // @[MemPrimitives.scala 96:27:@12715.4]
  assign Mem1D_6_clock = clock; // @[:@12485.4]
  assign Mem1D_6_reset = reset; // @[:@12486.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 131:28:@13267.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 132:32:@13268.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@12725.4]
  assign Mem1D_6_io_w_data_0 = _T_516[40:9]; // @[MemPrimitives.scala 95:29:@12726.4]
  assign Mem1D_6_io_w_en_0 = _T_516[41]; // @[MemPrimitives.scala 96:27:@12727.4]
  assign Mem1D_7_clock = clock; // @[:@12501.4]
  assign Mem1D_7_reset = reset; // @[:@12502.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 131:28:@13329.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 132:32:@13330.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@12737.4]
  assign Mem1D_7_io_w_data_0 = _T_527[40:9]; // @[MemPrimitives.scala 95:29:@12738.4]
  assign Mem1D_7_io_w_en_0 = _T_527[41]; // @[MemPrimitives.scala 96:27:@12739.4]
  assign Mem1D_8_clock = clock; // @[:@12517.4]
  assign Mem1D_8_reset = reset; // @[:@12518.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 131:28:@13391.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 132:32:@13392.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@12749.4]
  assign Mem1D_8_io_w_data_0 = _T_538[40:9]; // @[MemPrimitives.scala 95:29:@12750.4]
  assign Mem1D_8_io_w_en_0 = _T_538[41]; // @[MemPrimitives.scala 96:27:@12751.4]
  assign Mem1D_9_clock = clock; // @[:@12533.4]
  assign Mem1D_9_reset = reset; // @[:@12534.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 131:28:@13453.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 132:32:@13454.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@12761.4]
  assign Mem1D_9_io_w_data_0 = _T_549[40:9]; // @[MemPrimitives.scala 95:29:@12762.4]
  assign Mem1D_9_io_w_en_0 = _T_549[41]; // @[MemPrimitives.scala 96:27:@12763.4]
  assign Mem1D_10_clock = clock; // @[:@12549.4]
  assign Mem1D_10_reset = reset; // @[:@12550.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 131:28:@13515.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 132:32:@13516.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@12773.4]
  assign Mem1D_10_io_w_data_0 = _T_560[40:9]; // @[MemPrimitives.scala 95:29:@12774.4]
  assign Mem1D_10_io_w_en_0 = _T_560[41]; // @[MemPrimitives.scala 96:27:@12775.4]
  assign Mem1D_11_clock = clock; // @[:@12565.4]
  assign Mem1D_11_reset = reset; // @[:@12566.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@13577.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@13578.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@12785.4]
  assign Mem1D_11_io_w_data_0 = _T_571[40:9]; // @[MemPrimitives.scala 95:29:@12786.4]
  assign Mem1D_11_io_w_en_0 = _T_571[41]; // @[MemPrimitives.scala 96:27:@12787.4]
  assign Mem1D_12_clock = clock; // @[:@12581.4]
  assign Mem1D_12_reset = reset; // @[:@12582.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 131:28:@13639.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 132:32:@13640.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@12797.4]
  assign Mem1D_12_io_w_data_0 = _T_582[40:9]; // @[MemPrimitives.scala 95:29:@12798.4]
  assign Mem1D_12_io_w_en_0 = _T_582[41]; // @[MemPrimitives.scala 96:27:@12799.4]
  assign Mem1D_13_clock = clock; // @[:@12597.4]
  assign Mem1D_13_reset = reset; // @[:@12598.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 131:28:@13701.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 132:32:@13702.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@12809.4]
  assign Mem1D_13_io_w_data_0 = _T_593[40:9]; // @[MemPrimitives.scala 95:29:@12810.4]
  assign Mem1D_13_io_w_en_0 = _T_593[41]; // @[MemPrimitives.scala 96:27:@12811.4]
  assign Mem1D_14_clock = clock; // @[:@12613.4]
  assign Mem1D_14_reset = reset; // @[:@12614.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 131:28:@13763.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 132:32:@13764.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@12821.4]
  assign Mem1D_14_io_w_data_0 = _T_604[40:9]; // @[MemPrimitives.scala 95:29:@12822.4]
  assign Mem1D_14_io_w_en_0 = _T_604[41]; // @[MemPrimitives.scala 96:27:@12823.4]
  assign Mem1D_15_clock = clock; // @[:@12629.4]
  assign Mem1D_15_reset = reset; // @[:@12630.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 131:28:@13825.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 132:32:@13826.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@12833.4]
  assign Mem1D_15_io_w_data_0 = _T_615[40:9]; // @[MemPrimitives.scala 95:29:@12834.4]
  assign Mem1D_15_io_w_en_0 = _T_615[41]; // @[MemPrimitives.scala 96:27:@12835.4]
  assign StickySelects_clock = clock; // @[:@12861.4]
  assign StickySelects_reset = reset; // @[:@12862.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_623; // @[MemPrimitives.scala 125:64:@12863.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_629; // @[MemPrimitives.scala 125:64:@12864.4]
  assign StickySelects_io_ins_2 = io_rPort_3_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@12865.4]
  assign StickySelects_io_ins_3 = io_rPort_5_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@12866.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@12867.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@12868.4]
  assign StickySelects_1_clock = clock; // @[:@12923.4]
  assign StickySelects_1_reset = reset; // @[:@12924.4]
  assign StickySelects_1_io_ins_0 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@12925.4]
  assign StickySelects_1_io_ins_1 = io_rPort_4_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@12926.4]
  assign StickySelects_1_io_ins_2 = io_rPort_6_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@12927.4]
  assign StickySelects_1_io_ins_3 = io_rPort_7_en_0 & _T_703; // @[MemPrimitives.scala 125:64:@12928.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_709; // @[MemPrimitives.scala 125:64:@12929.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_715; // @[MemPrimitives.scala 125:64:@12930.4]
  assign StickySelects_2_clock = clock; // @[:@12985.4]
  assign StickySelects_2_reset = reset; // @[:@12986.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_747; // @[MemPrimitives.scala 125:64:@12987.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_753; // @[MemPrimitives.scala 125:64:@12988.4]
  assign StickySelects_2_io_ins_2 = io_rPort_3_en_0 & _T_759; // @[MemPrimitives.scala 125:64:@12989.4]
  assign StickySelects_2_io_ins_3 = io_rPort_5_en_0 & _T_765; // @[MemPrimitives.scala 125:64:@12990.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_771; // @[MemPrimitives.scala 125:64:@12991.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_777; // @[MemPrimitives.scala 125:64:@12992.4]
  assign StickySelects_3_clock = clock; // @[:@13047.4]
  assign StickySelects_3_reset = reset; // @[:@13048.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_809; // @[MemPrimitives.scala 125:64:@13049.4]
  assign StickySelects_3_io_ins_1 = io_rPort_4_en_0 & _T_815; // @[MemPrimitives.scala 125:64:@13050.4]
  assign StickySelects_3_io_ins_2 = io_rPort_6_en_0 & _T_821; // @[MemPrimitives.scala 125:64:@13051.4]
  assign StickySelects_3_io_ins_3 = io_rPort_7_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@13052.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@13053.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_839; // @[MemPrimitives.scala 125:64:@13054.4]
  assign StickySelects_4_clock = clock; // @[:@13109.4]
  assign StickySelects_4_reset = reset; // @[:@13110.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_871; // @[MemPrimitives.scala 125:64:@13111.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_877; // @[MemPrimitives.scala 125:64:@13112.4]
  assign StickySelects_4_io_ins_2 = io_rPort_3_en_0 & _T_883; // @[MemPrimitives.scala 125:64:@13113.4]
  assign StickySelects_4_io_ins_3 = io_rPort_5_en_0 & _T_889; // @[MemPrimitives.scala 125:64:@13114.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_895; // @[MemPrimitives.scala 125:64:@13115.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_901; // @[MemPrimitives.scala 125:64:@13116.4]
  assign StickySelects_5_clock = clock; // @[:@13171.4]
  assign StickySelects_5_reset = reset; // @[:@13172.4]
  assign StickySelects_5_io_ins_0 = io_rPort_1_en_0 & _T_933; // @[MemPrimitives.scala 125:64:@13173.4]
  assign StickySelects_5_io_ins_1 = io_rPort_4_en_0 & _T_939; // @[MemPrimitives.scala 125:64:@13174.4]
  assign StickySelects_5_io_ins_2 = io_rPort_6_en_0 & _T_945; // @[MemPrimitives.scala 125:64:@13175.4]
  assign StickySelects_5_io_ins_3 = io_rPort_7_en_0 & _T_951; // @[MemPrimitives.scala 125:64:@13176.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_957; // @[MemPrimitives.scala 125:64:@13177.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_963; // @[MemPrimitives.scala 125:64:@13178.4]
  assign StickySelects_6_clock = clock; // @[:@13233.4]
  assign StickySelects_6_reset = reset; // @[:@13234.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_995; // @[MemPrimitives.scala 125:64:@13235.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_1001; // @[MemPrimitives.scala 125:64:@13236.4]
  assign StickySelects_6_io_ins_2 = io_rPort_3_en_0 & _T_1007; // @[MemPrimitives.scala 125:64:@13237.4]
  assign StickySelects_6_io_ins_3 = io_rPort_5_en_0 & _T_1013; // @[MemPrimitives.scala 125:64:@13238.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1019; // @[MemPrimitives.scala 125:64:@13239.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1025; // @[MemPrimitives.scala 125:64:@13240.4]
  assign StickySelects_7_clock = clock; // @[:@13295.4]
  assign StickySelects_7_reset = reset; // @[:@13296.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1057; // @[MemPrimitives.scala 125:64:@13297.4]
  assign StickySelects_7_io_ins_1 = io_rPort_4_en_0 & _T_1063; // @[MemPrimitives.scala 125:64:@13298.4]
  assign StickySelects_7_io_ins_2 = io_rPort_6_en_0 & _T_1069; // @[MemPrimitives.scala 125:64:@13299.4]
  assign StickySelects_7_io_ins_3 = io_rPort_7_en_0 & _T_1075; // @[MemPrimitives.scala 125:64:@13300.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1081; // @[MemPrimitives.scala 125:64:@13301.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1087; // @[MemPrimitives.scala 125:64:@13302.4]
  assign StickySelects_8_clock = clock; // @[:@13357.4]
  assign StickySelects_8_reset = reset; // @[:@13358.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13359.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13360.4]
  assign StickySelects_8_io_ins_2 = io_rPort_3_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13361.4]
  assign StickySelects_8_io_ins_3 = io_rPort_5_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13362.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13363.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1149; // @[MemPrimitives.scala 125:64:@13364.4]
  assign StickySelects_9_clock = clock; // @[:@13419.4]
  assign StickySelects_9_reset = reset; // @[:@13420.4]
  assign StickySelects_9_io_ins_0 = io_rPort_1_en_0 & _T_1181; // @[MemPrimitives.scala 125:64:@13421.4]
  assign StickySelects_9_io_ins_1 = io_rPort_4_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13422.4]
  assign StickySelects_9_io_ins_2 = io_rPort_6_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13423.4]
  assign StickySelects_9_io_ins_3 = io_rPort_7_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13424.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13425.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13426.4]
  assign StickySelects_10_clock = clock; // @[:@13481.4]
  assign StickySelects_10_reset = reset; // @[:@13482.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1243; // @[MemPrimitives.scala 125:64:@13483.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_1249; // @[MemPrimitives.scala 125:64:@13484.4]
  assign StickySelects_10_io_ins_2 = io_rPort_3_en_0 & _T_1255; // @[MemPrimitives.scala 125:64:@13485.4]
  assign StickySelects_10_io_ins_3 = io_rPort_5_en_0 & _T_1261; // @[MemPrimitives.scala 125:64:@13486.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_1267; // @[MemPrimitives.scala 125:64:@13487.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_1273; // @[MemPrimitives.scala 125:64:@13488.4]
  assign StickySelects_11_clock = clock; // @[:@13543.4]
  assign StickySelects_11_reset = reset; // @[:@13544.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@13545.4]
  assign StickySelects_11_io_ins_1 = io_rPort_4_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@13546.4]
  assign StickySelects_11_io_ins_2 = io_rPort_6_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@13547.4]
  assign StickySelects_11_io_ins_3 = io_rPort_7_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@13548.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_1329; // @[MemPrimitives.scala 125:64:@13549.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1335; // @[MemPrimitives.scala 125:64:@13550.4]
  assign StickySelects_12_clock = clock; // @[:@13605.4]
  assign StickySelects_12_reset = reset; // @[:@13606.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@13607.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@13608.4]
  assign StickySelects_12_io_ins_2 = io_rPort_3_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@13609.4]
  assign StickySelects_12_io_ins_3 = io_rPort_5_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@13610.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@13611.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@13612.4]
  assign StickySelects_13_clock = clock; // @[:@13667.4]
  assign StickySelects_13_reset = reset; // @[:@13668.4]
  assign StickySelects_13_io_ins_0 = io_rPort_1_en_0 & _T_1429; // @[MemPrimitives.scala 125:64:@13669.4]
  assign StickySelects_13_io_ins_1 = io_rPort_4_en_0 & _T_1435; // @[MemPrimitives.scala 125:64:@13670.4]
  assign StickySelects_13_io_ins_2 = io_rPort_6_en_0 & _T_1441; // @[MemPrimitives.scala 125:64:@13671.4]
  assign StickySelects_13_io_ins_3 = io_rPort_7_en_0 & _T_1447; // @[MemPrimitives.scala 125:64:@13672.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_1453; // @[MemPrimitives.scala 125:64:@13673.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@13674.4]
  assign StickySelects_14_clock = clock; // @[:@13729.4]
  assign StickySelects_14_reset = reset; // @[:@13730.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_1491; // @[MemPrimitives.scala 125:64:@13731.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_1497; // @[MemPrimitives.scala 125:64:@13732.4]
  assign StickySelects_14_io_ins_2 = io_rPort_3_en_0 & _T_1503; // @[MemPrimitives.scala 125:64:@13733.4]
  assign StickySelects_14_io_ins_3 = io_rPort_5_en_0 & _T_1509; // @[MemPrimitives.scala 125:64:@13734.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_1515; // @[MemPrimitives.scala 125:64:@13735.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_1521; // @[MemPrimitives.scala 125:64:@13736.4]
  assign StickySelects_15_clock = clock; // @[:@13791.4]
  assign StickySelects_15_reset = reset; // @[:@13792.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1553; // @[MemPrimitives.scala 125:64:@13793.4]
  assign StickySelects_15_io_ins_1 = io_rPort_4_en_0 & _T_1559; // @[MemPrimitives.scala 125:64:@13794.4]
  assign StickySelects_15_io_ins_2 = io_rPort_6_en_0 & _T_1565; // @[MemPrimitives.scala 125:64:@13795.4]
  assign StickySelects_15_io_ins_3 = io_rPort_7_en_0 & _T_1571; // @[MemPrimitives.scala 125:64:@13796.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_1577; // @[MemPrimitives.scala 125:64:@13797.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1583; // @[MemPrimitives.scala 125:64:@13798.4]
  assign RetimeWrapper_clock = clock; // @[:@13854.4]
  assign RetimeWrapper_reset = reset; // @[:@13855.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13857.4]
  assign RetimeWrapper_io_in = _T_623 & io_rPort_0_en_0; // @[package.scala 94:16:@13856.4]
  assign RetimeWrapper_1_clock = clock; // @[:@13862.4]
  assign RetimeWrapper_1_reset = reset; // @[:@13863.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13865.4]
  assign RetimeWrapper_1_io_in = _T_747 & io_rPort_0_en_0; // @[package.scala 94:16:@13864.4]
  assign RetimeWrapper_2_clock = clock; // @[:@13870.4]
  assign RetimeWrapper_2_reset = reset; // @[:@13871.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13873.4]
  assign RetimeWrapper_2_io_in = _T_871 & io_rPort_0_en_0; // @[package.scala 94:16:@13872.4]
  assign RetimeWrapper_3_clock = clock; // @[:@13878.4]
  assign RetimeWrapper_3_reset = reset; // @[:@13879.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13881.4]
  assign RetimeWrapper_3_io_in = _T_995 & io_rPort_0_en_0; // @[package.scala 94:16:@13880.4]
  assign RetimeWrapper_4_clock = clock; // @[:@13886.4]
  assign RetimeWrapper_4_reset = reset; // @[:@13887.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13889.4]
  assign RetimeWrapper_4_io_in = _T_1119 & io_rPort_0_en_0; // @[package.scala 94:16:@13888.4]
  assign RetimeWrapper_5_clock = clock; // @[:@13894.4]
  assign RetimeWrapper_5_reset = reset; // @[:@13895.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13897.4]
  assign RetimeWrapper_5_io_in = _T_1243 & io_rPort_0_en_0; // @[package.scala 94:16:@13896.4]
  assign RetimeWrapper_6_clock = clock; // @[:@13902.4]
  assign RetimeWrapper_6_reset = reset; // @[:@13903.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13905.4]
  assign RetimeWrapper_6_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@13904.4]
  assign RetimeWrapper_7_clock = clock; // @[:@13910.4]
  assign RetimeWrapper_7_reset = reset; // @[:@13911.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13913.4]
  assign RetimeWrapper_7_io_in = _T_1491 & io_rPort_0_en_0; // @[package.scala 94:16:@13912.4]
  assign RetimeWrapper_8_clock = clock; // @[:@13950.4]
  assign RetimeWrapper_8_reset = reset; // @[:@13951.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13953.4]
  assign RetimeWrapper_8_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@13952.4]
  assign RetimeWrapper_9_clock = clock; // @[:@13958.4]
  assign RetimeWrapper_9_reset = reset; // @[:@13959.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13961.4]
  assign RetimeWrapper_9_io_in = _T_809 & io_rPort_1_en_0; // @[package.scala 94:16:@13960.4]
  assign RetimeWrapper_10_clock = clock; // @[:@13966.4]
  assign RetimeWrapper_10_reset = reset; // @[:@13967.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13969.4]
  assign RetimeWrapper_10_io_in = _T_933 & io_rPort_1_en_0; // @[package.scala 94:16:@13968.4]
  assign RetimeWrapper_11_clock = clock; // @[:@13974.4]
  assign RetimeWrapper_11_reset = reset; // @[:@13975.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13977.4]
  assign RetimeWrapper_11_io_in = _T_1057 & io_rPort_1_en_0; // @[package.scala 94:16:@13976.4]
  assign RetimeWrapper_12_clock = clock; // @[:@13982.4]
  assign RetimeWrapper_12_reset = reset; // @[:@13983.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13985.4]
  assign RetimeWrapper_12_io_in = _T_1181 & io_rPort_1_en_0; // @[package.scala 94:16:@13984.4]
  assign RetimeWrapper_13_clock = clock; // @[:@13990.4]
  assign RetimeWrapper_13_reset = reset; // @[:@13991.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13993.4]
  assign RetimeWrapper_13_io_in = _T_1305 & io_rPort_1_en_0; // @[package.scala 94:16:@13992.4]
  assign RetimeWrapper_14_clock = clock; // @[:@13998.4]
  assign RetimeWrapper_14_reset = reset; // @[:@13999.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14001.4]
  assign RetimeWrapper_14_io_in = _T_1429 & io_rPort_1_en_0; // @[package.scala 94:16:@14000.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14006.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14007.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14009.4]
  assign RetimeWrapper_15_io_in = _T_1553 & io_rPort_1_en_0; // @[package.scala 94:16:@14008.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14046.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14047.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14049.4]
  assign RetimeWrapper_16_io_in = _T_629 & io_rPort_2_en_0; // @[package.scala 94:16:@14048.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14054.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14055.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14057.4]
  assign RetimeWrapper_17_io_in = _T_753 & io_rPort_2_en_0; // @[package.scala 94:16:@14056.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14062.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14063.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14065.4]
  assign RetimeWrapper_18_io_in = _T_877 & io_rPort_2_en_0; // @[package.scala 94:16:@14064.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14070.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14071.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14073.4]
  assign RetimeWrapper_19_io_in = _T_1001 & io_rPort_2_en_0; // @[package.scala 94:16:@14072.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14078.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14079.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14081.4]
  assign RetimeWrapper_20_io_in = _T_1125 & io_rPort_2_en_0; // @[package.scala 94:16:@14080.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14086.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14087.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14089.4]
  assign RetimeWrapper_21_io_in = _T_1249 & io_rPort_2_en_0; // @[package.scala 94:16:@14088.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14094.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14095.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14097.4]
  assign RetimeWrapper_22_io_in = _T_1373 & io_rPort_2_en_0; // @[package.scala 94:16:@14096.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14102.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14103.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14105.4]
  assign RetimeWrapper_23_io_in = _T_1497 & io_rPort_2_en_0; // @[package.scala 94:16:@14104.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14142.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14143.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14145.4]
  assign RetimeWrapper_24_io_in = _T_635 & io_rPort_3_en_0; // @[package.scala 94:16:@14144.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14150.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14151.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14153.4]
  assign RetimeWrapper_25_io_in = _T_759 & io_rPort_3_en_0; // @[package.scala 94:16:@14152.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14158.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14159.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14161.4]
  assign RetimeWrapper_26_io_in = _T_883 & io_rPort_3_en_0; // @[package.scala 94:16:@14160.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14166.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14167.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14169.4]
  assign RetimeWrapper_27_io_in = _T_1007 & io_rPort_3_en_0; // @[package.scala 94:16:@14168.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14174.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14175.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14177.4]
  assign RetimeWrapper_28_io_in = _T_1131 & io_rPort_3_en_0; // @[package.scala 94:16:@14176.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14182.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14183.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14185.4]
  assign RetimeWrapper_29_io_in = _T_1255 & io_rPort_3_en_0; // @[package.scala 94:16:@14184.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14190.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14191.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14193.4]
  assign RetimeWrapper_30_io_in = _T_1379 & io_rPort_3_en_0; // @[package.scala 94:16:@14192.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14198.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14199.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14201.4]
  assign RetimeWrapper_31_io_in = _T_1503 & io_rPort_3_en_0; // @[package.scala 94:16:@14200.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14238.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14239.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14241.4]
  assign RetimeWrapper_32_io_in = _T_691 & io_rPort_4_en_0; // @[package.scala 94:16:@14240.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14246.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14247.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14249.4]
  assign RetimeWrapper_33_io_in = _T_815 & io_rPort_4_en_0; // @[package.scala 94:16:@14248.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14254.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14255.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14257.4]
  assign RetimeWrapper_34_io_in = _T_939 & io_rPort_4_en_0; // @[package.scala 94:16:@14256.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14262.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14263.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14265.4]
  assign RetimeWrapper_35_io_in = _T_1063 & io_rPort_4_en_0; // @[package.scala 94:16:@14264.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14270.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14271.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14273.4]
  assign RetimeWrapper_36_io_in = _T_1187 & io_rPort_4_en_0; // @[package.scala 94:16:@14272.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14278.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14279.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14281.4]
  assign RetimeWrapper_37_io_in = _T_1311 & io_rPort_4_en_0; // @[package.scala 94:16:@14280.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14286.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14287.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14289.4]
  assign RetimeWrapper_38_io_in = _T_1435 & io_rPort_4_en_0; // @[package.scala 94:16:@14288.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14294.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14295.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14297.4]
  assign RetimeWrapper_39_io_in = _T_1559 & io_rPort_4_en_0; // @[package.scala 94:16:@14296.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14334.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14335.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14337.4]
  assign RetimeWrapper_40_io_in = _T_641 & io_rPort_5_en_0; // @[package.scala 94:16:@14336.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14342.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14343.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14345.4]
  assign RetimeWrapper_41_io_in = _T_765 & io_rPort_5_en_0; // @[package.scala 94:16:@14344.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14350.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14351.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14353.4]
  assign RetimeWrapper_42_io_in = _T_889 & io_rPort_5_en_0; // @[package.scala 94:16:@14352.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14358.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14359.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14361.4]
  assign RetimeWrapper_43_io_in = _T_1013 & io_rPort_5_en_0; // @[package.scala 94:16:@14360.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14366.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14367.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14369.4]
  assign RetimeWrapper_44_io_in = _T_1137 & io_rPort_5_en_0; // @[package.scala 94:16:@14368.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14374.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14375.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14377.4]
  assign RetimeWrapper_45_io_in = _T_1261 & io_rPort_5_en_0; // @[package.scala 94:16:@14376.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14382.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14383.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14385.4]
  assign RetimeWrapper_46_io_in = _T_1385 & io_rPort_5_en_0; // @[package.scala 94:16:@14384.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14390.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14391.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14393.4]
  assign RetimeWrapper_47_io_in = _T_1509 & io_rPort_5_en_0; // @[package.scala 94:16:@14392.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14430.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14431.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14433.4]
  assign RetimeWrapper_48_io_in = _T_697 & io_rPort_6_en_0; // @[package.scala 94:16:@14432.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14438.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14439.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14441.4]
  assign RetimeWrapper_49_io_in = _T_821 & io_rPort_6_en_0; // @[package.scala 94:16:@14440.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14446.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14447.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14449.4]
  assign RetimeWrapper_50_io_in = _T_945 & io_rPort_6_en_0; // @[package.scala 94:16:@14448.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14454.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14455.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14457.4]
  assign RetimeWrapper_51_io_in = _T_1069 & io_rPort_6_en_0; // @[package.scala 94:16:@14456.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14462.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14463.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14465.4]
  assign RetimeWrapper_52_io_in = _T_1193 & io_rPort_6_en_0; // @[package.scala 94:16:@14464.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14470.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14471.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14473.4]
  assign RetimeWrapper_53_io_in = _T_1317 & io_rPort_6_en_0; // @[package.scala 94:16:@14472.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14478.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14479.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14481.4]
  assign RetimeWrapper_54_io_in = _T_1441 & io_rPort_6_en_0; // @[package.scala 94:16:@14480.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14486.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14487.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14489.4]
  assign RetimeWrapper_55_io_in = _T_1565 & io_rPort_6_en_0; // @[package.scala 94:16:@14488.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14526.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14527.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14529.4]
  assign RetimeWrapper_56_io_in = _T_703 & io_rPort_7_en_0; // @[package.scala 94:16:@14528.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14534.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14535.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14537.4]
  assign RetimeWrapper_57_io_in = _T_827 & io_rPort_7_en_0; // @[package.scala 94:16:@14536.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14542.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14543.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14545.4]
  assign RetimeWrapper_58_io_in = _T_951 & io_rPort_7_en_0; // @[package.scala 94:16:@14544.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14550.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14551.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14553.4]
  assign RetimeWrapper_59_io_in = _T_1075 & io_rPort_7_en_0; // @[package.scala 94:16:@14552.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14558.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14559.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14561.4]
  assign RetimeWrapper_60_io_in = _T_1199 & io_rPort_7_en_0; // @[package.scala 94:16:@14560.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14566.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14567.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14569.4]
  assign RetimeWrapper_61_io_in = _T_1323 & io_rPort_7_en_0; // @[package.scala 94:16:@14568.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14574.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14575.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14577.4]
  assign RetimeWrapper_62_io_in = _T_1447 & io_rPort_7_en_0; // @[package.scala 94:16:@14576.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14582.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14583.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14585.4]
  assign RetimeWrapper_63_io_in = _T_1571 & io_rPort_7_en_0; // @[package.scala 94:16:@14584.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14622.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14623.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14625.4]
  assign RetimeWrapper_64_io_in = _T_647 & io_rPort_8_en_0; // @[package.scala 94:16:@14624.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14630.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14631.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14633.4]
  assign RetimeWrapper_65_io_in = _T_771 & io_rPort_8_en_0; // @[package.scala 94:16:@14632.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14638.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14639.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14641.4]
  assign RetimeWrapper_66_io_in = _T_895 & io_rPort_8_en_0; // @[package.scala 94:16:@14640.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14646.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14647.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14649.4]
  assign RetimeWrapper_67_io_in = _T_1019 & io_rPort_8_en_0; // @[package.scala 94:16:@14648.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14654.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14655.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14657.4]
  assign RetimeWrapper_68_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@14656.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14662.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14663.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14665.4]
  assign RetimeWrapper_69_io_in = _T_1267 & io_rPort_8_en_0; // @[package.scala 94:16:@14664.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14670.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14671.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14673.4]
  assign RetimeWrapper_70_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@14672.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14678.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14679.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14681.4]
  assign RetimeWrapper_71_io_in = _T_1515 & io_rPort_8_en_0; // @[package.scala 94:16:@14680.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14718.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14719.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14721.4]
  assign RetimeWrapper_72_io_in = _T_709 & io_rPort_9_en_0; // @[package.scala 94:16:@14720.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14726.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14727.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14729.4]
  assign RetimeWrapper_73_io_in = _T_833 & io_rPort_9_en_0; // @[package.scala 94:16:@14728.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14734.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14735.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14737.4]
  assign RetimeWrapper_74_io_in = _T_957 & io_rPort_9_en_0; // @[package.scala 94:16:@14736.4]
  assign RetimeWrapper_75_clock = clock; // @[:@14742.4]
  assign RetimeWrapper_75_reset = reset; // @[:@14743.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14745.4]
  assign RetimeWrapper_75_io_in = _T_1081 & io_rPort_9_en_0; // @[package.scala 94:16:@14744.4]
  assign RetimeWrapper_76_clock = clock; // @[:@14750.4]
  assign RetimeWrapper_76_reset = reset; // @[:@14751.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14753.4]
  assign RetimeWrapper_76_io_in = _T_1205 & io_rPort_9_en_0; // @[package.scala 94:16:@14752.4]
  assign RetimeWrapper_77_clock = clock; // @[:@14758.4]
  assign RetimeWrapper_77_reset = reset; // @[:@14759.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14761.4]
  assign RetimeWrapper_77_io_in = _T_1329 & io_rPort_9_en_0; // @[package.scala 94:16:@14760.4]
  assign RetimeWrapper_78_clock = clock; // @[:@14766.4]
  assign RetimeWrapper_78_reset = reset; // @[:@14767.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14769.4]
  assign RetimeWrapper_78_io_in = _T_1453 & io_rPort_9_en_0; // @[package.scala 94:16:@14768.4]
  assign RetimeWrapper_79_clock = clock; // @[:@14774.4]
  assign RetimeWrapper_79_reset = reset; // @[:@14775.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14777.4]
  assign RetimeWrapper_79_io_in = _T_1577 & io_rPort_9_en_0; // @[package.scala 94:16:@14776.4]
  assign RetimeWrapper_80_clock = clock; // @[:@14814.4]
  assign RetimeWrapper_80_reset = reset; // @[:@14815.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14817.4]
  assign RetimeWrapper_80_io_in = _T_653 & io_rPort_10_en_0; // @[package.scala 94:16:@14816.4]
  assign RetimeWrapper_81_clock = clock; // @[:@14822.4]
  assign RetimeWrapper_81_reset = reset; // @[:@14823.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14825.4]
  assign RetimeWrapper_81_io_in = _T_777 & io_rPort_10_en_0; // @[package.scala 94:16:@14824.4]
  assign RetimeWrapper_82_clock = clock; // @[:@14830.4]
  assign RetimeWrapper_82_reset = reset; // @[:@14831.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14833.4]
  assign RetimeWrapper_82_io_in = _T_901 & io_rPort_10_en_0; // @[package.scala 94:16:@14832.4]
  assign RetimeWrapper_83_clock = clock; // @[:@14838.4]
  assign RetimeWrapper_83_reset = reset; // @[:@14839.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14841.4]
  assign RetimeWrapper_83_io_in = _T_1025 & io_rPort_10_en_0; // @[package.scala 94:16:@14840.4]
  assign RetimeWrapper_84_clock = clock; // @[:@14846.4]
  assign RetimeWrapper_84_reset = reset; // @[:@14847.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14849.4]
  assign RetimeWrapper_84_io_in = _T_1149 & io_rPort_10_en_0; // @[package.scala 94:16:@14848.4]
  assign RetimeWrapper_85_clock = clock; // @[:@14854.4]
  assign RetimeWrapper_85_reset = reset; // @[:@14855.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14857.4]
  assign RetimeWrapper_85_io_in = _T_1273 & io_rPort_10_en_0; // @[package.scala 94:16:@14856.4]
  assign RetimeWrapper_86_clock = clock; // @[:@14862.4]
  assign RetimeWrapper_86_reset = reset; // @[:@14863.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14865.4]
  assign RetimeWrapper_86_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@14864.4]
  assign RetimeWrapper_87_clock = clock; // @[:@14870.4]
  assign RetimeWrapper_87_reset = reset; // @[:@14871.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14873.4]
  assign RetimeWrapper_87_io_in = _T_1521 & io_rPort_10_en_0; // @[package.scala 94:16:@14872.4]
  assign RetimeWrapper_88_clock = clock; // @[:@14910.4]
  assign RetimeWrapper_88_reset = reset; // @[:@14911.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14913.4]
  assign RetimeWrapper_88_io_in = _T_715 & io_rPort_11_en_0; // @[package.scala 94:16:@14912.4]
  assign RetimeWrapper_89_clock = clock; // @[:@14918.4]
  assign RetimeWrapper_89_reset = reset; // @[:@14919.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14921.4]
  assign RetimeWrapper_89_io_in = _T_839 & io_rPort_11_en_0; // @[package.scala 94:16:@14920.4]
  assign RetimeWrapper_90_clock = clock; // @[:@14926.4]
  assign RetimeWrapper_90_reset = reset; // @[:@14927.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14929.4]
  assign RetimeWrapper_90_io_in = _T_963 & io_rPort_11_en_0; // @[package.scala 94:16:@14928.4]
  assign RetimeWrapper_91_clock = clock; // @[:@14934.4]
  assign RetimeWrapper_91_reset = reset; // @[:@14935.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14937.4]
  assign RetimeWrapper_91_io_in = _T_1087 & io_rPort_11_en_0; // @[package.scala 94:16:@14936.4]
  assign RetimeWrapper_92_clock = clock; // @[:@14942.4]
  assign RetimeWrapper_92_reset = reset; // @[:@14943.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14945.4]
  assign RetimeWrapper_92_io_in = _T_1211 & io_rPort_11_en_0; // @[package.scala 94:16:@14944.4]
  assign RetimeWrapper_93_clock = clock; // @[:@14950.4]
  assign RetimeWrapper_93_reset = reset; // @[:@14951.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14953.4]
  assign RetimeWrapper_93_io_in = _T_1335 & io_rPort_11_en_0; // @[package.scala 94:16:@14952.4]
  assign RetimeWrapper_94_clock = clock; // @[:@14958.4]
  assign RetimeWrapper_94_reset = reset; // @[:@14959.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14961.4]
  assign RetimeWrapper_94_io_in = _T_1459 & io_rPort_11_en_0; // @[package.scala 94:16:@14960.4]
  assign RetimeWrapper_95_clock = clock; // @[:@14966.4]
  assign RetimeWrapper_95_reset = reset; // @[:@14967.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14969.4]
  assign RetimeWrapper_95_io_in = _T_1583 & io_rPort_11_en_0; // @[package.scala 94:16:@14968.4]
endmodule
module StickySelects_17( // @[:@16693.2]
  input   clock, // @[:@16694.4]
  input   reset, // @[:@16695.4]
  input   io_ins_0, // @[:@16696.4]
  input   io_ins_1, // @[:@16696.4]
  output  io_outs_0, // @[:@16696.4]
  output  io_outs_1 // @[:@16696.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@16698.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@16699.4]
  reg [31:0] _RAND_1;
  wire  _T_23; // @[StickySelects.scala 49:53:@16700.4]
  wire  _T_24; // @[StickySelects.scala 49:21:@16701.4]
  wire  _T_25; // @[StickySelects.scala 49:53:@16703.4]
  wire  _T_26; // @[StickySelects.scala 49:21:@16704.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@16700.4]
  assign _T_24 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 49:21:@16701.4]
  assign _T_25 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@16703.4]
  assign _T_26 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 49:21:@16704.4]
  assign io_outs_0 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 53:57:@16706.4]
  assign io_outs_1 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 53:57:@16707.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_ins_1) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (io_ins_0) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_25;
      end
    end
  end
endmodule
module StickySelects_18( // @[:@16709.2]
  input   clock, // @[:@16710.4]
  input   reset, // @[:@16711.4]
  input   io_ins_0, // @[:@16712.4]
  input   io_ins_1, // @[:@16712.4]
  input   io_ins_2, // @[:@16712.4]
  input   io_ins_3, // @[:@16712.4]
  output  io_outs_0, // @[:@16712.4]
  output  io_outs_1, // @[:@16712.4]
  output  io_outs_2, // @[:@16712.4]
  output  io_outs_3 // @[:@16712.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@16714.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@16715.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@16716.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@16717.4]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[StickySelects.scala 47:46:@16718.4]
  wire  _T_30; // @[StickySelects.scala 47:46:@16719.4]
  wire  _T_31; // @[StickySelects.scala 49:53:@16720.4]
  wire  _T_32; // @[StickySelects.scala 49:21:@16721.4]
  wire  _T_33; // @[StickySelects.scala 47:46:@16723.4]
  wire  _T_34; // @[StickySelects.scala 47:46:@16724.4]
  wire  _T_35; // @[StickySelects.scala 49:53:@16725.4]
  wire  _T_36; // @[StickySelects.scala 49:21:@16726.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@16728.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@16729.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@16730.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@16731.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@16734.4]
  wire  _T_43; // @[StickySelects.scala 49:53:@16735.4]
  wire  _T_44; // @[StickySelects.scala 49:21:@16736.4]
  assign _T_29 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@16718.4]
  assign _T_30 = _T_29 | io_ins_3; // @[StickySelects.scala 47:46:@16719.4]
  assign _T_31 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@16720.4]
  assign _T_32 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 49:21:@16721.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@16723.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 47:46:@16724.4]
  assign _T_35 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@16725.4]
  assign _T_36 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 49:21:@16726.4]
  assign _T_37 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@16728.4]
  assign _T_38 = _T_37 | io_ins_3; // @[StickySelects.scala 47:46:@16729.4]
  assign _T_39 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@16730.4]
  assign _T_40 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 49:21:@16731.4]
  assign _T_42 = _T_37 | io_ins_2; // @[StickySelects.scala 47:46:@16734.4]
  assign _T_43 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@16735.4]
  assign _T_44 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 49:21:@16736.4]
  assign io_outs_0 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 53:57:@16738.4]
  assign io_outs_1 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 53:57:@16739.4]
  assign io_outs_2 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 53:57:@16740.4]
  assign io_outs_3 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 53:57:@16741.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_30) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_31;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_35;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_39;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_42) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_43;
      end
    end
  end
endmodule
module x302_lb2_0( // @[:@18629.2]
  input         clock, // @[:@18630.4]
  input         reset, // @[:@18631.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@18632.4]
  input         io_rPort_5_en_0, // @[:@18632.4]
  input         io_rPort_5_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_5_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@18632.4]
  input         io_rPort_4_en_0, // @[:@18632.4]
  input         io_rPort_4_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_4_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@18632.4]
  input         io_rPort_3_en_0, // @[:@18632.4]
  input         io_rPort_3_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_3_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@18632.4]
  input         io_rPort_2_en_0, // @[:@18632.4]
  input         io_rPort_2_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_2_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@18632.4]
  input         io_rPort_1_en_0, // @[:@18632.4]
  input         io_rPort_1_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_1_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@18632.4]
  input         io_rPort_0_en_0, // @[:@18632.4]
  input         io_rPort_0_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_0_output_0, // @[:@18632.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@18632.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@18632.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@18632.4]
  input  [31:0] io_wPort_1_data_0, // @[:@18632.4]
  input         io_wPort_1_en_0, // @[:@18632.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@18632.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@18632.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@18632.4]
  input  [31:0] io_wPort_0_data_0, // @[:@18632.4]
  input         io_wPort_0_en_0 // @[:@18632.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@20256.4]
  wire  _T_264; // @[MemPrimitives.scala 82:210:@18943.4]
  wire  _T_266; // @[MemPrimitives.scala 82:210:@18944.4]
  wire  _T_267; // @[MemPrimitives.scala 82:228:@18945.4]
  wire  _T_268; // @[MemPrimitives.scala 83:102:@18946.4]
  wire [41:0] _T_270; // @[Cat.scala 30:58:@18948.4]
  wire  _T_275; // @[MemPrimitives.scala 82:210:@18955.4]
  wire  _T_277; // @[MemPrimitives.scala 82:210:@18956.4]
  wire  _T_278; // @[MemPrimitives.scala 82:228:@18957.4]
  wire  _T_279; // @[MemPrimitives.scala 83:102:@18958.4]
  wire [41:0] _T_281; // @[Cat.scala 30:58:@18960.4]
  wire  _T_288; // @[MemPrimitives.scala 82:210:@18968.4]
  wire  _T_289; // @[MemPrimitives.scala 82:228:@18969.4]
  wire  _T_290; // @[MemPrimitives.scala 83:102:@18970.4]
  wire [41:0] _T_292; // @[Cat.scala 30:58:@18972.4]
  wire  _T_299; // @[MemPrimitives.scala 82:210:@18980.4]
  wire  _T_300; // @[MemPrimitives.scala 82:228:@18981.4]
  wire  _T_301; // @[MemPrimitives.scala 83:102:@18982.4]
  wire [41:0] _T_303; // @[Cat.scala 30:58:@18984.4]
  wire  _T_308; // @[MemPrimitives.scala 82:210:@18991.4]
  wire  _T_311; // @[MemPrimitives.scala 82:228:@18993.4]
  wire  _T_312; // @[MemPrimitives.scala 83:102:@18994.4]
  wire [41:0] _T_314; // @[Cat.scala 30:58:@18996.4]
  wire  _T_319; // @[MemPrimitives.scala 82:210:@19003.4]
  wire  _T_322; // @[MemPrimitives.scala 82:228:@19005.4]
  wire  _T_323; // @[MemPrimitives.scala 83:102:@19006.4]
  wire [41:0] _T_325; // @[Cat.scala 30:58:@19008.4]
  wire  _T_333; // @[MemPrimitives.scala 82:228:@19017.4]
  wire  _T_334; // @[MemPrimitives.scala 83:102:@19018.4]
  wire [41:0] _T_336; // @[Cat.scala 30:58:@19020.4]
  wire  _T_344; // @[MemPrimitives.scala 82:228:@19029.4]
  wire  _T_345; // @[MemPrimitives.scala 83:102:@19030.4]
  wire [41:0] _T_347; // @[Cat.scala 30:58:@19032.4]
  wire  _T_352; // @[MemPrimitives.scala 82:210:@19039.4]
  wire  _T_355; // @[MemPrimitives.scala 82:228:@19041.4]
  wire  _T_356; // @[MemPrimitives.scala 83:102:@19042.4]
  wire [41:0] _T_358; // @[Cat.scala 30:58:@19044.4]
  wire  _T_363; // @[MemPrimitives.scala 82:210:@19051.4]
  wire  _T_366; // @[MemPrimitives.scala 82:228:@19053.4]
  wire  _T_367; // @[MemPrimitives.scala 83:102:@19054.4]
  wire [41:0] _T_369; // @[Cat.scala 30:58:@19056.4]
  wire  _T_377; // @[MemPrimitives.scala 82:228:@19065.4]
  wire  _T_378; // @[MemPrimitives.scala 83:102:@19066.4]
  wire [41:0] _T_380; // @[Cat.scala 30:58:@19068.4]
  wire  _T_388; // @[MemPrimitives.scala 82:228:@19077.4]
  wire  _T_389; // @[MemPrimitives.scala 83:102:@19078.4]
  wire [41:0] _T_391; // @[Cat.scala 30:58:@19080.4]
  wire  _T_396; // @[MemPrimitives.scala 82:210:@19087.4]
  wire  _T_399; // @[MemPrimitives.scala 82:228:@19089.4]
  wire  _T_400; // @[MemPrimitives.scala 83:102:@19090.4]
  wire [41:0] _T_402; // @[Cat.scala 30:58:@19092.4]
  wire  _T_407; // @[MemPrimitives.scala 82:210:@19099.4]
  wire  _T_410; // @[MemPrimitives.scala 82:228:@19101.4]
  wire  _T_411; // @[MemPrimitives.scala 83:102:@19102.4]
  wire [41:0] _T_413; // @[Cat.scala 30:58:@19104.4]
  wire  _T_421; // @[MemPrimitives.scala 82:228:@19113.4]
  wire  _T_422; // @[MemPrimitives.scala 83:102:@19114.4]
  wire [41:0] _T_424; // @[Cat.scala 30:58:@19116.4]
  wire  _T_432; // @[MemPrimitives.scala 82:228:@19125.4]
  wire  _T_433; // @[MemPrimitives.scala 83:102:@19126.4]
  wire [41:0] _T_435; // @[Cat.scala 30:58:@19128.4]
  wire  _T_440; // @[MemPrimitives.scala 110:210:@19135.4]
  wire  _T_442; // @[MemPrimitives.scala 110:210:@19136.4]
  wire  _T_443; // @[MemPrimitives.scala 110:228:@19137.4]
  wire  _T_446; // @[MemPrimitives.scala 110:210:@19139.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@19140.4]
  wire  _T_449; // @[MemPrimitives.scala 110:228:@19141.4]
  wire  _T_451; // @[MemPrimitives.scala 126:35:@19148.4]
  wire  _T_452; // @[MemPrimitives.scala 126:35:@19149.4]
  wire [10:0] _T_454; // @[Cat.scala 30:58:@19151.4]
  wire [10:0] _T_456; // @[Cat.scala 30:58:@19153.4]
  wire [10:0] _T_457; // @[Mux.scala 31:69:@19154.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@19161.4]
  wire  _T_464; // @[MemPrimitives.scala 110:210:@19162.4]
  wire  _T_465; // @[MemPrimitives.scala 110:228:@19163.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@19165.4]
  wire  _T_470; // @[MemPrimitives.scala 110:210:@19166.4]
  wire  _T_471; // @[MemPrimitives.scala 110:228:@19167.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@19169.4]
  wire  _T_476; // @[MemPrimitives.scala 110:210:@19170.4]
  wire  _T_477; // @[MemPrimitives.scala 110:228:@19171.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@19173.4]
  wire  _T_482; // @[MemPrimitives.scala 110:210:@19174.4]
  wire  _T_483; // @[MemPrimitives.scala 110:228:@19175.4]
  wire  _T_485; // @[MemPrimitives.scala 126:35:@19184.4]
  wire  _T_486; // @[MemPrimitives.scala 126:35:@19185.4]
  wire  _T_487; // @[MemPrimitives.scala 126:35:@19186.4]
  wire  _T_488; // @[MemPrimitives.scala 126:35:@19187.4]
  wire [10:0] _T_490; // @[Cat.scala 30:58:@19189.4]
  wire [10:0] _T_492; // @[Cat.scala 30:58:@19191.4]
  wire [10:0] _T_494; // @[Cat.scala 30:58:@19193.4]
  wire [10:0] _T_496; // @[Cat.scala 30:58:@19195.4]
  wire [10:0] _T_497; // @[Mux.scala 31:69:@19196.4]
  wire [10:0] _T_498; // @[Mux.scala 31:69:@19197.4]
  wire [10:0] _T_499; // @[Mux.scala 31:69:@19198.4]
  wire  _T_506; // @[MemPrimitives.scala 110:210:@19206.4]
  wire  _T_507; // @[MemPrimitives.scala 110:228:@19207.4]
  wire  _T_512; // @[MemPrimitives.scala 110:210:@19210.4]
  wire  _T_513; // @[MemPrimitives.scala 110:228:@19211.4]
  wire  _T_515; // @[MemPrimitives.scala 126:35:@19218.4]
  wire  _T_516; // @[MemPrimitives.scala 126:35:@19219.4]
  wire [10:0] _T_518; // @[Cat.scala 30:58:@19221.4]
  wire [10:0] _T_520; // @[Cat.scala 30:58:@19223.4]
  wire [10:0] _T_521; // @[Mux.scala 31:69:@19224.4]
  wire  _T_528; // @[MemPrimitives.scala 110:210:@19232.4]
  wire  _T_529; // @[MemPrimitives.scala 110:228:@19233.4]
  wire  _T_534; // @[MemPrimitives.scala 110:210:@19236.4]
  wire  _T_535; // @[MemPrimitives.scala 110:228:@19237.4]
  wire  _T_540; // @[MemPrimitives.scala 110:210:@19240.4]
  wire  _T_541; // @[MemPrimitives.scala 110:228:@19241.4]
  wire  _T_546; // @[MemPrimitives.scala 110:210:@19244.4]
  wire  _T_547; // @[MemPrimitives.scala 110:228:@19245.4]
  wire  _T_549; // @[MemPrimitives.scala 126:35:@19254.4]
  wire  _T_550; // @[MemPrimitives.scala 126:35:@19255.4]
  wire  _T_551; // @[MemPrimitives.scala 126:35:@19256.4]
  wire  _T_552; // @[MemPrimitives.scala 126:35:@19257.4]
  wire [10:0] _T_554; // @[Cat.scala 30:58:@19259.4]
  wire [10:0] _T_556; // @[Cat.scala 30:58:@19261.4]
  wire [10:0] _T_558; // @[Cat.scala 30:58:@19263.4]
  wire [10:0] _T_560; // @[Cat.scala 30:58:@19265.4]
  wire [10:0] _T_561; // @[Mux.scala 31:69:@19266.4]
  wire [10:0] _T_562; // @[Mux.scala 31:69:@19267.4]
  wire [10:0] _T_563; // @[Mux.scala 31:69:@19268.4]
  wire  _T_568; // @[MemPrimitives.scala 110:210:@19275.4]
  wire  _T_571; // @[MemPrimitives.scala 110:228:@19277.4]
  wire  _T_574; // @[MemPrimitives.scala 110:210:@19279.4]
  wire  _T_577; // @[MemPrimitives.scala 110:228:@19281.4]
  wire  _T_579; // @[MemPrimitives.scala 126:35:@19288.4]
  wire  _T_580; // @[MemPrimitives.scala 126:35:@19289.4]
  wire [10:0] _T_582; // @[Cat.scala 30:58:@19291.4]
  wire [10:0] _T_584; // @[Cat.scala 30:58:@19293.4]
  wire [10:0] _T_585; // @[Mux.scala 31:69:@19294.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@19301.4]
  wire  _T_593; // @[MemPrimitives.scala 110:228:@19303.4]
  wire  _T_596; // @[MemPrimitives.scala 110:210:@19305.4]
  wire  _T_599; // @[MemPrimitives.scala 110:228:@19307.4]
  wire  _T_602; // @[MemPrimitives.scala 110:210:@19309.4]
  wire  _T_605; // @[MemPrimitives.scala 110:228:@19311.4]
  wire  _T_608; // @[MemPrimitives.scala 110:210:@19313.4]
  wire  _T_611; // @[MemPrimitives.scala 110:228:@19315.4]
  wire  _T_613; // @[MemPrimitives.scala 126:35:@19324.4]
  wire  _T_614; // @[MemPrimitives.scala 126:35:@19325.4]
  wire  _T_615; // @[MemPrimitives.scala 126:35:@19326.4]
  wire  _T_616; // @[MemPrimitives.scala 126:35:@19327.4]
  wire [10:0] _T_618; // @[Cat.scala 30:58:@19329.4]
  wire [10:0] _T_620; // @[Cat.scala 30:58:@19331.4]
  wire [10:0] _T_622; // @[Cat.scala 30:58:@19333.4]
  wire [10:0] _T_624; // @[Cat.scala 30:58:@19335.4]
  wire [10:0] _T_625; // @[Mux.scala 31:69:@19336.4]
  wire [10:0] _T_626; // @[Mux.scala 31:69:@19337.4]
  wire [10:0] _T_627; // @[Mux.scala 31:69:@19338.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@19347.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@19351.4]
  wire  _T_643; // @[MemPrimitives.scala 126:35:@19358.4]
  wire  _T_644; // @[MemPrimitives.scala 126:35:@19359.4]
  wire [10:0] _T_646; // @[Cat.scala 30:58:@19361.4]
  wire [10:0] _T_648; // @[Cat.scala 30:58:@19363.4]
  wire [10:0] _T_649; // @[Mux.scala 31:69:@19364.4]
  wire  _T_657; // @[MemPrimitives.scala 110:228:@19373.4]
  wire  _T_663; // @[MemPrimitives.scala 110:228:@19377.4]
  wire  _T_669; // @[MemPrimitives.scala 110:228:@19381.4]
  wire  _T_675; // @[MemPrimitives.scala 110:228:@19385.4]
  wire  _T_677; // @[MemPrimitives.scala 126:35:@19394.4]
  wire  _T_678; // @[MemPrimitives.scala 126:35:@19395.4]
  wire  _T_679; // @[MemPrimitives.scala 126:35:@19396.4]
  wire  _T_680; // @[MemPrimitives.scala 126:35:@19397.4]
  wire [10:0] _T_682; // @[Cat.scala 30:58:@19399.4]
  wire [10:0] _T_684; // @[Cat.scala 30:58:@19401.4]
  wire [10:0] _T_686; // @[Cat.scala 30:58:@19403.4]
  wire [10:0] _T_688; // @[Cat.scala 30:58:@19405.4]
  wire [10:0] _T_689; // @[Mux.scala 31:69:@19406.4]
  wire [10:0] _T_690; // @[Mux.scala 31:69:@19407.4]
  wire [10:0] _T_691; // @[Mux.scala 31:69:@19408.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@19415.4]
  wire  _T_699; // @[MemPrimitives.scala 110:228:@19417.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@19419.4]
  wire  _T_705; // @[MemPrimitives.scala 110:228:@19421.4]
  wire  _T_707; // @[MemPrimitives.scala 126:35:@19428.4]
  wire  _T_708; // @[MemPrimitives.scala 126:35:@19429.4]
  wire [10:0] _T_710; // @[Cat.scala 30:58:@19431.4]
  wire [10:0] _T_712; // @[Cat.scala 30:58:@19433.4]
  wire [10:0] _T_713; // @[Mux.scala 31:69:@19434.4]
  wire  _T_718; // @[MemPrimitives.scala 110:210:@19441.4]
  wire  _T_721; // @[MemPrimitives.scala 110:228:@19443.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@19445.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@19447.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@19449.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@19451.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@19453.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@19455.4]
  wire  _T_741; // @[MemPrimitives.scala 126:35:@19464.4]
  wire  _T_742; // @[MemPrimitives.scala 126:35:@19465.4]
  wire  _T_743; // @[MemPrimitives.scala 126:35:@19466.4]
  wire  _T_744; // @[MemPrimitives.scala 126:35:@19467.4]
  wire [10:0] _T_746; // @[Cat.scala 30:58:@19469.4]
  wire [10:0] _T_748; // @[Cat.scala 30:58:@19471.4]
  wire [10:0] _T_750; // @[Cat.scala 30:58:@19473.4]
  wire [10:0] _T_752; // @[Cat.scala 30:58:@19475.4]
  wire [10:0] _T_753; // @[Mux.scala 31:69:@19476.4]
  wire [10:0] _T_754; // @[Mux.scala 31:69:@19477.4]
  wire [10:0] _T_755; // @[Mux.scala 31:69:@19478.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@19487.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@19491.4]
  wire  _T_771; // @[MemPrimitives.scala 126:35:@19498.4]
  wire  _T_772; // @[MemPrimitives.scala 126:35:@19499.4]
  wire [10:0] _T_774; // @[Cat.scala 30:58:@19501.4]
  wire [10:0] _T_776; // @[Cat.scala 30:58:@19503.4]
  wire [10:0] _T_777; // @[Mux.scala 31:69:@19504.4]
  wire  _T_785; // @[MemPrimitives.scala 110:228:@19513.4]
  wire  _T_791; // @[MemPrimitives.scala 110:228:@19517.4]
  wire  _T_797; // @[MemPrimitives.scala 110:228:@19521.4]
  wire  _T_803; // @[MemPrimitives.scala 110:228:@19525.4]
  wire  _T_805; // @[MemPrimitives.scala 126:35:@19534.4]
  wire  _T_806; // @[MemPrimitives.scala 126:35:@19535.4]
  wire  _T_807; // @[MemPrimitives.scala 126:35:@19536.4]
  wire  _T_808; // @[MemPrimitives.scala 126:35:@19537.4]
  wire [10:0] _T_810; // @[Cat.scala 30:58:@19539.4]
  wire [10:0] _T_812; // @[Cat.scala 30:58:@19541.4]
  wire [10:0] _T_814; // @[Cat.scala 30:58:@19543.4]
  wire [10:0] _T_816; // @[Cat.scala 30:58:@19545.4]
  wire [10:0] _T_817; // @[Mux.scala 31:69:@19546.4]
  wire [10:0] _T_818; // @[Mux.scala 31:69:@19547.4]
  wire [10:0] _T_819; // @[Mux.scala 31:69:@19548.4]
  wire  _T_824; // @[MemPrimitives.scala 110:210:@19555.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@19557.4]
  wire  _T_830; // @[MemPrimitives.scala 110:210:@19559.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@19561.4]
  wire  _T_835; // @[MemPrimitives.scala 126:35:@19568.4]
  wire  _T_836; // @[MemPrimitives.scala 126:35:@19569.4]
  wire [10:0] _T_838; // @[Cat.scala 30:58:@19571.4]
  wire [10:0] _T_840; // @[Cat.scala 30:58:@19573.4]
  wire [10:0] _T_841; // @[Mux.scala 31:69:@19574.4]
  wire  _T_846; // @[MemPrimitives.scala 110:210:@19581.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@19583.4]
  wire  _T_852; // @[MemPrimitives.scala 110:210:@19585.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@19587.4]
  wire  _T_858; // @[MemPrimitives.scala 110:210:@19589.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@19591.4]
  wire  _T_864; // @[MemPrimitives.scala 110:210:@19593.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@19595.4]
  wire  _T_869; // @[MemPrimitives.scala 126:35:@19604.4]
  wire  _T_870; // @[MemPrimitives.scala 126:35:@19605.4]
  wire  _T_871; // @[MemPrimitives.scala 126:35:@19606.4]
  wire  _T_872; // @[MemPrimitives.scala 126:35:@19607.4]
  wire [10:0] _T_874; // @[Cat.scala 30:58:@19609.4]
  wire [10:0] _T_876; // @[Cat.scala 30:58:@19611.4]
  wire [10:0] _T_878; // @[Cat.scala 30:58:@19613.4]
  wire [10:0] _T_880; // @[Cat.scala 30:58:@19615.4]
  wire [10:0] _T_881; // @[Mux.scala 31:69:@19616.4]
  wire [10:0] _T_882; // @[Mux.scala 31:69:@19617.4]
  wire [10:0] _T_883; // @[Mux.scala 31:69:@19618.4]
  wire  _T_891; // @[MemPrimitives.scala 110:228:@19627.4]
  wire  _T_897; // @[MemPrimitives.scala 110:228:@19631.4]
  wire  _T_899; // @[MemPrimitives.scala 126:35:@19638.4]
  wire  _T_900; // @[MemPrimitives.scala 126:35:@19639.4]
  wire [10:0] _T_902; // @[Cat.scala 30:58:@19641.4]
  wire [10:0] _T_904; // @[Cat.scala 30:58:@19643.4]
  wire [10:0] _T_905; // @[Mux.scala 31:69:@19644.4]
  wire  _T_913; // @[MemPrimitives.scala 110:228:@19653.4]
  wire  _T_919; // @[MemPrimitives.scala 110:228:@19657.4]
  wire  _T_925; // @[MemPrimitives.scala 110:228:@19661.4]
  wire  _T_931; // @[MemPrimitives.scala 110:228:@19665.4]
  wire  _T_933; // @[MemPrimitives.scala 126:35:@19674.4]
  wire  _T_934; // @[MemPrimitives.scala 126:35:@19675.4]
  wire  _T_935; // @[MemPrimitives.scala 126:35:@19676.4]
  wire  _T_936; // @[MemPrimitives.scala 126:35:@19677.4]
  wire [10:0] _T_938; // @[Cat.scala 30:58:@19679.4]
  wire [10:0] _T_940; // @[Cat.scala 30:58:@19681.4]
  wire [10:0] _T_942; // @[Cat.scala 30:58:@19683.4]
  wire [10:0] _T_944; // @[Cat.scala 30:58:@19685.4]
  wire [10:0] _T_945; // @[Mux.scala 31:69:@19686.4]
  wire [10:0] _T_946; // @[Mux.scala 31:69:@19687.4]
  wire [10:0] _T_947; // @[Mux.scala 31:69:@19688.4]
  wire  _T_1011; // @[package.scala 96:25:@19773.4 package.scala 96:25:@19774.4]
  wire [31:0] _T_1015; // @[Mux.scala 31:69:@19783.4]
  wire  _T_1008; // @[package.scala 96:25:@19765.4 package.scala 96:25:@19766.4]
  wire [31:0] _T_1016; // @[Mux.scala 31:69:@19784.4]
  wire  _T_1005; // @[package.scala 96:25:@19757.4 package.scala 96:25:@19758.4]
  wire [31:0] _T_1017; // @[Mux.scala 31:69:@19785.4]
  wire  _T_1002; // @[package.scala 96:25:@19749.4 package.scala 96:25:@19750.4]
  wire [31:0] _T_1018; // @[Mux.scala 31:69:@19786.4]
  wire  _T_999; // @[package.scala 96:25:@19741.4 package.scala 96:25:@19742.4]
  wire [31:0] _T_1019; // @[Mux.scala 31:69:@19787.4]
  wire  _T_996; // @[package.scala 96:25:@19733.4 package.scala 96:25:@19734.4]
  wire [31:0] _T_1020; // @[Mux.scala 31:69:@19788.4]
  wire  _T_993; // @[package.scala 96:25:@19725.4 package.scala 96:25:@19726.4]
  wire  _T_1082; // @[package.scala 96:25:@19869.4 package.scala 96:25:@19870.4]
  wire [31:0] _T_1086; // @[Mux.scala 31:69:@19879.4]
  wire  _T_1079; // @[package.scala 96:25:@19861.4 package.scala 96:25:@19862.4]
  wire [31:0] _T_1087; // @[Mux.scala 31:69:@19880.4]
  wire  _T_1076; // @[package.scala 96:25:@19853.4 package.scala 96:25:@19854.4]
  wire [31:0] _T_1088; // @[Mux.scala 31:69:@19881.4]
  wire  _T_1073; // @[package.scala 96:25:@19845.4 package.scala 96:25:@19846.4]
  wire [31:0] _T_1089; // @[Mux.scala 31:69:@19882.4]
  wire  _T_1070; // @[package.scala 96:25:@19837.4 package.scala 96:25:@19838.4]
  wire [31:0] _T_1090; // @[Mux.scala 31:69:@19883.4]
  wire  _T_1067; // @[package.scala 96:25:@19829.4 package.scala 96:25:@19830.4]
  wire [31:0] _T_1091; // @[Mux.scala 31:69:@19884.4]
  wire  _T_1064; // @[package.scala 96:25:@19821.4 package.scala 96:25:@19822.4]
  wire  _T_1153; // @[package.scala 96:25:@19965.4 package.scala 96:25:@19966.4]
  wire [31:0] _T_1157; // @[Mux.scala 31:69:@19975.4]
  wire  _T_1150; // @[package.scala 96:25:@19957.4 package.scala 96:25:@19958.4]
  wire [31:0] _T_1158; // @[Mux.scala 31:69:@19976.4]
  wire  _T_1147; // @[package.scala 96:25:@19949.4 package.scala 96:25:@19950.4]
  wire [31:0] _T_1159; // @[Mux.scala 31:69:@19977.4]
  wire  _T_1144; // @[package.scala 96:25:@19941.4 package.scala 96:25:@19942.4]
  wire [31:0] _T_1160; // @[Mux.scala 31:69:@19978.4]
  wire  _T_1141; // @[package.scala 96:25:@19933.4 package.scala 96:25:@19934.4]
  wire [31:0] _T_1161; // @[Mux.scala 31:69:@19979.4]
  wire  _T_1138; // @[package.scala 96:25:@19925.4 package.scala 96:25:@19926.4]
  wire [31:0] _T_1162; // @[Mux.scala 31:69:@19980.4]
  wire  _T_1135; // @[package.scala 96:25:@19917.4 package.scala 96:25:@19918.4]
  wire  _T_1224; // @[package.scala 96:25:@20061.4 package.scala 96:25:@20062.4]
  wire [31:0] _T_1228; // @[Mux.scala 31:69:@20071.4]
  wire  _T_1221; // @[package.scala 96:25:@20053.4 package.scala 96:25:@20054.4]
  wire [31:0] _T_1229; // @[Mux.scala 31:69:@20072.4]
  wire  _T_1218; // @[package.scala 96:25:@20045.4 package.scala 96:25:@20046.4]
  wire [31:0] _T_1230; // @[Mux.scala 31:69:@20073.4]
  wire  _T_1215; // @[package.scala 96:25:@20037.4 package.scala 96:25:@20038.4]
  wire [31:0] _T_1231; // @[Mux.scala 31:69:@20074.4]
  wire  _T_1212; // @[package.scala 96:25:@20029.4 package.scala 96:25:@20030.4]
  wire [31:0] _T_1232; // @[Mux.scala 31:69:@20075.4]
  wire  _T_1209; // @[package.scala 96:25:@20021.4 package.scala 96:25:@20022.4]
  wire [31:0] _T_1233; // @[Mux.scala 31:69:@20076.4]
  wire  _T_1206; // @[package.scala 96:25:@20013.4 package.scala 96:25:@20014.4]
  wire  _T_1295; // @[package.scala 96:25:@20157.4 package.scala 96:25:@20158.4]
  wire [31:0] _T_1299; // @[Mux.scala 31:69:@20167.4]
  wire  _T_1292; // @[package.scala 96:25:@20149.4 package.scala 96:25:@20150.4]
  wire [31:0] _T_1300; // @[Mux.scala 31:69:@20168.4]
  wire  _T_1289; // @[package.scala 96:25:@20141.4 package.scala 96:25:@20142.4]
  wire [31:0] _T_1301; // @[Mux.scala 31:69:@20169.4]
  wire  _T_1286; // @[package.scala 96:25:@20133.4 package.scala 96:25:@20134.4]
  wire [31:0] _T_1302; // @[Mux.scala 31:69:@20170.4]
  wire  _T_1283; // @[package.scala 96:25:@20125.4 package.scala 96:25:@20126.4]
  wire [31:0] _T_1303; // @[Mux.scala 31:69:@20171.4]
  wire  _T_1280; // @[package.scala 96:25:@20117.4 package.scala 96:25:@20118.4]
  wire [31:0] _T_1304; // @[Mux.scala 31:69:@20172.4]
  wire  _T_1277; // @[package.scala 96:25:@20109.4 package.scala 96:25:@20110.4]
  wire  _T_1366; // @[package.scala 96:25:@20253.4 package.scala 96:25:@20254.4]
  wire [31:0] _T_1370; // @[Mux.scala 31:69:@20263.4]
  wire  _T_1363; // @[package.scala 96:25:@20245.4 package.scala 96:25:@20246.4]
  wire [31:0] _T_1371; // @[Mux.scala 31:69:@20264.4]
  wire  _T_1360; // @[package.scala 96:25:@20237.4 package.scala 96:25:@20238.4]
  wire [31:0] _T_1372; // @[Mux.scala 31:69:@20265.4]
  wire  _T_1357; // @[package.scala 96:25:@20229.4 package.scala 96:25:@20230.4]
  wire [31:0] _T_1373; // @[Mux.scala 31:69:@20266.4]
  wire  _T_1354; // @[package.scala 96:25:@20221.4 package.scala 96:25:@20222.4]
  wire [31:0] _T_1374; // @[Mux.scala 31:69:@20267.4]
  wire  _T_1351; // @[package.scala 96:25:@20213.4 package.scala 96:25:@20214.4]
  wire [31:0] _T_1375; // @[Mux.scala 31:69:@20268.4]
  wire  _T_1348; // @[package.scala 96:25:@20205.4 package.scala 96:25:@20206.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@18687.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@18703.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@18719.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@18735.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@18751.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@18767.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@18783.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@18799.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@18815.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@18831.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@18847.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@18863.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@18879.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@18895.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@18911.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@18927.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_17 StickySelects ( // @[MemPrimitives.scala 124:33:@19143.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1)
  );
  StickySelects_18 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@19177.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_17 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@19213.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1)
  );
  StickySelects_18 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@19247.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3)
  );
  StickySelects_17 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@19283.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1)
  );
  StickySelects_18 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@19317.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_17 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@19353.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1)
  );
  StickySelects_18 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@19387.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3)
  );
  StickySelects_17 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@19423.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1)
  );
  StickySelects_18 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@19457.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_17 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@19493.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1)
  );
  StickySelects_18 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@19527.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3)
  );
  StickySelects_17 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@19563.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1)
  );
  StickySelects_18 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@19597.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3)
  );
  StickySelects_17 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@19633.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1)
  );
  StickySelects_18 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@19667.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@19720.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@19728.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@19736.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@19744.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@19752.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@19760.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@19768.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@19776.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@19816.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@19824.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@19832.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@19840.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@19848.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@19856.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@19864.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@19872.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@19912.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@19920.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@19928.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@19936.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@19944.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@19952.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@19960.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@19968.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@20008.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@20016.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@20024.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@20032.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@20040.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@20048.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@20056.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@20064.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@20104.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@20112.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@20120.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@20128.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@20136.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@20144.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@20152.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@20160.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@20200.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@20208.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@20216.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@20224.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@20232.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@20240.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@20248.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@20256.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  assign _T_264 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@18943.4]
  assign _T_266 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@18944.4]
  assign _T_267 = _T_264 & _T_266; // @[MemPrimitives.scala 82:228:@18945.4]
  assign _T_268 = io_wPort_0_en_0 & _T_267; // @[MemPrimitives.scala 83:102:@18946.4]
  assign _T_270 = {_T_268,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18948.4]
  assign _T_275 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@18955.4]
  assign _T_277 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@18956.4]
  assign _T_278 = _T_275 & _T_277; // @[MemPrimitives.scala 82:228:@18957.4]
  assign _T_279 = io_wPort_1_en_0 & _T_278; // @[MemPrimitives.scala 83:102:@18958.4]
  assign _T_281 = {_T_279,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@18960.4]
  assign _T_288 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@18968.4]
  assign _T_289 = _T_264 & _T_288; // @[MemPrimitives.scala 82:228:@18969.4]
  assign _T_290 = io_wPort_0_en_0 & _T_289; // @[MemPrimitives.scala 83:102:@18970.4]
  assign _T_292 = {_T_290,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18972.4]
  assign _T_299 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@18980.4]
  assign _T_300 = _T_275 & _T_299; // @[MemPrimitives.scala 82:228:@18981.4]
  assign _T_301 = io_wPort_1_en_0 & _T_300; // @[MemPrimitives.scala 83:102:@18982.4]
  assign _T_303 = {_T_301,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@18984.4]
  assign _T_308 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@18991.4]
  assign _T_311 = _T_308 & _T_266; // @[MemPrimitives.scala 82:228:@18993.4]
  assign _T_312 = io_wPort_0_en_0 & _T_311; // @[MemPrimitives.scala 83:102:@18994.4]
  assign _T_314 = {_T_312,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18996.4]
  assign _T_319 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@19003.4]
  assign _T_322 = _T_319 & _T_277; // @[MemPrimitives.scala 82:228:@19005.4]
  assign _T_323 = io_wPort_1_en_0 & _T_322; // @[MemPrimitives.scala 83:102:@19006.4]
  assign _T_325 = {_T_323,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19008.4]
  assign _T_333 = _T_308 & _T_288; // @[MemPrimitives.scala 82:228:@19017.4]
  assign _T_334 = io_wPort_0_en_0 & _T_333; // @[MemPrimitives.scala 83:102:@19018.4]
  assign _T_336 = {_T_334,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19020.4]
  assign _T_344 = _T_319 & _T_299; // @[MemPrimitives.scala 82:228:@19029.4]
  assign _T_345 = io_wPort_1_en_0 & _T_344; // @[MemPrimitives.scala 83:102:@19030.4]
  assign _T_347 = {_T_345,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19032.4]
  assign _T_352 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@19039.4]
  assign _T_355 = _T_352 & _T_266; // @[MemPrimitives.scala 82:228:@19041.4]
  assign _T_356 = io_wPort_0_en_0 & _T_355; // @[MemPrimitives.scala 83:102:@19042.4]
  assign _T_358 = {_T_356,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19044.4]
  assign _T_363 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@19051.4]
  assign _T_366 = _T_363 & _T_277; // @[MemPrimitives.scala 82:228:@19053.4]
  assign _T_367 = io_wPort_1_en_0 & _T_366; // @[MemPrimitives.scala 83:102:@19054.4]
  assign _T_369 = {_T_367,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19056.4]
  assign _T_377 = _T_352 & _T_288; // @[MemPrimitives.scala 82:228:@19065.4]
  assign _T_378 = io_wPort_0_en_0 & _T_377; // @[MemPrimitives.scala 83:102:@19066.4]
  assign _T_380 = {_T_378,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19068.4]
  assign _T_388 = _T_363 & _T_299; // @[MemPrimitives.scala 82:228:@19077.4]
  assign _T_389 = io_wPort_1_en_0 & _T_388; // @[MemPrimitives.scala 83:102:@19078.4]
  assign _T_391 = {_T_389,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19080.4]
  assign _T_396 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@19087.4]
  assign _T_399 = _T_396 & _T_266; // @[MemPrimitives.scala 82:228:@19089.4]
  assign _T_400 = io_wPort_0_en_0 & _T_399; // @[MemPrimitives.scala 83:102:@19090.4]
  assign _T_402 = {_T_400,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19092.4]
  assign _T_407 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@19099.4]
  assign _T_410 = _T_407 & _T_277; // @[MemPrimitives.scala 82:228:@19101.4]
  assign _T_411 = io_wPort_1_en_0 & _T_410; // @[MemPrimitives.scala 83:102:@19102.4]
  assign _T_413 = {_T_411,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19104.4]
  assign _T_421 = _T_396 & _T_288; // @[MemPrimitives.scala 82:228:@19113.4]
  assign _T_422 = io_wPort_0_en_0 & _T_421; // @[MemPrimitives.scala 83:102:@19114.4]
  assign _T_424 = {_T_422,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19116.4]
  assign _T_432 = _T_407 & _T_299; // @[MemPrimitives.scala 82:228:@19125.4]
  assign _T_433 = io_wPort_1_en_0 & _T_432; // @[MemPrimitives.scala 83:102:@19126.4]
  assign _T_435 = {_T_433,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19128.4]
  assign _T_440 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19135.4]
  assign _T_442 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@19136.4]
  assign _T_443 = _T_440 & _T_442; // @[MemPrimitives.scala 110:228:@19137.4]
  assign _T_446 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19139.4]
  assign _T_448 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@19140.4]
  assign _T_449 = _T_446 & _T_448; // @[MemPrimitives.scala 110:228:@19141.4]
  assign _T_451 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@19148.4]
  assign _T_452 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@19149.4]
  assign _T_454 = {_T_451,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19151.4]
  assign _T_456 = {_T_452,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19153.4]
  assign _T_457 = _T_451 ? _T_454 : _T_456; // @[Mux.scala 31:69:@19154.4]
  assign _T_462 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19161.4]
  assign _T_464 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19162.4]
  assign _T_465 = _T_462 & _T_464; // @[MemPrimitives.scala 110:228:@19163.4]
  assign _T_468 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19165.4]
  assign _T_470 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19166.4]
  assign _T_471 = _T_468 & _T_470; // @[MemPrimitives.scala 110:228:@19167.4]
  assign _T_474 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19169.4]
  assign _T_476 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19170.4]
  assign _T_477 = _T_474 & _T_476; // @[MemPrimitives.scala 110:228:@19171.4]
  assign _T_480 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19173.4]
  assign _T_482 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19174.4]
  assign _T_483 = _T_480 & _T_482; // @[MemPrimitives.scala 110:228:@19175.4]
  assign _T_485 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@19184.4]
  assign _T_486 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@19185.4]
  assign _T_487 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@19186.4]
  assign _T_488 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@19187.4]
  assign _T_490 = {_T_485,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19189.4]
  assign _T_492 = {_T_486,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19191.4]
  assign _T_494 = {_T_487,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19193.4]
  assign _T_496 = {_T_488,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19195.4]
  assign _T_497 = _T_487 ? _T_494 : _T_496; // @[Mux.scala 31:69:@19196.4]
  assign _T_498 = _T_486 ? _T_492 : _T_497; // @[Mux.scala 31:69:@19197.4]
  assign _T_499 = _T_485 ? _T_490 : _T_498; // @[Mux.scala 31:69:@19198.4]
  assign _T_506 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@19206.4]
  assign _T_507 = _T_440 & _T_506; // @[MemPrimitives.scala 110:228:@19207.4]
  assign _T_512 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@19210.4]
  assign _T_513 = _T_446 & _T_512; // @[MemPrimitives.scala 110:228:@19211.4]
  assign _T_515 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@19218.4]
  assign _T_516 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@19219.4]
  assign _T_518 = {_T_515,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19221.4]
  assign _T_520 = {_T_516,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19223.4]
  assign _T_521 = _T_515 ? _T_518 : _T_520; // @[Mux.scala 31:69:@19224.4]
  assign _T_528 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19232.4]
  assign _T_529 = _T_462 & _T_528; // @[MemPrimitives.scala 110:228:@19233.4]
  assign _T_534 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19236.4]
  assign _T_535 = _T_468 & _T_534; // @[MemPrimitives.scala 110:228:@19237.4]
  assign _T_540 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19240.4]
  assign _T_541 = _T_474 & _T_540; // @[MemPrimitives.scala 110:228:@19241.4]
  assign _T_546 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19244.4]
  assign _T_547 = _T_480 & _T_546; // @[MemPrimitives.scala 110:228:@19245.4]
  assign _T_549 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@19254.4]
  assign _T_550 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@19255.4]
  assign _T_551 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@19256.4]
  assign _T_552 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@19257.4]
  assign _T_554 = {_T_549,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19259.4]
  assign _T_556 = {_T_550,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19261.4]
  assign _T_558 = {_T_551,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19263.4]
  assign _T_560 = {_T_552,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19265.4]
  assign _T_561 = _T_551 ? _T_558 : _T_560; // @[Mux.scala 31:69:@19266.4]
  assign _T_562 = _T_550 ? _T_556 : _T_561; // @[Mux.scala 31:69:@19267.4]
  assign _T_563 = _T_549 ? _T_554 : _T_562; // @[Mux.scala 31:69:@19268.4]
  assign _T_568 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19275.4]
  assign _T_571 = _T_568 & _T_442; // @[MemPrimitives.scala 110:228:@19277.4]
  assign _T_574 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19279.4]
  assign _T_577 = _T_574 & _T_448; // @[MemPrimitives.scala 110:228:@19281.4]
  assign _T_579 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@19288.4]
  assign _T_580 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@19289.4]
  assign _T_582 = {_T_579,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19291.4]
  assign _T_584 = {_T_580,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19293.4]
  assign _T_585 = _T_579 ? _T_582 : _T_584; // @[Mux.scala 31:69:@19294.4]
  assign _T_590 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19301.4]
  assign _T_593 = _T_590 & _T_464; // @[MemPrimitives.scala 110:228:@19303.4]
  assign _T_596 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19305.4]
  assign _T_599 = _T_596 & _T_470; // @[MemPrimitives.scala 110:228:@19307.4]
  assign _T_602 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19309.4]
  assign _T_605 = _T_602 & _T_476; // @[MemPrimitives.scala 110:228:@19311.4]
  assign _T_608 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19313.4]
  assign _T_611 = _T_608 & _T_482; // @[MemPrimitives.scala 110:228:@19315.4]
  assign _T_613 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@19324.4]
  assign _T_614 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@19325.4]
  assign _T_615 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@19326.4]
  assign _T_616 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@19327.4]
  assign _T_618 = {_T_613,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19329.4]
  assign _T_620 = {_T_614,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19331.4]
  assign _T_622 = {_T_615,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19333.4]
  assign _T_624 = {_T_616,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19335.4]
  assign _T_625 = _T_615 ? _T_622 : _T_624; // @[Mux.scala 31:69:@19336.4]
  assign _T_626 = _T_614 ? _T_620 : _T_625; // @[Mux.scala 31:69:@19337.4]
  assign _T_627 = _T_613 ? _T_618 : _T_626; // @[Mux.scala 31:69:@19338.4]
  assign _T_635 = _T_568 & _T_506; // @[MemPrimitives.scala 110:228:@19347.4]
  assign _T_641 = _T_574 & _T_512; // @[MemPrimitives.scala 110:228:@19351.4]
  assign _T_643 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@19358.4]
  assign _T_644 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@19359.4]
  assign _T_646 = {_T_643,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19361.4]
  assign _T_648 = {_T_644,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19363.4]
  assign _T_649 = _T_643 ? _T_646 : _T_648; // @[Mux.scala 31:69:@19364.4]
  assign _T_657 = _T_590 & _T_528; // @[MemPrimitives.scala 110:228:@19373.4]
  assign _T_663 = _T_596 & _T_534; // @[MemPrimitives.scala 110:228:@19377.4]
  assign _T_669 = _T_602 & _T_540; // @[MemPrimitives.scala 110:228:@19381.4]
  assign _T_675 = _T_608 & _T_546; // @[MemPrimitives.scala 110:228:@19385.4]
  assign _T_677 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@19394.4]
  assign _T_678 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@19395.4]
  assign _T_679 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@19396.4]
  assign _T_680 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@19397.4]
  assign _T_682 = {_T_677,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19399.4]
  assign _T_684 = {_T_678,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19401.4]
  assign _T_686 = {_T_679,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19403.4]
  assign _T_688 = {_T_680,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19405.4]
  assign _T_689 = _T_679 ? _T_686 : _T_688; // @[Mux.scala 31:69:@19406.4]
  assign _T_690 = _T_678 ? _T_684 : _T_689; // @[Mux.scala 31:69:@19407.4]
  assign _T_691 = _T_677 ? _T_682 : _T_690; // @[Mux.scala 31:69:@19408.4]
  assign _T_696 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19415.4]
  assign _T_699 = _T_696 & _T_442; // @[MemPrimitives.scala 110:228:@19417.4]
  assign _T_702 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19419.4]
  assign _T_705 = _T_702 & _T_448; // @[MemPrimitives.scala 110:228:@19421.4]
  assign _T_707 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@19428.4]
  assign _T_708 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@19429.4]
  assign _T_710 = {_T_707,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19431.4]
  assign _T_712 = {_T_708,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19433.4]
  assign _T_713 = _T_707 ? _T_710 : _T_712; // @[Mux.scala 31:69:@19434.4]
  assign _T_718 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19441.4]
  assign _T_721 = _T_718 & _T_464; // @[MemPrimitives.scala 110:228:@19443.4]
  assign _T_724 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19445.4]
  assign _T_727 = _T_724 & _T_470; // @[MemPrimitives.scala 110:228:@19447.4]
  assign _T_730 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19449.4]
  assign _T_733 = _T_730 & _T_476; // @[MemPrimitives.scala 110:228:@19451.4]
  assign _T_736 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19453.4]
  assign _T_739 = _T_736 & _T_482; // @[MemPrimitives.scala 110:228:@19455.4]
  assign _T_741 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@19464.4]
  assign _T_742 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@19465.4]
  assign _T_743 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@19466.4]
  assign _T_744 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@19467.4]
  assign _T_746 = {_T_741,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19469.4]
  assign _T_748 = {_T_742,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19471.4]
  assign _T_750 = {_T_743,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19473.4]
  assign _T_752 = {_T_744,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19475.4]
  assign _T_753 = _T_743 ? _T_750 : _T_752; // @[Mux.scala 31:69:@19476.4]
  assign _T_754 = _T_742 ? _T_748 : _T_753; // @[Mux.scala 31:69:@19477.4]
  assign _T_755 = _T_741 ? _T_746 : _T_754; // @[Mux.scala 31:69:@19478.4]
  assign _T_763 = _T_696 & _T_506; // @[MemPrimitives.scala 110:228:@19487.4]
  assign _T_769 = _T_702 & _T_512; // @[MemPrimitives.scala 110:228:@19491.4]
  assign _T_771 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@19498.4]
  assign _T_772 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@19499.4]
  assign _T_774 = {_T_771,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19501.4]
  assign _T_776 = {_T_772,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19503.4]
  assign _T_777 = _T_771 ? _T_774 : _T_776; // @[Mux.scala 31:69:@19504.4]
  assign _T_785 = _T_718 & _T_528; // @[MemPrimitives.scala 110:228:@19513.4]
  assign _T_791 = _T_724 & _T_534; // @[MemPrimitives.scala 110:228:@19517.4]
  assign _T_797 = _T_730 & _T_540; // @[MemPrimitives.scala 110:228:@19521.4]
  assign _T_803 = _T_736 & _T_546; // @[MemPrimitives.scala 110:228:@19525.4]
  assign _T_805 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@19534.4]
  assign _T_806 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@19535.4]
  assign _T_807 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@19536.4]
  assign _T_808 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@19537.4]
  assign _T_810 = {_T_805,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19539.4]
  assign _T_812 = {_T_806,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19541.4]
  assign _T_814 = {_T_807,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19543.4]
  assign _T_816 = {_T_808,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19545.4]
  assign _T_817 = _T_807 ? _T_814 : _T_816; // @[Mux.scala 31:69:@19546.4]
  assign _T_818 = _T_806 ? _T_812 : _T_817; // @[Mux.scala 31:69:@19547.4]
  assign _T_819 = _T_805 ? _T_810 : _T_818; // @[Mux.scala 31:69:@19548.4]
  assign _T_824 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19555.4]
  assign _T_827 = _T_824 & _T_442; // @[MemPrimitives.scala 110:228:@19557.4]
  assign _T_830 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19559.4]
  assign _T_833 = _T_830 & _T_448; // @[MemPrimitives.scala 110:228:@19561.4]
  assign _T_835 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@19568.4]
  assign _T_836 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@19569.4]
  assign _T_838 = {_T_835,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19571.4]
  assign _T_840 = {_T_836,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19573.4]
  assign _T_841 = _T_835 ? _T_838 : _T_840; // @[Mux.scala 31:69:@19574.4]
  assign _T_846 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19581.4]
  assign _T_849 = _T_846 & _T_464; // @[MemPrimitives.scala 110:228:@19583.4]
  assign _T_852 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19585.4]
  assign _T_855 = _T_852 & _T_470; // @[MemPrimitives.scala 110:228:@19587.4]
  assign _T_858 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19589.4]
  assign _T_861 = _T_858 & _T_476; // @[MemPrimitives.scala 110:228:@19591.4]
  assign _T_864 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19593.4]
  assign _T_867 = _T_864 & _T_482; // @[MemPrimitives.scala 110:228:@19595.4]
  assign _T_869 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@19604.4]
  assign _T_870 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@19605.4]
  assign _T_871 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@19606.4]
  assign _T_872 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@19607.4]
  assign _T_874 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19609.4]
  assign _T_876 = {_T_870,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19611.4]
  assign _T_878 = {_T_871,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19613.4]
  assign _T_880 = {_T_872,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19615.4]
  assign _T_881 = _T_871 ? _T_878 : _T_880; // @[Mux.scala 31:69:@19616.4]
  assign _T_882 = _T_870 ? _T_876 : _T_881; // @[Mux.scala 31:69:@19617.4]
  assign _T_883 = _T_869 ? _T_874 : _T_882; // @[Mux.scala 31:69:@19618.4]
  assign _T_891 = _T_824 & _T_506; // @[MemPrimitives.scala 110:228:@19627.4]
  assign _T_897 = _T_830 & _T_512; // @[MemPrimitives.scala 110:228:@19631.4]
  assign _T_899 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@19638.4]
  assign _T_900 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@19639.4]
  assign _T_902 = {_T_899,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19641.4]
  assign _T_904 = {_T_900,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19643.4]
  assign _T_905 = _T_899 ? _T_902 : _T_904; // @[Mux.scala 31:69:@19644.4]
  assign _T_913 = _T_846 & _T_528; // @[MemPrimitives.scala 110:228:@19653.4]
  assign _T_919 = _T_852 & _T_534; // @[MemPrimitives.scala 110:228:@19657.4]
  assign _T_925 = _T_858 & _T_540; // @[MemPrimitives.scala 110:228:@19661.4]
  assign _T_931 = _T_864 & _T_546; // @[MemPrimitives.scala 110:228:@19665.4]
  assign _T_933 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@19674.4]
  assign _T_934 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@19675.4]
  assign _T_935 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@19676.4]
  assign _T_936 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@19677.4]
  assign _T_938 = {_T_933,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19679.4]
  assign _T_940 = {_T_934,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19681.4]
  assign _T_942 = {_T_935,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19683.4]
  assign _T_944 = {_T_936,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19685.4]
  assign _T_945 = _T_935 ? _T_942 : _T_944; // @[Mux.scala 31:69:@19686.4]
  assign _T_946 = _T_934 ? _T_940 : _T_945; // @[Mux.scala 31:69:@19687.4]
  assign _T_947 = _T_933 ? _T_938 : _T_946; // @[Mux.scala 31:69:@19688.4]
  assign _T_1011 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@19773.4 package.scala 96:25:@19774.4]
  assign _T_1015 = _T_1011 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@19783.4]
  assign _T_1008 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@19765.4 package.scala 96:25:@19766.4]
  assign _T_1016 = _T_1008 ? Mem1D_11_io_output : _T_1015; // @[Mux.scala 31:69:@19784.4]
  assign _T_1005 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@19757.4 package.scala 96:25:@19758.4]
  assign _T_1017 = _T_1005 ? Mem1D_9_io_output : _T_1016; // @[Mux.scala 31:69:@19785.4]
  assign _T_1002 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@19749.4 package.scala 96:25:@19750.4]
  assign _T_1018 = _T_1002 ? Mem1D_7_io_output : _T_1017; // @[Mux.scala 31:69:@19786.4]
  assign _T_999 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@19741.4 package.scala 96:25:@19742.4]
  assign _T_1019 = _T_999 ? Mem1D_5_io_output : _T_1018; // @[Mux.scala 31:69:@19787.4]
  assign _T_996 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@19733.4 package.scala 96:25:@19734.4]
  assign _T_1020 = _T_996 ? Mem1D_3_io_output : _T_1019; // @[Mux.scala 31:69:@19788.4]
  assign _T_993 = RetimeWrapper_io_out; // @[package.scala 96:25:@19725.4 package.scala 96:25:@19726.4]
  assign _T_1082 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@19869.4 package.scala 96:25:@19870.4]
  assign _T_1086 = _T_1082 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@19879.4]
  assign _T_1079 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@19861.4 package.scala 96:25:@19862.4]
  assign _T_1087 = _T_1079 ? Mem1D_10_io_output : _T_1086; // @[Mux.scala 31:69:@19880.4]
  assign _T_1076 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@19853.4 package.scala 96:25:@19854.4]
  assign _T_1088 = _T_1076 ? Mem1D_8_io_output : _T_1087; // @[Mux.scala 31:69:@19881.4]
  assign _T_1073 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@19845.4 package.scala 96:25:@19846.4]
  assign _T_1089 = _T_1073 ? Mem1D_6_io_output : _T_1088; // @[Mux.scala 31:69:@19882.4]
  assign _T_1070 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@19837.4 package.scala 96:25:@19838.4]
  assign _T_1090 = _T_1070 ? Mem1D_4_io_output : _T_1089; // @[Mux.scala 31:69:@19883.4]
  assign _T_1067 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@19829.4 package.scala 96:25:@19830.4]
  assign _T_1091 = _T_1067 ? Mem1D_2_io_output : _T_1090; // @[Mux.scala 31:69:@19884.4]
  assign _T_1064 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@19821.4 package.scala 96:25:@19822.4]
  assign _T_1153 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@19965.4 package.scala 96:25:@19966.4]
  assign _T_1157 = _T_1153 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@19975.4]
  assign _T_1150 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@19957.4 package.scala 96:25:@19958.4]
  assign _T_1158 = _T_1150 ? Mem1D_10_io_output : _T_1157; // @[Mux.scala 31:69:@19976.4]
  assign _T_1147 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@19949.4 package.scala 96:25:@19950.4]
  assign _T_1159 = _T_1147 ? Mem1D_8_io_output : _T_1158; // @[Mux.scala 31:69:@19977.4]
  assign _T_1144 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@19941.4 package.scala 96:25:@19942.4]
  assign _T_1160 = _T_1144 ? Mem1D_6_io_output : _T_1159; // @[Mux.scala 31:69:@19978.4]
  assign _T_1141 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@19933.4 package.scala 96:25:@19934.4]
  assign _T_1161 = _T_1141 ? Mem1D_4_io_output : _T_1160; // @[Mux.scala 31:69:@19979.4]
  assign _T_1138 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@19925.4 package.scala 96:25:@19926.4]
  assign _T_1162 = _T_1138 ? Mem1D_2_io_output : _T_1161; // @[Mux.scala 31:69:@19980.4]
  assign _T_1135 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@19917.4 package.scala 96:25:@19918.4]
  assign _T_1224 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@20061.4 package.scala 96:25:@20062.4]
  assign _T_1228 = _T_1224 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@20071.4]
  assign _T_1221 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@20053.4 package.scala 96:25:@20054.4]
  assign _T_1229 = _T_1221 ? Mem1D_11_io_output : _T_1228; // @[Mux.scala 31:69:@20072.4]
  assign _T_1218 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@20045.4 package.scala 96:25:@20046.4]
  assign _T_1230 = _T_1218 ? Mem1D_9_io_output : _T_1229; // @[Mux.scala 31:69:@20073.4]
  assign _T_1215 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@20037.4 package.scala 96:25:@20038.4]
  assign _T_1231 = _T_1215 ? Mem1D_7_io_output : _T_1230; // @[Mux.scala 31:69:@20074.4]
  assign _T_1212 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@20029.4 package.scala 96:25:@20030.4]
  assign _T_1232 = _T_1212 ? Mem1D_5_io_output : _T_1231; // @[Mux.scala 31:69:@20075.4]
  assign _T_1209 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@20021.4 package.scala 96:25:@20022.4]
  assign _T_1233 = _T_1209 ? Mem1D_3_io_output : _T_1232; // @[Mux.scala 31:69:@20076.4]
  assign _T_1206 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@20013.4 package.scala 96:25:@20014.4]
  assign _T_1295 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@20157.4 package.scala 96:25:@20158.4]
  assign _T_1299 = _T_1295 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@20167.4]
  assign _T_1292 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@20149.4 package.scala 96:25:@20150.4]
  assign _T_1300 = _T_1292 ? Mem1D_11_io_output : _T_1299; // @[Mux.scala 31:69:@20168.4]
  assign _T_1289 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@20141.4 package.scala 96:25:@20142.4]
  assign _T_1301 = _T_1289 ? Mem1D_9_io_output : _T_1300; // @[Mux.scala 31:69:@20169.4]
  assign _T_1286 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@20133.4 package.scala 96:25:@20134.4]
  assign _T_1302 = _T_1286 ? Mem1D_7_io_output : _T_1301; // @[Mux.scala 31:69:@20170.4]
  assign _T_1283 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@20125.4 package.scala 96:25:@20126.4]
  assign _T_1303 = _T_1283 ? Mem1D_5_io_output : _T_1302; // @[Mux.scala 31:69:@20171.4]
  assign _T_1280 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@20117.4 package.scala 96:25:@20118.4]
  assign _T_1304 = _T_1280 ? Mem1D_3_io_output : _T_1303; // @[Mux.scala 31:69:@20172.4]
  assign _T_1277 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@20109.4 package.scala 96:25:@20110.4]
  assign _T_1366 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@20253.4 package.scala 96:25:@20254.4]
  assign _T_1370 = _T_1366 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@20263.4]
  assign _T_1363 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@20245.4 package.scala 96:25:@20246.4]
  assign _T_1371 = _T_1363 ? Mem1D_11_io_output : _T_1370; // @[Mux.scala 31:69:@20264.4]
  assign _T_1360 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@20237.4 package.scala 96:25:@20238.4]
  assign _T_1372 = _T_1360 ? Mem1D_9_io_output : _T_1371; // @[Mux.scala 31:69:@20265.4]
  assign _T_1357 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@20229.4 package.scala 96:25:@20230.4]
  assign _T_1373 = _T_1357 ? Mem1D_7_io_output : _T_1372; // @[Mux.scala 31:69:@20266.4]
  assign _T_1354 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@20221.4 package.scala 96:25:@20222.4]
  assign _T_1374 = _T_1354 ? Mem1D_5_io_output : _T_1373; // @[Mux.scala 31:69:@20267.4]
  assign _T_1351 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@20213.4 package.scala 96:25:@20214.4]
  assign _T_1375 = _T_1351 ? Mem1D_3_io_output : _T_1374; // @[Mux.scala 31:69:@20268.4]
  assign _T_1348 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@20205.4 package.scala 96:25:@20206.4]
  assign io_rPort_5_output_0 = _T_1348 ? Mem1D_1_io_output : _T_1375; // @[MemPrimitives.scala 152:13:@20270.4]
  assign io_rPort_4_output_0 = _T_1277 ? Mem1D_1_io_output : _T_1304; // @[MemPrimitives.scala 152:13:@20174.4]
  assign io_rPort_3_output_0 = _T_1206 ? Mem1D_1_io_output : _T_1233; // @[MemPrimitives.scala 152:13:@20078.4]
  assign io_rPort_2_output_0 = _T_1135 ? Mem1D_io_output : _T_1162; // @[MemPrimitives.scala 152:13:@19982.4]
  assign io_rPort_1_output_0 = _T_1064 ? Mem1D_io_output : _T_1091; // @[MemPrimitives.scala 152:13:@19886.4]
  assign io_rPort_0_output_0 = _T_993 ? Mem1D_1_io_output : _T_1020; // @[MemPrimitives.scala 152:13:@19790.4]
  assign Mem1D_clock = clock; // @[:@18688.4]
  assign Mem1D_reset = reset; // @[:@18689.4]
  assign Mem1D_io_r_ofs_0 = _T_457[8:0]; // @[MemPrimitives.scala 131:28:@19158.4]
  assign Mem1D_io_r_backpressure = _T_457[9]; // @[MemPrimitives.scala 132:32:@19159.4]
  assign Mem1D_io_w_ofs_0 = _T_270[8:0]; // @[MemPrimitives.scala 94:28:@18952.4]
  assign Mem1D_io_w_data_0 = _T_270[40:9]; // @[MemPrimitives.scala 95:29:@18953.4]
  assign Mem1D_io_w_en_0 = _T_270[41]; // @[MemPrimitives.scala 96:27:@18954.4]
  assign Mem1D_1_clock = clock; // @[:@18704.4]
  assign Mem1D_1_reset = reset; // @[:@18705.4]
  assign Mem1D_1_io_r_ofs_0 = _T_499[8:0]; // @[MemPrimitives.scala 131:28:@19202.4]
  assign Mem1D_1_io_r_backpressure = _T_499[9]; // @[MemPrimitives.scala 132:32:@19203.4]
  assign Mem1D_1_io_w_ofs_0 = _T_281[8:0]; // @[MemPrimitives.scala 94:28:@18964.4]
  assign Mem1D_1_io_w_data_0 = _T_281[40:9]; // @[MemPrimitives.scala 95:29:@18965.4]
  assign Mem1D_1_io_w_en_0 = _T_281[41]; // @[MemPrimitives.scala 96:27:@18966.4]
  assign Mem1D_2_clock = clock; // @[:@18720.4]
  assign Mem1D_2_reset = reset; // @[:@18721.4]
  assign Mem1D_2_io_r_ofs_0 = _T_521[8:0]; // @[MemPrimitives.scala 131:28:@19228.4]
  assign Mem1D_2_io_r_backpressure = _T_521[9]; // @[MemPrimitives.scala 132:32:@19229.4]
  assign Mem1D_2_io_w_ofs_0 = _T_292[8:0]; // @[MemPrimitives.scala 94:28:@18976.4]
  assign Mem1D_2_io_w_data_0 = _T_292[40:9]; // @[MemPrimitives.scala 95:29:@18977.4]
  assign Mem1D_2_io_w_en_0 = _T_292[41]; // @[MemPrimitives.scala 96:27:@18978.4]
  assign Mem1D_3_clock = clock; // @[:@18736.4]
  assign Mem1D_3_reset = reset; // @[:@18737.4]
  assign Mem1D_3_io_r_ofs_0 = _T_563[8:0]; // @[MemPrimitives.scala 131:28:@19272.4]
  assign Mem1D_3_io_r_backpressure = _T_563[9]; // @[MemPrimitives.scala 132:32:@19273.4]
  assign Mem1D_3_io_w_ofs_0 = _T_303[8:0]; // @[MemPrimitives.scala 94:28:@18988.4]
  assign Mem1D_3_io_w_data_0 = _T_303[40:9]; // @[MemPrimitives.scala 95:29:@18989.4]
  assign Mem1D_3_io_w_en_0 = _T_303[41]; // @[MemPrimitives.scala 96:27:@18990.4]
  assign Mem1D_4_clock = clock; // @[:@18752.4]
  assign Mem1D_4_reset = reset; // @[:@18753.4]
  assign Mem1D_4_io_r_ofs_0 = _T_585[8:0]; // @[MemPrimitives.scala 131:28:@19298.4]
  assign Mem1D_4_io_r_backpressure = _T_585[9]; // @[MemPrimitives.scala 132:32:@19299.4]
  assign Mem1D_4_io_w_ofs_0 = _T_314[8:0]; // @[MemPrimitives.scala 94:28:@19000.4]
  assign Mem1D_4_io_w_data_0 = _T_314[40:9]; // @[MemPrimitives.scala 95:29:@19001.4]
  assign Mem1D_4_io_w_en_0 = _T_314[41]; // @[MemPrimitives.scala 96:27:@19002.4]
  assign Mem1D_5_clock = clock; // @[:@18768.4]
  assign Mem1D_5_reset = reset; // @[:@18769.4]
  assign Mem1D_5_io_r_ofs_0 = _T_627[8:0]; // @[MemPrimitives.scala 131:28:@19342.4]
  assign Mem1D_5_io_r_backpressure = _T_627[9]; // @[MemPrimitives.scala 132:32:@19343.4]
  assign Mem1D_5_io_w_ofs_0 = _T_325[8:0]; // @[MemPrimitives.scala 94:28:@19012.4]
  assign Mem1D_5_io_w_data_0 = _T_325[40:9]; // @[MemPrimitives.scala 95:29:@19013.4]
  assign Mem1D_5_io_w_en_0 = _T_325[41]; // @[MemPrimitives.scala 96:27:@19014.4]
  assign Mem1D_6_clock = clock; // @[:@18784.4]
  assign Mem1D_6_reset = reset; // @[:@18785.4]
  assign Mem1D_6_io_r_ofs_0 = _T_649[8:0]; // @[MemPrimitives.scala 131:28:@19368.4]
  assign Mem1D_6_io_r_backpressure = _T_649[9]; // @[MemPrimitives.scala 132:32:@19369.4]
  assign Mem1D_6_io_w_ofs_0 = _T_336[8:0]; // @[MemPrimitives.scala 94:28:@19024.4]
  assign Mem1D_6_io_w_data_0 = _T_336[40:9]; // @[MemPrimitives.scala 95:29:@19025.4]
  assign Mem1D_6_io_w_en_0 = _T_336[41]; // @[MemPrimitives.scala 96:27:@19026.4]
  assign Mem1D_7_clock = clock; // @[:@18800.4]
  assign Mem1D_7_reset = reset; // @[:@18801.4]
  assign Mem1D_7_io_r_ofs_0 = _T_691[8:0]; // @[MemPrimitives.scala 131:28:@19412.4]
  assign Mem1D_7_io_r_backpressure = _T_691[9]; // @[MemPrimitives.scala 132:32:@19413.4]
  assign Mem1D_7_io_w_ofs_0 = _T_347[8:0]; // @[MemPrimitives.scala 94:28:@19036.4]
  assign Mem1D_7_io_w_data_0 = _T_347[40:9]; // @[MemPrimitives.scala 95:29:@19037.4]
  assign Mem1D_7_io_w_en_0 = _T_347[41]; // @[MemPrimitives.scala 96:27:@19038.4]
  assign Mem1D_8_clock = clock; // @[:@18816.4]
  assign Mem1D_8_reset = reset; // @[:@18817.4]
  assign Mem1D_8_io_r_ofs_0 = _T_713[8:0]; // @[MemPrimitives.scala 131:28:@19438.4]
  assign Mem1D_8_io_r_backpressure = _T_713[9]; // @[MemPrimitives.scala 132:32:@19439.4]
  assign Mem1D_8_io_w_ofs_0 = _T_358[8:0]; // @[MemPrimitives.scala 94:28:@19048.4]
  assign Mem1D_8_io_w_data_0 = _T_358[40:9]; // @[MemPrimitives.scala 95:29:@19049.4]
  assign Mem1D_8_io_w_en_0 = _T_358[41]; // @[MemPrimitives.scala 96:27:@19050.4]
  assign Mem1D_9_clock = clock; // @[:@18832.4]
  assign Mem1D_9_reset = reset; // @[:@18833.4]
  assign Mem1D_9_io_r_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 131:28:@19482.4]
  assign Mem1D_9_io_r_backpressure = _T_755[9]; // @[MemPrimitives.scala 132:32:@19483.4]
  assign Mem1D_9_io_w_ofs_0 = _T_369[8:0]; // @[MemPrimitives.scala 94:28:@19060.4]
  assign Mem1D_9_io_w_data_0 = _T_369[40:9]; // @[MemPrimitives.scala 95:29:@19061.4]
  assign Mem1D_9_io_w_en_0 = _T_369[41]; // @[MemPrimitives.scala 96:27:@19062.4]
  assign Mem1D_10_clock = clock; // @[:@18848.4]
  assign Mem1D_10_reset = reset; // @[:@18849.4]
  assign Mem1D_10_io_r_ofs_0 = _T_777[8:0]; // @[MemPrimitives.scala 131:28:@19508.4]
  assign Mem1D_10_io_r_backpressure = _T_777[9]; // @[MemPrimitives.scala 132:32:@19509.4]
  assign Mem1D_10_io_w_ofs_0 = _T_380[8:0]; // @[MemPrimitives.scala 94:28:@19072.4]
  assign Mem1D_10_io_w_data_0 = _T_380[40:9]; // @[MemPrimitives.scala 95:29:@19073.4]
  assign Mem1D_10_io_w_en_0 = _T_380[41]; // @[MemPrimitives.scala 96:27:@19074.4]
  assign Mem1D_11_clock = clock; // @[:@18864.4]
  assign Mem1D_11_reset = reset; // @[:@18865.4]
  assign Mem1D_11_io_r_ofs_0 = _T_819[8:0]; // @[MemPrimitives.scala 131:28:@19552.4]
  assign Mem1D_11_io_r_backpressure = _T_819[9]; // @[MemPrimitives.scala 132:32:@19553.4]
  assign Mem1D_11_io_w_ofs_0 = _T_391[8:0]; // @[MemPrimitives.scala 94:28:@19084.4]
  assign Mem1D_11_io_w_data_0 = _T_391[40:9]; // @[MemPrimitives.scala 95:29:@19085.4]
  assign Mem1D_11_io_w_en_0 = _T_391[41]; // @[MemPrimitives.scala 96:27:@19086.4]
  assign Mem1D_12_clock = clock; // @[:@18880.4]
  assign Mem1D_12_reset = reset; // @[:@18881.4]
  assign Mem1D_12_io_r_ofs_0 = _T_841[8:0]; // @[MemPrimitives.scala 131:28:@19578.4]
  assign Mem1D_12_io_r_backpressure = _T_841[9]; // @[MemPrimitives.scala 132:32:@19579.4]
  assign Mem1D_12_io_w_ofs_0 = _T_402[8:0]; // @[MemPrimitives.scala 94:28:@19096.4]
  assign Mem1D_12_io_w_data_0 = _T_402[40:9]; // @[MemPrimitives.scala 95:29:@19097.4]
  assign Mem1D_12_io_w_en_0 = _T_402[41]; // @[MemPrimitives.scala 96:27:@19098.4]
  assign Mem1D_13_clock = clock; // @[:@18896.4]
  assign Mem1D_13_reset = reset; // @[:@18897.4]
  assign Mem1D_13_io_r_ofs_0 = _T_883[8:0]; // @[MemPrimitives.scala 131:28:@19622.4]
  assign Mem1D_13_io_r_backpressure = _T_883[9]; // @[MemPrimitives.scala 132:32:@19623.4]
  assign Mem1D_13_io_w_ofs_0 = _T_413[8:0]; // @[MemPrimitives.scala 94:28:@19108.4]
  assign Mem1D_13_io_w_data_0 = _T_413[40:9]; // @[MemPrimitives.scala 95:29:@19109.4]
  assign Mem1D_13_io_w_en_0 = _T_413[41]; // @[MemPrimitives.scala 96:27:@19110.4]
  assign Mem1D_14_clock = clock; // @[:@18912.4]
  assign Mem1D_14_reset = reset; // @[:@18913.4]
  assign Mem1D_14_io_r_ofs_0 = _T_905[8:0]; // @[MemPrimitives.scala 131:28:@19648.4]
  assign Mem1D_14_io_r_backpressure = _T_905[9]; // @[MemPrimitives.scala 132:32:@19649.4]
  assign Mem1D_14_io_w_ofs_0 = _T_424[8:0]; // @[MemPrimitives.scala 94:28:@19120.4]
  assign Mem1D_14_io_w_data_0 = _T_424[40:9]; // @[MemPrimitives.scala 95:29:@19121.4]
  assign Mem1D_14_io_w_en_0 = _T_424[41]; // @[MemPrimitives.scala 96:27:@19122.4]
  assign Mem1D_15_clock = clock; // @[:@18928.4]
  assign Mem1D_15_reset = reset; // @[:@18929.4]
  assign Mem1D_15_io_r_ofs_0 = _T_947[8:0]; // @[MemPrimitives.scala 131:28:@19692.4]
  assign Mem1D_15_io_r_backpressure = _T_947[9]; // @[MemPrimitives.scala 132:32:@19693.4]
  assign Mem1D_15_io_w_ofs_0 = _T_435[8:0]; // @[MemPrimitives.scala 94:28:@19132.4]
  assign Mem1D_15_io_w_data_0 = _T_435[40:9]; // @[MemPrimitives.scala 95:29:@19133.4]
  assign Mem1D_15_io_w_en_0 = _T_435[41]; // @[MemPrimitives.scala 96:27:@19134.4]
  assign StickySelects_clock = clock; // @[:@19144.4]
  assign StickySelects_reset = reset; // @[:@19145.4]
  assign StickySelects_io_ins_0 = io_rPort_1_en_0 & _T_443; // @[MemPrimitives.scala 125:64:@19146.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_449; // @[MemPrimitives.scala 125:64:@19147.4]
  assign StickySelects_1_clock = clock; // @[:@19178.4]
  assign StickySelects_1_reset = reset; // @[:@19179.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_465; // @[MemPrimitives.scala 125:64:@19180.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_471; // @[MemPrimitives.scala 125:64:@19181.4]
  assign StickySelects_1_io_ins_2 = io_rPort_4_en_0 & _T_477; // @[MemPrimitives.scala 125:64:@19182.4]
  assign StickySelects_1_io_ins_3 = io_rPort_5_en_0 & _T_483; // @[MemPrimitives.scala 125:64:@19183.4]
  assign StickySelects_2_clock = clock; // @[:@19214.4]
  assign StickySelects_2_reset = reset; // @[:@19215.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_507; // @[MemPrimitives.scala 125:64:@19216.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_513; // @[MemPrimitives.scala 125:64:@19217.4]
  assign StickySelects_3_clock = clock; // @[:@19248.4]
  assign StickySelects_3_reset = reset; // @[:@19249.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_529; // @[MemPrimitives.scala 125:64:@19250.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_535; // @[MemPrimitives.scala 125:64:@19251.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_541; // @[MemPrimitives.scala 125:64:@19252.4]
  assign StickySelects_3_io_ins_3 = io_rPort_5_en_0 & _T_547; // @[MemPrimitives.scala 125:64:@19253.4]
  assign StickySelects_4_clock = clock; // @[:@19284.4]
  assign StickySelects_4_reset = reset; // @[:@19285.4]
  assign StickySelects_4_io_ins_0 = io_rPort_1_en_0 & _T_571; // @[MemPrimitives.scala 125:64:@19286.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_577; // @[MemPrimitives.scala 125:64:@19287.4]
  assign StickySelects_5_clock = clock; // @[:@19318.4]
  assign StickySelects_5_reset = reset; // @[:@19319.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_593; // @[MemPrimitives.scala 125:64:@19320.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_599; // @[MemPrimitives.scala 125:64:@19321.4]
  assign StickySelects_5_io_ins_2 = io_rPort_4_en_0 & _T_605; // @[MemPrimitives.scala 125:64:@19322.4]
  assign StickySelects_5_io_ins_3 = io_rPort_5_en_0 & _T_611; // @[MemPrimitives.scala 125:64:@19323.4]
  assign StickySelects_6_clock = clock; // @[:@19354.4]
  assign StickySelects_6_reset = reset; // @[:@19355.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@19356.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@19357.4]
  assign StickySelects_7_clock = clock; // @[:@19388.4]
  assign StickySelects_7_reset = reset; // @[:@19389.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_657; // @[MemPrimitives.scala 125:64:@19390.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_663; // @[MemPrimitives.scala 125:64:@19391.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_669; // @[MemPrimitives.scala 125:64:@19392.4]
  assign StickySelects_7_io_ins_3 = io_rPort_5_en_0 & _T_675; // @[MemPrimitives.scala 125:64:@19393.4]
  assign StickySelects_8_clock = clock; // @[:@19424.4]
  assign StickySelects_8_reset = reset; // @[:@19425.4]
  assign StickySelects_8_io_ins_0 = io_rPort_1_en_0 & _T_699; // @[MemPrimitives.scala 125:64:@19426.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_705; // @[MemPrimitives.scala 125:64:@19427.4]
  assign StickySelects_9_clock = clock; // @[:@19458.4]
  assign StickySelects_9_reset = reset; // @[:@19459.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_721; // @[MemPrimitives.scala 125:64:@19460.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@19461.4]
  assign StickySelects_9_io_ins_2 = io_rPort_4_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@19462.4]
  assign StickySelects_9_io_ins_3 = io_rPort_5_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@19463.4]
  assign StickySelects_10_clock = clock; // @[:@19494.4]
  assign StickySelects_10_reset = reset; // @[:@19495.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@19496.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@19497.4]
  assign StickySelects_11_clock = clock; // @[:@19528.4]
  assign StickySelects_11_reset = reset; // @[:@19529.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_785; // @[MemPrimitives.scala 125:64:@19530.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_791; // @[MemPrimitives.scala 125:64:@19531.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_797; // @[MemPrimitives.scala 125:64:@19532.4]
  assign StickySelects_11_io_ins_3 = io_rPort_5_en_0 & _T_803; // @[MemPrimitives.scala 125:64:@19533.4]
  assign StickySelects_12_clock = clock; // @[:@19564.4]
  assign StickySelects_12_reset = reset; // @[:@19565.4]
  assign StickySelects_12_io_ins_0 = io_rPort_1_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@19566.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@19567.4]
  assign StickySelects_13_clock = clock; // @[:@19598.4]
  assign StickySelects_13_reset = reset; // @[:@19599.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_849; // @[MemPrimitives.scala 125:64:@19600.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_855; // @[MemPrimitives.scala 125:64:@19601.4]
  assign StickySelects_13_io_ins_2 = io_rPort_4_en_0 & _T_861; // @[MemPrimitives.scala 125:64:@19602.4]
  assign StickySelects_13_io_ins_3 = io_rPort_5_en_0 & _T_867; // @[MemPrimitives.scala 125:64:@19603.4]
  assign StickySelects_14_clock = clock; // @[:@19634.4]
  assign StickySelects_14_reset = reset; // @[:@19635.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_891; // @[MemPrimitives.scala 125:64:@19636.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_897; // @[MemPrimitives.scala 125:64:@19637.4]
  assign StickySelects_15_clock = clock; // @[:@19668.4]
  assign StickySelects_15_reset = reset; // @[:@19669.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_913; // @[MemPrimitives.scala 125:64:@19670.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_919; // @[MemPrimitives.scala 125:64:@19671.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_925; // @[MemPrimitives.scala 125:64:@19672.4]
  assign StickySelects_15_io_ins_3 = io_rPort_5_en_0 & _T_931; // @[MemPrimitives.scala 125:64:@19673.4]
  assign RetimeWrapper_clock = clock; // @[:@19721.4]
  assign RetimeWrapper_reset = reset; // @[:@19722.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19724.4]
  assign RetimeWrapper_io_in = _T_465 & io_rPort_0_en_0; // @[package.scala 94:16:@19723.4]
  assign RetimeWrapper_1_clock = clock; // @[:@19729.4]
  assign RetimeWrapper_1_reset = reset; // @[:@19730.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19732.4]
  assign RetimeWrapper_1_io_in = _T_529 & io_rPort_0_en_0; // @[package.scala 94:16:@19731.4]
  assign RetimeWrapper_2_clock = clock; // @[:@19737.4]
  assign RetimeWrapper_2_reset = reset; // @[:@19738.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19740.4]
  assign RetimeWrapper_2_io_in = _T_593 & io_rPort_0_en_0; // @[package.scala 94:16:@19739.4]
  assign RetimeWrapper_3_clock = clock; // @[:@19745.4]
  assign RetimeWrapper_3_reset = reset; // @[:@19746.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19748.4]
  assign RetimeWrapper_3_io_in = _T_657 & io_rPort_0_en_0; // @[package.scala 94:16:@19747.4]
  assign RetimeWrapper_4_clock = clock; // @[:@19753.4]
  assign RetimeWrapper_4_reset = reset; // @[:@19754.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19756.4]
  assign RetimeWrapper_4_io_in = _T_721 & io_rPort_0_en_0; // @[package.scala 94:16:@19755.4]
  assign RetimeWrapper_5_clock = clock; // @[:@19761.4]
  assign RetimeWrapper_5_reset = reset; // @[:@19762.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19764.4]
  assign RetimeWrapper_5_io_in = _T_785 & io_rPort_0_en_0; // @[package.scala 94:16:@19763.4]
  assign RetimeWrapper_6_clock = clock; // @[:@19769.4]
  assign RetimeWrapper_6_reset = reset; // @[:@19770.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19772.4]
  assign RetimeWrapper_6_io_in = _T_849 & io_rPort_0_en_0; // @[package.scala 94:16:@19771.4]
  assign RetimeWrapper_7_clock = clock; // @[:@19777.4]
  assign RetimeWrapper_7_reset = reset; // @[:@19778.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19780.4]
  assign RetimeWrapper_7_io_in = _T_913 & io_rPort_0_en_0; // @[package.scala 94:16:@19779.4]
  assign RetimeWrapper_8_clock = clock; // @[:@19817.4]
  assign RetimeWrapper_8_reset = reset; // @[:@19818.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19820.4]
  assign RetimeWrapper_8_io_in = _T_443 & io_rPort_1_en_0; // @[package.scala 94:16:@19819.4]
  assign RetimeWrapper_9_clock = clock; // @[:@19825.4]
  assign RetimeWrapper_9_reset = reset; // @[:@19826.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19828.4]
  assign RetimeWrapper_9_io_in = _T_507 & io_rPort_1_en_0; // @[package.scala 94:16:@19827.4]
  assign RetimeWrapper_10_clock = clock; // @[:@19833.4]
  assign RetimeWrapper_10_reset = reset; // @[:@19834.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19836.4]
  assign RetimeWrapper_10_io_in = _T_571 & io_rPort_1_en_0; // @[package.scala 94:16:@19835.4]
  assign RetimeWrapper_11_clock = clock; // @[:@19841.4]
  assign RetimeWrapper_11_reset = reset; // @[:@19842.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19844.4]
  assign RetimeWrapper_11_io_in = _T_635 & io_rPort_1_en_0; // @[package.scala 94:16:@19843.4]
  assign RetimeWrapper_12_clock = clock; // @[:@19849.4]
  assign RetimeWrapper_12_reset = reset; // @[:@19850.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19852.4]
  assign RetimeWrapper_12_io_in = _T_699 & io_rPort_1_en_0; // @[package.scala 94:16:@19851.4]
  assign RetimeWrapper_13_clock = clock; // @[:@19857.4]
  assign RetimeWrapper_13_reset = reset; // @[:@19858.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19860.4]
  assign RetimeWrapper_13_io_in = _T_763 & io_rPort_1_en_0; // @[package.scala 94:16:@19859.4]
  assign RetimeWrapper_14_clock = clock; // @[:@19865.4]
  assign RetimeWrapper_14_reset = reset; // @[:@19866.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19868.4]
  assign RetimeWrapper_14_io_in = _T_827 & io_rPort_1_en_0; // @[package.scala 94:16:@19867.4]
  assign RetimeWrapper_15_clock = clock; // @[:@19873.4]
  assign RetimeWrapper_15_reset = reset; // @[:@19874.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19876.4]
  assign RetimeWrapper_15_io_in = _T_891 & io_rPort_1_en_0; // @[package.scala 94:16:@19875.4]
  assign RetimeWrapper_16_clock = clock; // @[:@19913.4]
  assign RetimeWrapper_16_reset = reset; // @[:@19914.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19916.4]
  assign RetimeWrapper_16_io_in = _T_449 & io_rPort_2_en_0; // @[package.scala 94:16:@19915.4]
  assign RetimeWrapper_17_clock = clock; // @[:@19921.4]
  assign RetimeWrapper_17_reset = reset; // @[:@19922.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19924.4]
  assign RetimeWrapper_17_io_in = _T_513 & io_rPort_2_en_0; // @[package.scala 94:16:@19923.4]
  assign RetimeWrapper_18_clock = clock; // @[:@19929.4]
  assign RetimeWrapper_18_reset = reset; // @[:@19930.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19932.4]
  assign RetimeWrapper_18_io_in = _T_577 & io_rPort_2_en_0; // @[package.scala 94:16:@19931.4]
  assign RetimeWrapper_19_clock = clock; // @[:@19937.4]
  assign RetimeWrapper_19_reset = reset; // @[:@19938.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19940.4]
  assign RetimeWrapper_19_io_in = _T_641 & io_rPort_2_en_0; // @[package.scala 94:16:@19939.4]
  assign RetimeWrapper_20_clock = clock; // @[:@19945.4]
  assign RetimeWrapper_20_reset = reset; // @[:@19946.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19948.4]
  assign RetimeWrapper_20_io_in = _T_705 & io_rPort_2_en_0; // @[package.scala 94:16:@19947.4]
  assign RetimeWrapper_21_clock = clock; // @[:@19953.4]
  assign RetimeWrapper_21_reset = reset; // @[:@19954.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19956.4]
  assign RetimeWrapper_21_io_in = _T_769 & io_rPort_2_en_0; // @[package.scala 94:16:@19955.4]
  assign RetimeWrapper_22_clock = clock; // @[:@19961.4]
  assign RetimeWrapper_22_reset = reset; // @[:@19962.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19964.4]
  assign RetimeWrapper_22_io_in = _T_833 & io_rPort_2_en_0; // @[package.scala 94:16:@19963.4]
  assign RetimeWrapper_23_clock = clock; // @[:@19969.4]
  assign RetimeWrapper_23_reset = reset; // @[:@19970.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19972.4]
  assign RetimeWrapper_23_io_in = _T_897 & io_rPort_2_en_0; // @[package.scala 94:16:@19971.4]
  assign RetimeWrapper_24_clock = clock; // @[:@20009.4]
  assign RetimeWrapper_24_reset = reset; // @[:@20010.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20012.4]
  assign RetimeWrapper_24_io_in = _T_471 & io_rPort_3_en_0; // @[package.scala 94:16:@20011.4]
  assign RetimeWrapper_25_clock = clock; // @[:@20017.4]
  assign RetimeWrapper_25_reset = reset; // @[:@20018.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20020.4]
  assign RetimeWrapper_25_io_in = _T_535 & io_rPort_3_en_0; // @[package.scala 94:16:@20019.4]
  assign RetimeWrapper_26_clock = clock; // @[:@20025.4]
  assign RetimeWrapper_26_reset = reset; // @[:@20026.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20028.4]
  assign RetimeWrapper_26_io_in = _T_599 & io_rPort_3_en_0; // @[package.scala 94:16:@20027.4]
  assign RetimeWrapper_27_clock = clock; // @[:@20033.4]
  assign RetimeWrapper_27_reset = reset; // @[:@20034.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20036.4]
  assign RetimeWrapper_27_io_in = _T_663 & io_rPort_3_en_0; // @[package.scala 94:16:@20035.4]
  assign RetimeWrapper_28_clock = clock; // @[:@20041.4]
  assign RetimeWrapper_28_reset = reset; // @[:@20042.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20044.4]
  assign RetimeWrapper_28_io_in = _T_727 & io_rPort_3_en_0; // @[package.scala 94:16:@20043.4]
  assign RetimeWrapper_29_clock = clock; // @[:@20049.4]
  assign RetimeWrapper_29_reset = reset; // @[:@20050.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20052.4]
  assign RetimeWrapper_29_io_in = _T_791 & io_rPort_3_en_0; // @[package.scala 94:16:@20051.4]
  assign RetimeWrapper_30_clock = clock; // @[:@20057.4]
  assign RetimeWrapper_30_reset = reset; // @[:@20058.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20060.4]
  assign RetimeWrapper_30_io_in = _T_855 & io_rPort_3_en_0; // @[package.scala 94:16:@20059.4]
  assign RetimeWrapper_31_clock = clock; // @[:@20065.4]
  assign RetimeWrapper_31_reset = reset; // @[:@20066.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20068.4]
  assign RetimeWrapper_31_io_in = _T_919 & io_rPort_3_en_0; // @[package.scala 94:16:@20067.4]
  assign RetimeWrapper_32_clock = clock; // @[:@20105.4]
  assign RetimeWrapper_32_reset = reset; // @[:@20106.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20108.4]
  assign RetimeWrapper_32_io_in = _T_477 & io_rPort_4_en_0; // @[package.scala 94:16:@20107.4]
  assign RetimeWrapper_33_clock = clock; // @[:@20113.4]
  assign RetimeWrapper_33_reset = reset; // @[:@20114.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20116.4]
  assign RetimeWrapper_33_io_in = _T_541 & io_rPort_4_en_0; // @[package.scala 94:16:@20115.4]
  assign RetimeWrapper_34_clock = clock; // @[:@20121.4]
  assign RetimeWrapper_34_reset = reset; // @[:@20122.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20124.4]
  assign RetimeWrapper_34_io_in = _T_605 & io_rPort_4_en_0; // @[package.scala 94:16:@20123.4]
  assign RetimeWrapper_35_clock = clock; // @[:@20129.4]
  assign RetimeWrapper_35_reset = reset; // @[:@20130.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20132.4]
  assign RetimeWrapper_35_io_in = _T_669 & io_rPort_4_en_0; // @[package.scala 94:16:@20131.4]
  assign RetimeWrapper_36_clock = clock; // @[:@20137.4]
  assign RetimeWrapper_36_reset = reset; // @[:@20138.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20140.4]
  assign RetimeWrapper_36_io_in = _T_733 & io_rPort_4_en_0; // @[package.scala 94:16:@20139.4]
  assign RetimeWrapper_37_clock = clock; // @[:@20145.4]
  assign RetimeWrapper_37_reset = reset; // @[:@20146.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20148.4]
  assign RetimeWrapper_37_io_in = _T_797 & io_rPort_4_en_0; // @[package.scala 94:16:@20147.4]
  assign RetimeWrapper_38_clock = clock; // @[:@20153.4]
  assign RetimeWrapper_38_reset = reset; // @[:@20154.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20156.4]
  assign RetimeWrapper_38_io_in = _T_861 & io_rPort_4_en_0; // @[package.scala 94:16:@20155.4]
  assign RetimeWrapper_39_clock = clock; // @[:@20161.4]
  assign RetimeWrapper_39_reset = reset; // @[:@20162.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20164.4]
  assign RetimeWrapper_39_io_in = _T_925 & io_rPort_4_en_0; // @[package.scala 94:16:@20163.4]
  assign RetimeWrapper_40_clock = clock; // @[:@20201.4]
  assign RetimeWrapper_40_reset = reset; // @[:@20202.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20204.4]
  assign RetimeWrapper_40_io_in = _T_483 & io_rPort_5_en_0; // @[package.scala 94:16:@20203.4]
  assign RetimeWrapper_41_clock = clock; // @[:@20209.4]
  assign RetimeWrapper_41_reset = reset; // @[:@20210.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20212.4]
  assign RetimeWrapper_41_io_in = _T_547 & io_rPort_5_en_0; // @[package.scala 94:16:@20211.4]
  assign RetimeWrapper_42_clock = clock; // @[:@20217.4]
  assign RetimeWrapper_42_reset = reset; // @[:@20218.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20220.4]
  assign RetimeWrapper_42_io_in = _T_611 & io_rPort_5_en_0; // @[package.scala 94:16:@20219.4]
  assign RetimeWrapper_43_clock = clock; // @[:@20225.4]
  assign RetimeWrapper_43_reset = reset; // @[:@20226.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20228.4]
  assign RetimeWrapper_43_io_in = _T_675 & io_rPort_5_en_0; // @[package.scala 94:16:@20227.4]
  assign RetimeWrapper_44_clock = clock; // @[:@20233.4]
  assign RetimeWrapper_44_reset = reset; // @[:@20234.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20236.4]
  assign RetimeWrapper_44_io_in = _T_739 & io_rPort_5_en_0; // @[package.scala 94:16:@20235.4]
  assign RetimeWrapper_45_clock = clock; // @[:@20241.4]
  assign RetimeWrapper_45_reset = reset; // @[:@20242.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20244.4]
  assign RetimeWrapper_45_io_in = _T_803 & io_rPort_5_en_0; // @[package.scala 94:16:@20243.4]
  assign RetimeWrapper_46_clock = clock; // @[:@20249.4]
  assign RetimeWrapper_46_reset = reset; // @[:@20250.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20252.4]
  assign RetimeWrapper_46_io_in = _T_867 & io_rPort_5_en_0; // @[package.scala 94:16:@20251.4]
  assign RetimeWrapper_47_clock = clock; // @[:@20257.4]
  assign RetimeWrapper_47_reset = reset; // @[:@20258.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20260.4]
  assign RetimeWrapper_47_io_in = _T_931 & io_rPort_5_en_0; // @[package.scala 94:16:@20259.4]
endmodule
module RetimeWrapper_233( // @[:@20771.2]
  input         clock, // @[:@20772.4]
  input         reset, // @[:@20773.4]
  input         io_flow, // @[:@20774.4]
  input  [31:0] io_in, // @[:@20774.4]
  output [31:0] io_out // @[:@20774.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20776.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20776.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20776.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20776.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20776.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20776.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@20776.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20789.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20788.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20787.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20786.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20785.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20783.4]
endmodule
module RetimeWrapper_235( // @[:@20835.2]
  input         clock, // @[:@20836.4]
  input         reset, // @[:@20837.4]
  input         io_flow, // @[:@20838.4]
  input  [31:0] io_in, // @[:@20838.4]
  output [31:0] io_out // @[:@20838.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20840.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20840.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20840.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20840.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20840.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20840.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@20840.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20853.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20852.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20851.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20850.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20849.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20847.4]
endmodule
module RetimeWrapper_243( // @[:@21385.2]
  input         clock, // @[:@21386.4]
  input         reset, // @[:@21387.4]
  input         io_flow, // @[:@21388.4]
  input  [31:0] io_in, // @[:@21388.4]
  output [31:0] io_out // @[:@21388.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@21390.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21403.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21402.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21401.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21400.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21399.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21397.4]
endmodule
module RetimeWrapper_246( // @[:@21481.2]
  input         clock, // @[:@21482.4]
  input         reset, // @[:@21483.4]
  input         io_flow, // @[:@21484.4]
  input  [31:0] io_in, // @[:@21484.4]
  output [31:0] io_out // @[:@21484.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@21486.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21499.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21498.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21497.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21496.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21495.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21493.4]
endmodule
module RetimeWrapper_247( // @[:@21513.2]
  input   clock, // @[:@21514.4]
  input   reset, // @[:@21515.4]
  input   io_flow, // @[:@21516.4]
  input   io_in, // @[:@21516.4]
  output  io_out // @[:@21516.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21518.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21518.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21518.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21518.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21518.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21518.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@21518.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21531.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21530.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21529.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21528.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21527.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21525.4]
endmodule
module RetimeWrapper_248( // @[:@21545.2]
  input         clock, // @[:@21546.4]
  input         reset, // @[:@21547.4]
  input         io_flow, // @[:@21548.4]
  input  [31:0] io_in, // @[:@21548.4]
  output [31:0] io_out // @[:@21548.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@21550.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21563.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21562.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21561.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21560.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21559.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21557.4]
endmodule
module RetimeWrapper_251( // @[:@21641.2]
  input         clock, // @[:@21642.4]
  input         reset, // @[:@21643.4]
  input         io_flow, // @[:@21644.4]
  input  [31:0] io_in, // @[:@21644.4]
  output [31:0] io_out // @[:@21644.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21646.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21646.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21646.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21646.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21646.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21646.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@21646.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21659.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21658.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21657.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21656.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21655.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21653.4]
endmodule
module RetimeWrapper_306( // @[:@25757.2]
  input         clock, // @[:@25758.4]
  input         reset, // @[:@25759.4]
  input         io_flow, // @[:@25760.4]
  input  [32:0] io_in, // @[:@25760.4]
  output [32:0] io_out // @[:@25760.4]
);
  wire [32:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25762.4]
  wire [32:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25762.4]
  wire [32:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25762.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25762.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25762.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25762.4]
  RetimeShiftRegister #(.WIDTH(33), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@25762.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25775.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25774.4]
  assign sr_init = 33'h0; // @[RetimeShiftRegister.scala 19:16:@25773.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25772.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25771.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25769.4]
endmodule
module RetimeWrapper_308( // @[:@25821.2]
  input         clock, // @[:@25822.4]
  input         reset, // @[:@25823.4]
  input         io_flow, // @[:@25824.4]
  input  [33:0] io_in, // @[:@25824.4]
  output [33:0] io_out // @[:@25824.4]
);
  wire [33:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25826.4]
  wire [33:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25826.4]
  wire [33:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25826.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25826.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25826.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25826.4]
  RetimeShiftRegister #(.WIDTH(34), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@25826.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25839.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25838.4]
  assign sr_init = 34'h0; // @[RetimeShiftRegister.scala 19:16:@25837.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25836.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25835.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25833.4]
endmodule
module fix2fixBox_78( // @[:@25937.2]
  input  [31:0] io_a, // @[:@25940.4]
  output [32:0] io_b // @[:@25940.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@25954.4]
endmodule
module __52( // @[:@25956.2]
  input  [31:0] io_b, // @[:@25959.4]
  output [32:0] io_result // @[:@25959.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@25964.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@25964.4]
  fix2fixBox_78 fix2fixBox ( // @[BigIPZynq.scala 219:30:@25964.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@25972.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@25967.4]
endmodule
module x406_x7( // @[:@26068.2]
  input         clock, // @[:@26069.4]
  input         reset, // @[:@26070.4]
  input  [31:0] io_a, // @[:@26071.4]
  input  [31:0] io_b, // @[:@26071.4]
  input         io_flow, // @[:@26071.4]
  output [31:0] io_result // @[:@26071.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@26079.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@26079.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@26086.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@26086.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@26096.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@26096.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@26096.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@26096.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@26096.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@26084.4 Math.scala 724:14:@26085.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@26091.4 Math.scala 724:14:@26092.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@26093.4]
  __52 _ ( // @[Math.scala 720:24:@26079.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __52 __1 ( // @[Math.scala 720:24:@26086.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@26096.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@26084.4 Math.scala 724:14:@26085.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@26091.4 Math.scala 724:14:@26092.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@26093.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@26104.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@26082.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@26089.4]
  assign fix2fixBox_clock = clock; // @[:@26097.4]
  assign fix2fixBox_reset = reset; // @[:@26098.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@26099.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@26102.4]
endmodule
module RetimeWrapper_321( // @[:@27196.2]
  input         clock, // @[:@27197.4]
  input         reset, // @[:@27198.4]
  input         io_flow, // @[:@27199.4]
  input  [31:0] io_in, // @[:@27199.4]
  output [31:0] io_out // @[:@27199.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27201.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27201.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27201.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27201.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27201.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27201.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@27201.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27214.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27213.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27212.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27211.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27210.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27208.4]
endmodule
module fix2fixBox_102( // @[:@27385.2]
  input  [31:0] io_a, // @[:@27388.4]
  output [31:0] io_b // @[:@27388.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@27398.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@27398.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@27401.4]
endmodule
module x414( // @[:@27403.2]
  input  [31:0] io_b, // @[:@27406.4]
  output [31:0] io_result // @[:@27406.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@27411.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@27411.4]
  fix2fixBox_102 fix2fixBox ( // @[BigIPZynq.scala 219:30:@27411.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@27419.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@27414.4]
endmodule
module Multiplier( // @[:@27431.2]
  input         clock, // @[:@27432.4]
  input         io_flow, // @[:@27434.4]
  input  [38:0] io_a, // @[:@27434.4]
  input  [38:0] io_b, // @[:@27434.4]
  output [38:0] io_out // @[:@27434.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@27436.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@27436.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@27436.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@27436.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@27436.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@27436.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@27446.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@27444.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@27443.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@27445.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@27442.4]
endmodule
module fix2fixBox_103( // @[:@27448.2]
  input  [38:0] io_a, // @[:@27451.4]
  output [31:0] io_b // @[:@27451.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@27459.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@27462.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@27459.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@27462.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@27465.4]
endmodule
module x415_mul( // @[:@27467.2]
  input         clock, // @[:@27468.4]
  input  [31:0] io_a, // @[:@27470.4]
  input  [31:0] io_b, // @[:@27470.4]
  input         io_flow, // @[:@27470.4]
  output [31:0] io_result // @[:@27470.4]
);
  wire  x415_mul_clock; // @[BigIPZynq.scala 63:21:@27485.4]
  wire  x415_mul_io_flow; // @[BigIPZynq.scala 63:21:@27485.4]
  wire [38:0] x415_mul_io_a; // @[BigIPZynq.scala 63:21:@27485.4]
  wire [38:0] x415_mul_io_b; // @[BigIPZynq.scala 63:21:@27485.4]
  wire [38:0] x415_mul_io_out; // @[BigIPZynq.scala 63:21:@27485.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@27493.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@27493.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@27477.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@27479.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@27481.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@27483.4]
  Multiplier x415_mul ( // @[BigIPZynq.scala 63:21:@27485.4]
    .clock(x415_mul_clock),
    .io_flow(x415_mul_io_flow),
    .io_a(x415_mul_io_a),
    .io_b(x415_mul_io_b),
    .io_out(x415_mul_io_out)
  );
  fix2fixBox_103 fix2fixBox ( // @[Math.scala 253:30:@27493.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@27477.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@27479.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@27481.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@27483.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@27501.4]
  assign x415_mul_clock = clock; // @[:@27486.4]
  assign x415_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@27490.4]
  assign x415_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@27488.4]
  assign x415_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@27489.4]
  assign fix2fixBox_io_a = x415_mul_io_out; // @[Math.scala 254:23:@27496.4]
endmodule
module fix2fixBox_104( // @[:@27503.2]
  input  [31:0] io_a, // @[:@27506.4]
  output [31:0] io_b // @[:@27506.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@27518.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@27518.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@27521.4]
endmodule
module x416( // @[:@27523.2]
  input  [31:0] io_b, // @[:@27526.4]
  output [31:0] io_result // @[:@27526.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@27531.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@27531.4]
  fix2fixBox_104 fix2fixBox ( // @[BigIPZynq.scala 219:30:@27531.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@27539.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@27534.4]
endmodule
module RetimeWrapper_340( // @[:@29349.2]
  input   clock, // @[:@29350.4]
  input   reset, // @[:@29351.4]
  input   io_flow, // @[:@29352.4]
  input   io_in, // @[:@29352.4]
  output  io_out // @[:@29352.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29354.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29354.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29354.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29354.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29354.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29354.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@29354.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29367.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29366.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29365.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29364.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29363.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29361.4]
endmodule
module RetimeWrapper_341( // @[:@29381.2]
  input         clock, // @[:@29382.4]
  input         reset, // @[:@29383.4]
  input         io_flow, // @[:@29384.4]
  input  [31:0] io_in, // @[:@29384.4]
  output [31:0] io_out // @[:@29384.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29386.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29386.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29386.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29386.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29386.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29386.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@29386.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29399.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29398.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29397.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29396.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29395.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29393.4]
endmodule
module RetimeWrapper_343( // @[:@29445.2]
  input         clock, // @[:@29446.4]
  input         reset, // @[:@29447.4]
  input         io_flow, // @[:@29448.4]
  input  [31:0] io_in, // @[:@29448.4]
  output [31:0] io_out // @[:@29448.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29450.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29450.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29450.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29450.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29450.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29450.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@29450.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29463.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29462.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29461.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29460.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29459.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29457.4]
endmodule
module RetimeWrapper_348( // @[:@29605.2]
  input         clock, // @[:@29606.4]
  input         reset, // @[:@29607.4]
  input         io_flow, // @[:@29608.4]
  input  [31:0] io_in, // @[:@29608.4]
  output [31:0] io_out // @[:@29608.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29610.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29610.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29610.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29610.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29610.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29610.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@29610.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29623.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29622.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29621.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29620.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29619.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29617.4]
endmodule
module RetimeWrapper_352( // @[:@29733.2]
  input   clock, // @[:@29734.4]
  input   reset, // @[:@29735.4]
  input   io_flow, // @[:@29736.4]
  input   io_in, // @[:@29736.4]
  output  io_out // @[:@29736.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29738.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29738.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29738.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29738.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29738.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29738.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@29738.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29751.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29750.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29749.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29748.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29747.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29745.4]
endmodule
module RetimeWrapper_355( // @[:@29829.2]
  input   clock, // @[:@29830.4]
  input   reset, // @[:@29831.4]
  input   io_flow, // @[:@29832.4]
  input   io_in, // @[:@29832.4]
  output  io_out // @[:@29832.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29834.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29834.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29834.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29834.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29834.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29834.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@29834.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29847.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29846.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29845.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29844.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29843.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29841.4]
endmodule
module RetimeWrapper_356( // @[:@29861.2]
  input         clock, // @[:@29862.4]
  input         reset, // @[:@29863.4]
  input         io_flow, // @[:@29864.4]
  input  [31:0] io_in, // @[:@29864.4]
  output [31:0] io_out // @[:@29864.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29866.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29866.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29866.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29866.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29866.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29866.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@29866.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29879.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29878.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@29877.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29876.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29875.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29873.4]
endmodule
module RetimeWrapper_358( // @[:@29925.2]
  input   clock, // @[:@29926.4]
  input   reset, // @[:@29927.4]
  input   io_flow, // @[:@29928.4]
  input   io_in, // @[:@29928.4]
  output  io_out // @[:@29928.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@29930.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@29930.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@29930.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29930.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29930.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29930.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@29930.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29943.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29942.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@29941.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29940.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29939.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29937.4]
endmodule
module RetimeWrapper_363( // @[:@30085.2]
  input         clock, // @[:@30086.4]
  input         reset, // @[:@30087.4]
  input         io_flow, // @[:@30088.4]
  input  [31:0] io_in, // @[:@30088.4]
  output [31:0] io_out // @[:@30088.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30090.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30090.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30090.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30090.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30090.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30090.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@30090.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30103.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30102.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30101.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30100.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30099.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30097.4]
endmodule
module RetimeWrapper_364( // @[:@30117.2]
  input         clock, // @[:@30118.4]
  input         reset, // @[:@30119.4]
  input         io_flow, // @[:@30120.4]
  input  [31:0] io_in, // @[:@30120.4]
  output [31:0] io_out // @[:@30120.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30122.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30122.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30122.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30122.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30122.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30122.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(16)) sr ( // @[RetimeShiftRegister.scala 15:20:@30122.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30135.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30134.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30133.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30132.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30131.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30129.4]
endmodule
module RetimeWrapper_367( // @[:@30213.2]
  input         clock, // @[:@30214.4]
  input         reset, // @[:@30215.4]
  input         io_flow, // @[:@30216.4]
  input  [31:0] io_in, // @[:@30216.4]
  output [31:0] io_out // @[:@30216.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30218.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30218.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30218.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30218.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30218.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30218.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(15)) sr ( // @[RetimeShiftRegister.scala 15:20:@30218.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30231.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30230.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30229.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30228.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30227.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30225.4]
endmodule
module RetimeWrapper_382( // @[:@31827.2]
  input         clock, // @[:@31828.4]
  input         reset, // @[:@31829.4]
  input         io_flow, // @[:@31830.4]
  input  [63:0] io_in, // @[:@31830.4]
  output [63:0] io_out // @[:@31830.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31832.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31832.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31832.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31832.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31832.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31832.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@31832.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31845.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31844.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@31843.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31842.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31841.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31839.4]
endmodule
module RetimeWrapper_383( // @[:@31859.2]
  input   clock, // @[:@31860.4]
  input   reset, // @[:@31861.4]
  input   io_flow, // @[:@31862.4]
  input   io_in, // @[:@31862.4]
  output  io_out // @[:@31862.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@31864.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@31864.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@31864.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31864.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31864.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31864.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@31864.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31877.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31876.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@31875.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31874.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31873.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31871.4]
endmodule
module x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@31943.2]
  input          clock, // @[:@31944.4]
  input          reset, // @[:@31945.4]
  output         io_in_x266_TREADY, // @[:@31946.4]
  input  [255:0] io_in_x266_TDATA, // @[:@31946.4]
  input  [7:0]   io_in_x266_TID, // @[:@31946.4]
  input  [7:0]   io_in_x266_TDEST, // @[:@31946.4]
  output         io_in_x267_TVALID, // @[:@31946.4]
  input          io_in_x267_TREADY, // @[:@31946.4]
  output [255:0] io_in_x267_TDATA, // @[:@31946.4]
  input          io_sigsIn_backpressure, // @[:@31946.4]
  input          io_sigsIn_datapathEn, // @[:@31946.4]
  input          io_sigsIn_break, // @[:@31946.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@31946.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@31946.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@31946.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@31946.4]
  input          io_rr // @[:@31946.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@31960.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@31960.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@31972.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@31972.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31995.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31995.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31995.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@31995.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@31995.4]
  wire  x301_lb_0_clock; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_reset; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_11_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_11_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_11_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_11_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_11_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_11_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_10_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_10_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_10_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_10_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_10_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_10_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_9_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_9_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_9_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_9_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_9_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_9_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_8_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_8_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_8_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_8_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_8_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_8_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_7_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_7_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_7_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_7_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_7_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_7_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_6_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_6_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_6_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_6_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_6_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_6_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_5_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_5_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_5_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_5_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_5_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_5_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_4_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_4_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_4_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_4_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_4_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_4_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_3_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_3_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_3_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_3_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_3_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_3_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_2_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_2_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_2_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_2_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_2_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_2_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_1_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_1_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_1_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_1_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_1_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_1_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_0_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_rPort_0_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_rPort_0_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_0_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_rPort_0_backpressure; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_rPort_0_output_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_wPort_1_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_wPort_1_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_wPort_1_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_wPort_1_data_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_wPort_1_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_wPort_0_banks_1; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [2:0] x301_lb_0_io_wPort_0_banks_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [8:0] x301_lb_0_io_wPort_0_ofs_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire [31:0] x301_lb_0_io_wPort_0_data_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x301_lb_0_io_wPort_0_en_0; // @[m_x301_lb_0.scala 39:17:@32005.4]
  wire  x302_lb2_0_clock; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_reset; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_5_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_5_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_rPort_5_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_5_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_5_backpressure; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_rPort_5_output_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_4_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_4_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_rPort_4_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_4_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_4_backpressure; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_rPort_4_output_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_3_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_3_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_rPort_3_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_3_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_3_backpressure; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_rPort_3_output_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_2_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_2_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_rPort_2_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_2_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_2_backpressure; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_rPort_2_output_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_1_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_1_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_rPort_1_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_1_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_1_backpressure; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_rPort_1_output_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_0_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_rPort_0_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_rPort_0_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_0_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_rPort_0_backpressure; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_rPort_0_output_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_wPort_1_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_wPort_1_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_wPort_1_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_wPort_1_data_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_wPort_1_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_wPort_0_banks_1; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [2:0] x302_lb2_0_io_wPort_0_banks_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [8:0] x302_lb2_0_io_wPort_0_ofs_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire [31:0] x302_lb2_0_io_wPort_0_data_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x302_lb2_0_io_wPort_0_en_0; // @[m_x302_lb2_0.scala 33:17:@32098.4]
  wire  x528_sub_1_clock; // @[Math.scala 191:24:@32225.4]
  wire  x528_sub_1_reset; // @[Math.scala 191:24:@32225.4]
  wire [31:0] x528_sub_1_io_a; // @[Math.scala 191:24:@32225.4]
  wire [31:0] x528_sub_1_io_b; // @[Math.scala 191:24:@32225.4]
  wire  x528_sub_1_io_flow; // @[Math.scala 191:24:@32225.4]
  wire [31:0] x528_sub_1_io_result; // @[Math.scala 191:24:@32225.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32252.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32252.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32252.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@32252.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@32252.4]
  wire  x311_sum_1_clock; // @[Math.scala 150:24:@32261.4]
  wire  x311_sum_1_reset; // @[Math.scala 150:24:@32261.4]
  wire [31:0] x311_sum_1_io_a; // @[Math.scala 150:24:@32261.4]
  wire [31:0] x311_sum_1_io_b; // @[Math.scala 150:24:@32261.4]
  wire  x311_sum_1_io_flow; // @[Math.scala 150:24:@32261.4]
  wire [31:0] x311_sum_1_io_result; // @[Math.scala 150:24:@32261.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32271.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32271.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32271.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32271.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32271.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32280.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32280.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32280.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@32280.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@32280.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@32298.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@32298.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@32298.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@32298.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@32298.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@32307.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@32307.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@32307.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@32307.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@32307.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@32316.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@32316.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@32316.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@32316.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@32316.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@32327.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@32327.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@32327.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@32327.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@32327.4]
  wire  x313_rdcol_1_clock; // @[Math.scala 150:24:@32350.4]
  wire  x313_rdcol_1_reset; // @[Math.scala 150:24:@32350.4]
  wire [31:0] x313_rdcol_1_io_a; // @[Math.scala 150:24:@32350.4]
  wire [31:0] x313_rdcol_1_io_b; // @[Math.scala 150:24:@32350.4]
  wire  x313_rdcol_1_io_flow; // @[Math.scala 150:24:@32350.4]
  wire [31:0] x313_rdcol_1_io_result; // @[Math.scala 150:24:@32350.4]
  wire  x317_sum_1_clock; // @[Math.scala 150:24:@32390.4]
  wire  x317_sum_1_reset; // @[Math.scala 150:24:@32390.4]
  wire [31:0] x317_sum_1_io_a; // @[Math.scala 150:24:@32390.4]
  wire [31:0] x317_sum_1_io_b; // @[Math.scala 150:24:@32390.4]
  wire  x317_sum_1_io_flow; // @[Math.scala 150:24:@32390.4]
  wire [31:0] x317_sum_1_io_result; // @[Math.scala 150:24:@32390.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@32400.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@32400.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@32400.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@32400.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@32400.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@32409.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@32409.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@32409.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@32409.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@32409.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@32418.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@32418.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@32418.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@32418.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@32418.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@32429.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@32429.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@32429.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@32429.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@32429.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@32450.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@32450.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@32466.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@32466.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@32466.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@32466.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@32466.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@32482.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@32482.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@32482.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@32482.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@32482.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@32497.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@32497.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@32497.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@32497.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@32497.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@32506.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@32506.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@32506.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@32506.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@32506.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@32515.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@32515.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@32524.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@32524.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@32524.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@32524.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@32524.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@32533.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@32533.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@32533.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@32533.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@32533.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@32542.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@32542.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@32542.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@32542.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@32542.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@32554.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@32554.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@32554.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@32554.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@32554.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@32575.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@32575.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@32575.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@32575.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@32575.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@32599.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@32599.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@32599.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@32599.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@32599.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@32608.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@32608.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@32608.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@32608.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@32608.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@32617.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@32617.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@32629.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@32629.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@32629.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@32629.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@32629.4]
  wire  x331_rdcol_1_clock; // @[Math.scala 150:24:@32652.4]
  wire  x331_rdcol_1_reset; // @[Math.scala 150:24:@32652.4]
  wire [31:0] x331_rdcol_1_io_a; // @[Math.scala 150:24:@32652.4]
  wire [31:0] x331_rdcol_1_io_b; // @[Math.scala 150:24:@32652.4]
  wire  x331_rdcol_1_io_flow; // @[Math.scala 150:24:@32652.4]
  wire [31:0] x331_rdcol_1_io_result; // @[Math.scala 150:24:@32652.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@32703.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@32703.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@32703.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@32703.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@32703.4]
  wire  x337_sum_1_clock; // @[Math.scala 150:24:@32712.4]
  wire  x337_sum_1_reset; // @[Math.scala 150:24:@32712.4]
  wire [31:0] x337_sum_1_io_a; // @[Math.scala 150:24:@32712.4]
  wire [31:0] x337_sum_1_io_b; // @[Math.scala 150:24:@32712.4]
  wire  x337_sum_1_io_flow; // @[Math.scala 150:24:@32712.4]
  wire [31:0] x337_sum_1_io_result; // @[Math.scala 150:24:@32712.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@32722.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@32722.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@32722.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@32722.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@32722.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@32731.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@32731.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@32731.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@32731.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@32731.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@32740.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@32740.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@32740.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@32740.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@32740.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@32752.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@32752.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@32752.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@32752.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@32752.4]
  wire  x340_rdcol_1_clock; // @[Math.scala 150:24:@32775.4]
  wire  x340_rdcol_1_reset; // @[Math.scala 150:24:@32775.4]
  wire [31:0] x340_rdcol_1_io_a; // @[Math.scala 150:24:@32775.4]
  wire [31:0] x340_rdcol_1_io_b; // @[Math.scala 150:24:@32775.4]
  wire  x340_rdcol_1_io_flow; // @[Math.scala 150:24:@32775.4]
  wire [31:0] x340_rdcol_1_io_result; // @[Math.scala 150:24:@32775.4]
  wire  x346_sum_1_clock; // @[Math.scala 150:24:@32826.4]
  wire  x346_sum_1_reset; // @[Math.scala 150:24:@32826.4]
  wire [31:0] x346_sum_1_io_a; // @[Math.scala 150:24:@32826.4]
  wire [31:0] x346_sum_1_io_b; // @[Math.scala 150:24:@32826.4]
  wire  x346_sum_1_io_flow; // @[Math.scala 150:24:@32826.4]
  wire [31:0] x346_sum_1_io_result; // @[Math.scala 150:24:@32826.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@32836.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@32836.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@32836.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@32836.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@32836.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@32845.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@32845.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@32854.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@32854.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@32854.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@32854.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@32854.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@32866.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@32866.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@32866.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@32866.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@32866.4]
  wire  x349_rdrow_1_clock; // @[Math.scala 191:24:@32889.4]
  wire  x349_rdrow_1_reset; // @[Math.scala 191:24:@32889.4]
  wire [31:0] x349_rdrow_1_io_a; // @[Math.scala 191:24:@32889.4]
  wire [31:0] x349_rdrow_1_io_b; // @[Math.scala 191:24:@32889.4]
  wire  x349_rdrow_1_io_flow; // @[Math.scala 191:24:@32889.4]
  wire [31:0] x349_rdrow_1_io_result; // @[Math.scala 191:24:@32889.4]
  wire  x536_sub_1_clock; // @[Math.scala 191:24:@32961.4]
  wire  x536_sub_1_reset; // @[Math.scala 191:24:@32961.4]
  wire [31:0] x536_sub_1_io_a; // @[Math.scala 191:24:@32961.4]
  wire [31:0] x536_sub_1_io_b; // @[Math.scala 191:24:@32961.4]
  wire  x536_sub_1_io_flow; // @[Math.scala 191:24:@32961.4]
  wire [31:0] x536_sub_1_io_result; // @[Math.scala 191:24:@32961.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@32971.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@32971.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@32971.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@32971.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@32971.4]
  wire  x357_sum_1_clock; // @[Math.scala 150:24:@32980.4]
  wire  x357_sum_1_reset; // @[Math.scala 150:24:@32980.4]
  wire [31:0] x357_sum_1_io_a; // @[Math.scala 150:24:@32980.4]
  wire [31:0] x357_sum_1_io_b; // @[Math.scala 150:24:@32980.4]
  wire  x357_sum_1_io_flow; // @[Math.scala 150:24:@32980.4]
  wire [31:0] x357_sum_1_io_result; // @[Math.scala 150:24:@32980.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@32990.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@32990.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@32990.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@32990.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@32990.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@32999.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@33011.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@33011.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@33011.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@33011.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@33011.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@33032.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@33032.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@33032.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@33032.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@33032.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@33047.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@33047.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@33047.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@33047.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@33047.4]
  wire  x362_sum_1_clock; // @[Math.scala 150:24:@33058.4]
  wire  x362_sum_1_reset; // @[Math.scala 150:24:@33058.4]
  wire [31:0] x362_sum_1_io_a; // @[Math.scala 150:24:@33058.4]
  wire [31:0] x362_sum_1_io_b; // @[Math.scala 150:24:@33058.4]
  wire  x362_sum_1_io_flow; // @[Math.scala 150:24:@33058.4]
  wire [31:0] x362_sum_1_io_result; // @[Math.scala 150:24:@33058.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@33068.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@33068.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@33068.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@33068.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@33068.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@33080.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@33107.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@33107.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@33107.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@33107.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@33107.4]
  wire  x367_sum_1_clock; // @[Math.scala 150:24:@33116.4]
  wire  x367_sum_1_reset; // @[Math.scala 150:24:@33116.4]
  wire [31:0] x367_sum_1_io_a; // @[Math.scala 150:24:@33116.4]
  wire [31:0] x367_sum_1_io_b; // @[Math.scala 150:24:@33116.4]
  wire  x367_sum_1_io_flow; // @[Math.scala 150:24:@33116.4]
  wire [31:0] x367_sum_1_io_result; // @[Math.scala 150:24:@33116.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@33126.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@33126.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@33126.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@33126.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@33126.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@33138.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@33138.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@33138.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@33138.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@33138.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@33165.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@33165.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@33165.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@33165.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@33165.4]
  wire  x372_sum_1_clock; // @[Math.scala 150:24:@33174.4]
  wire  x372_sum_1_reset; // @[Math.scala 150:24:@33174.4]
  wire [31:0] x372_sum_1_io_a; // @[Math.scala 150:24:@33174.4]
  wire [31:0] x372_sum_1_io_b; // @[Math.scala 150:24:@33174.4]
  wire  x372_sum_1_io_flow; // @[Math.scala 150:24:@33174.4]
  wire [31:0] x372_sum_1_io_result; // @[Math.scala 150:24:@33174.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@33184.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@33184.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@33184.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@33184.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@33184.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@33196.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@33196.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@33196.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@33196.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@33196.4]
  wire  x375_rdrow_1_clock; // @[Math.scala 191:24:@33219.4]
  wire  x375_rdrow_1_reset; // @[Math.scala 191:24:@33219.4]
  wire [31:0] x375_rdrow_1_io_a; // @[Math.scala 191:24:@33219.4]
  wire [31:0] x375_rdrow_1_io_b; // @[Math.scala 191:24:@33219.4]
  wire  x375_rdrow_1_io_flow; // @[Math.scala 191:24:@33219.4]
  wire [31:0] x375_rdrow_1_io_result; // @[Math.scala 191:24:@33219.4]
  wire  x541_sub_1_clock; // @[Math.scala 191:24:@33291.4]
  wire  x541_sub_1_reset; // @[Math.scala 191:24:@33291.4]
  wire [31:0] x541_sub_1_io_a; // @[Math.scala 191:24:@33291.4]
  wire [31:0] x541_sub_1_io_b; // @[Math.scala 191:24:@33291.4]
  wire  x541_sub_1_io_flow; // @[Math.scala 191:24:@33291.4]
  wire [31:0] x541_sub_1_io_result; // @[Math.scala 191:24:@33291.4]
  wire  x383_sum_1_clock; // @[Math.scala 150:24:@33301.4]
  wire  x383_sum_1_reset; // @[Math.scala 150:24:@33301.4]
  wire [31:0] x383_sum_1_io_a; // @[Math.scala 150:24:@33301.4]
  wire [31:0] x383_sum_1_io_b; // @[Math.scala 150:24:@33301.4]
  wire  x383_sum_1_io_flow; // @[Math.scala 150:24:@33301.4]
  wire [31:0] x383_sum_1_io_result; // @[Math.scala 150:24:@33301.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@33311.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@33311.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@33311.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@33311.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@33311.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@33320.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@33320.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@33332.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@33332.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@33332.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@33332.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@33332.4]
  wire  x388_sum_1_clock; // @[Math.scala 150:24:@33359.4]
  wire  x388_sum_1_reset; // @[Math.scala 150:24:@33359.4]
  wire [31:0] x388_sum_1_io_a; // @[Math.scala 150:24:@33359.4]
  wire [31:0] x388_sum_1_io_b; // @[Math.scala 150:24:@33359.4]
  wire  x388_sum_1_io_flow; // @[Math.scala 150:24:@33359.4]
  wire [31:0] x388_sum_1_io_result; // @[Math.scala 150:24:@33359.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@33369.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@33369.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@33369.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@33369.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@33369.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@33381.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@33381.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@33381.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@33381.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@33381.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@33408.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@33408.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@33408.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@33408.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@33408.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@33408.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@33430.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@33430.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@33430.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@33430.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@33430.4]
  wire  x398_sum_1_clock; // @[Math.scala 150:24:@33459.4]
  wire  x398_sum_1_reset; // @[Math.scala 150:24:@33459.4]
  wire [31:0] x398_sum_1_io_a; // @[Math.scala 150:24:@33459.4]
  wire [31:0] x398_sum_1_io_b; // @[Math.scala 150:24:@33459.4]
  wire  x398_sum_1_io_flow; // @[Math.scala 150:24:@33459.4]
  wire [31:0] x398_sum_1_io_result; // @[Math.scala 150:24:@33459.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@33469.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@33469.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@33469.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@33469.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@33469.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@33481.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@33481.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@33481.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@33481.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@33481.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@33504.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@33504.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@33504.4]
  wire [32:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@33504.4]
  wire [32:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@33504.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@33516.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@33516.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@33516.4]
  wire [32:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@33516.4]
  wire [32:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@33516.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@33528.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@33528.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@33528.4]
  wire [33:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@33528.4]
  wire [33:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@33528.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@33540.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@33540.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@33540.4]
  wire [32:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@33540.4]
  wire [32:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@33540.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@33552.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@33552.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@33552.4]
  wire [32:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@33552.4]
  wire [32:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@33552.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@33562.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@33562.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@33562.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@33562.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@33562.4]
  wire  x406_x7_1_clock; // @[Math.scala 150:24:@33571.4]
  wire  x406_x7_1_reset; // @[Math.scala 150:24:@33571.4]
  wire [31:0] x406_x7_1_io_a; // @[Math.scala 150:24:@33571.4]
  wire [31:0] x406_x7_1_io_b; // @[Math.scala 150:24:@33571.4]
  wire  x406_x7_1_io_flow; // @[Math.scala 150:24:@33571.4]
  wire [31:0] x406_x7_1_io_result; // @[Math.scala 150:24:@33571.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@33581.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@33581.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@33581.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@33581.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@33581.4]
  wire  x407_x8_1_clock; // @[Math.scala 150:24:@33590.4]
  wire  x407_x8_1_reset; // @[Math.scala 150:24:@33590.4]
  wire [31:0] x407_x8_1_io_a; // @[Math.scala 150:24:@33590.4]
  wire [31:0] x407_x8_1_io_b; // @[Math.scala 150:24:@33590.4]
  wire  x407_x8_1_io_flow; // @[Math.scala 150:24:@33590.4]
  wire [31:0] x407_x8_1_io_result; // @[Math.scala 150:24:@33590.4]
  wire  x408_x7_1_clock; // @[Math.scala 150:24:@33600.4]
  wire  x408_x7_1_reset; // @[Math.scala 150:24:@33600.4]
  wire [31:0] x408_x7_1_io_a; // @[Math.scala 150:24:@33600.4]
  wire [31:0] x408_x7_1_io_b; // @[Math.scala 150:24:@33600.4]
  wire  x408_x7_1_io_flow; // @[Math.scala 150:24:@33600.4]
  wire [31:0] x408_x7_1_io_result; // @[Math.scala 150:24:@33600.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@33610.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@33610.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@33610.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@33610.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@33610.4]
  wire  x409_x8_1_clock; // @[Math.scala 150:24:@33619.4]
  wire  x409_x8_1_reset; // @[Math.scala 150:24:@33619.4]
  wire [31:0] x409_x8_1_io_a; // @[Math.scala 150:24:@33619.4]
  wire [31:0] x409_x8_1_io_b; // @[Math.scala 150:24:@33619.4]
  wire  x409_x8_1_io_flow; // @[Math.scala 150:24:@33619.4]
  wire [31:0] x409_x8_1_io_result; // @[Math.scala 150:24:@33619.4]
  wire  x410_x7_1_clock; // @[Math.scala 150:24:@33629.4]
  wire  x410_x7_1_reset; // @[Math.scala 150:24:@33629.4]
  wire [31:0] x410_x7_1_io_a; // @[Math.scala 150:24:@33629.4]
  wire [31:0] x410_x7_1_io_b; // @[Math.scala 150:24:@33629.4]
  wire  x410_x7_1_io_flow; // @[Math.scala 150:24:@33629.4]
  wire [31:0] x410_x7_1_io_result; // @[Math.scala 150:24:@33629.4]
  wire  x411_x8_1_clock; // @[Math.scala 150:24:@33639.4]
  wire  x411_x8_1_reset; // @[Math.scala 150:24:@33639.4]
  wire [31:0] x411_x8_1_io_a; // @[Math.scala 150:24:@33639.4]
  wire [31:0] x411_x8_1_io_b; // @[Math.scala 150:24:@33639.4]
  wire  x411_x8_1_io_flow; // @[Math.scala 150:24:@33639.4]
  wire [31:0] x411_x8_1_io_result; // @[Math.scala 150:24:@33639.4]
  wire  x412_x7_1_clock; // @[Math.scala 150:24:@33649.4]
  wire  x412_x7_1_reset; // @[Math.scala 150:24:@33649.4]
  wire [31:0] x412_x7_1_io_a; // @[Math.scala 150:24:@33649.4]
  wire [31:0] x412_x7_1_io_b; // @[Math.scala 150:24:@33649.4]
  wire  x412_x7_1_io_flow; // @[Math.scala 150:24:@33649.4]
  wire [31:0] x412_x7_1_io_result; // @[Math.scala 150:24:@33649.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@33659.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@33659.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@33659.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@33659.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@33659.4]
  wire  x413_sum_1_clock; // @[Math.scala 150:24:@33668.4]
  wire  x413_sum_1_reset; // @[Math.scala 150:24:@33668.4]
  wire [31:0] x413_sum_1_io_a; // @[Math.scala 150:24:@33668.4]
  wire [31:0] x413_sum_1_io_b; // @[Math.scala 150:24:@33668.4]
  wire  x413_sum_1_io_flow; // @[Math.scala 150:24:@33668.4]
  wire [31:0] x413_sum_1_io_result; // @[Math.scala 150:24:@33668.4]
  wire [31:0] x414_1_io_b; // @[Math.scala 720:24:@33678.4]
  wire [31:0] x414_1_io_result; // @[Math.scala 720:24:@33678.4]
  wire  x415_mul_1_clock; // @[Math.scala 262:24:@33689.4]
  wire [31:0] x415_mul_1_io_a; // @[Math.scala 262:24:@33689.4]
  wire [31:0] x415_mul_1_io_b; // @[Math.scala 262:24:@33689.4]
  wire  x415_mul_1_io_flow; // @[Math.scala 262:24:@33689.4]
  wire [31:0] x415_mul_1_io_result; // @[Math.scala 262:24:@33689.4]
  wire [31:0] x416_1_io_b; // @[Math.scala 720:24:@33699.4]
  wire [31:0] x416_1_io_result; // @[Math.scala 720:24:@33699.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@33710.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@33710.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@33710.4]
  wire [32:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@33710.4]
  wire [32:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@33710.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@33722.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@33722.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@33722.4]
  wire [32:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@33722.4]
  wire [32:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@33722.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@33734.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@33734.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@33734.4]
  wire [33:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@33734.4]
  wire [33:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@33734.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@33746.4]
  wire [32:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@33746.4]
  wire [32:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@33746.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@33758.4]
  wire [32:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@33758.4]
  wire [32:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@33768.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@33768.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@33768.4]
  wire [31:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@33768.4]
  wire [31:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@33768.4]
  wire  x422_x7_1_clock; // @[Math.scala 150:24:@33777.4]
  wire  x422_x7_1_reset; // @[Math.scala 150:24:@33777.4]
  wire [31:0] x422_x7_1_io_a; // @[Math.scala 150:24:@33777.4]
  wire [31:0] x422_x7_1_io_b; // @[Math.scala 150:24:@33777.4]
  wire  x422_x7_1_io_flow; // @[Math.scala 150:24:@33777.4]
  wire [31:0] x422_x7_1_io_result; // @[Math.scala 150:24:@33777.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@33787.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@33787.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@33787.4]
  wire [31:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@33787.4]
  wire [31:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@33787.4]
  wire  x423_x8_1_clock; // @[Math.scala 150:24:@33796.4]
  wire  x423_x8_1_reset; // @[Math.scala 150:24:@33796.4]
  wire [31:0] x423_x8_1_io_a; // @[Math.scala 150:24:@33796.4]
  wire [31:0] x423_x8_1_io_b; // @[Math.scala 150:24:@33796.4]
  wire  x423_x8_1_io_flow; // @[Math.scala 150:24:@33796.4]
  wire [31:0] x423_x8_1_io_result; // @[Math.scala 150:24:@33796.4]
  wire  x424_x7_1_clock; // @[Math.scala 150:24:@33806.4]
  wire  x424_x7_1_reset; // @[Math.scala 150:24:@33806.4]
  wire [31:0] x424_x7_1_io_a; // @[Math.scala 150:24:@33806.4]
  wire [31:0] x424_x7_1_io_b; // @[Math.scala 150:24:@33806.4]
  wire  x424_x7_1_io_flow; // @[Math.scala 150:24:@33806.4]
  wire [31:0] x424_x7_1_io_result; // @[Math.scala 150:24:@33806.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@33816.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@33816.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@33816.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@33816.4]
  wire  x425_x8_1_clock; // @[Math.scala 150:24:@33825.4]
  wire  x425_x8_1_reset; // @[Math.scala 150:24:@33825.4]
  wire [31:0] x425_x8_1_io_a; // @[Math.scala 150:24:@33825.4]
  wire [31:0] x425_x8_1_io_b; // @[Math.scala 150:24:@33825.4]
  wire  x425_x8_1_io_flow; // @[Math.scala 150:24:@33825.4]
  wire [31:0] x425_x8_1_io_result; // @[Math.scala 150:24:@33825.4]
  wire  x426_x7_1_clock; // @[Math.scala 150:24:@33835.4]
  wire  x426_x7_1_reset; // @[Math.scala 150:24:@33835.4]
  wire [31:0] x426_x7_1_io_a; // @[Math.scala 150:24:@33835.4]
  wire [31:0] x426_x7_1_io_b; // @[Math.scala 150:24:@33835.4]
  wire  x426_x7_1_io_flow; // @[Math.scala 150:24:@33835.4]
  wire [31:0] x426_x7_1_io_result; // @[Math.scala 150:24:@33835.4]
  wire  x427_x8_1_clock; // @[Math.scala 150:24:@33845.4]
  wire  x427_x8_1_reset; // @[Math.scala 150:24:@33845.4]
  wire [31:0] x427_x8_1_io_a; // @[Math.scala 150:24:@33845.4]
  wire [31:0] x427_x8_1_io_b; // @[Math.scala 150:24:@33845.4]
  wire  x427_x8_1_io_flow; // @[Math.scala 150:24:@33845.4]
  wire [31:0] x427_x8_1_io_result; // @[Math.scala 150:24:@33845.4]
  wire  x428_x7_1_clock; // @[Math.scala 150:24:@33855.4]
  wire  x428_x7_1_reset; // @[Math.scala 150:24:@33855.4]
  wire [31:0] x428_x7_1_io_a; // @[Math.scala 150:24:@33855.4]
  wire [31:0] x428_x7_1_io_b; // @[Math.scala 150:24:@33855.4]
  wire  x428_x7_1_io_flow; // @[Math.scala 150:24:@33855.4]
  wire [31:0] x428_x7_1_io_result; // @[Math.scala 150:24:@33855.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@33865.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@33865.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@33865.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@33865.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@33865.4]
  wire  x429_sum_1_clock; // @[Math.scala 150:24:@33874.4]
  wire  x429_sum_1_reset; // @[Math.scala 150:24:@33874.4]
  wire [31:0] x429_sum_1_io_a; // @[Math.scala 150:24:@33874.4]
  wire [31:0] x429_sum_1_io_b; // @[Math.scala 150:24:@33874.4]
  wire  x429_sum_1_io_flow; // @[Math.scala 150:24:@33874.4]
  wire [31:0] x429_sum_1_io_result; // @[Math.scala 150:24:@33874.4]
  wire [31:0] x430_1_io_b; // @[Math.scala 720:24:@33884.4]
  wire [31:0] x430_1_io_result; // @[Math.scala 720:24:@33884.4]
  wire  x431_mul_1_clock; // @[Math.scala 262:24:@33895.4]
  wire [31:0] x431_mul_1_io_a; // @[Math.scala 262:24:@33895.4]
  wire [31:0] x431_mul_1_io_b; // @[Math.scala 262:24:@33895.4]
  wire  x431_mul_1_io_flow; // @[Math.scala 262:24:@33895.4]
  wire [31:0] x431_mul_1_io_result; // @[Math.scala 262:24:@33895.4]
  wire [31:0] x432_1_io_b; // @[Math.scala 720:24:@33905.4]
  wire [31:0] x432_1_io_result; // @[Math.scala 720:24:@33905.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@33914.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@33923.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@33923.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@33923.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@33932.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@33941.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@33941.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@33941.4]
  wire [31:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@33941.4]
  wire [31:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@33941.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@33950.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@33950.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@33950.4]
  wire [31:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@33950.4]
  wire [31:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@33950.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@33959.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@33959.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@33959.4]
  wire [31:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@33959.4]
  wire [31:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@33959.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@33991.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@33991.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@33991.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@34000.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@34000.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@34000.4]
  wire [31:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@34000.4]
  wire [31:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@34000.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@34009.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@34009.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@34009.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@34009.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@34009.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@34041.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@34041.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@34050.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@34050.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@34050.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@34050.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@34050.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@34059.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@34059.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@34059.4]
  wire [31:0] RetimeWrapper_91_io_in; // @[package.scala 93:22:@34059.4]
  wire [31:0] RetimeWrapper_91_io_out; // @[package.scala 93:22:@34059.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@34068.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@34068.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@34068.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@34068.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@34068.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@34077.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@34077.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@34077.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@34077.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@34077.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@34086.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@34086.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@34086.4]
  wire [31:0] RetimeWrapper_94_io_in; // @[package.scala 93:22:@34086.4]
  wire [31:0] RetimeWrapper_94_io_out; // @[package.scala 93:22:@34086.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@34098.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@34098.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@34098.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@34098.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@34098.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@34119.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@34119.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@34119.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@34119.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@34119.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@34128.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@34128.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@34128.4]
  wire [31:0] RetimeWrapper_97_io_in; // @[package.scala 93:22:@34128.4]
  wire [31:0] RetimeWrapper_97_io_out; // @[package.scala 93:22:@34128.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@34137.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@34137.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@34137.4]
  wire [31:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@34137.4]
  wire [31:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@34137.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@34149.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@34149.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@34149.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@34149.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@34149.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@34170.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@34170.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@34170.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@34170.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@34170.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@34179.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@34179.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@34179.4]
  wire [31:0] RetimeWrapper_101_io_in; // @[package.scala 93:22:@34179.4]
  wire [31:0] RetimeWrapper_101_io_out; // @[package.scala 93:22:@34179.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@34188.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@34188.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@34188.4]
  wire [31:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@34188.4]
  wire [31:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@34188.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@34200.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@34221.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@34221.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@34221.4]
  wire [31:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@34221.4]
  wire [31:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@34221.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@34230.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@34230.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@34230.4]
  wire [31:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@34230.4]
  wire [31:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@34230.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@34239.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@34239.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@34239.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@34239.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@34239.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@34251.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@34272.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@34272.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@34272.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@34272.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@34272.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@34281.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@34281.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@34281.4]
  wire [31:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@34281.4]
  wire [31:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@34281.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@34293.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@34293.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@34293.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@34293.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@34293.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@34314.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@34323.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@34323.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@34323.4]
  wire [31:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@34323.4]
  wire [31:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@34323.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@34335.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@34335.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@34335.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@34335.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@34335.4]
  wire  x451_x9_1_clock; // @[Math.scala 150:24:@34368.4]
  wire  x451_x9_1_reset; // @[Math.scala 150:24:@34368.4]
  wire [31:0] x451_x9_1_io_a; // @[Math.scala 150:24:@34368.4]
  wire [31:0] x451_x9_1_io_b; // @[Math.scala 150:24:@34368.4]
  wire  x451_x9_1_io_flow; // @[Math.scala 150:24:@34368.4]
  wire [31:0] x451_x9_1_io_result; // @[Math.scala 150:24:@34368.4]
  wire  x452_x10_1_clock; // @[Math.scala 150:24:@34378.4]
  wire  x452_x10_1_reset; // @[Math.scala 150:24:@34378.4]
  wire [31:0] x452_x10_1_io_a; // @[Math.scala 150:24:@34378.4]
  wire [31:0] x452_x10_1_io_b; // @[Math.scala 150:24:@34378.4]
  wire  x452_x10_1_io_flow; // @[Math.scala 150:24:@34378.4]
  wire [31:0] x452_x10_1_io_result; // @[Math.scala 150:24:@34378.4]
  wire  x453_sum_1_clock; // @[Math.scala 150:24:@34388.4]
  wire  x453_sum_1_reset; // @[Math.scala 150:24:@34388.4]
  wire [31:0] x453_sum_1_io_a; // @[Math.scala 150:24:@34388.4]
  wire [31:0] x453_sum_1_io_b; // @[Math.scala 150:24:@34388.4]
  wire  x453_sum_1_io_flow; // @[Math.scala 150:24:@34388.4]
  wire [31:0] x453_sum_1_io_result; // @[Math.scala 150:24:@34388.4]
  wire [31:0] x454_1_io_b; // @[Math.scala 720:24:@34398.4]
  wire [31:0] x454_1_io_result; // @[Math.scala 720:24:@34398.4]
  wire  x455_mul_1_clock; // @[Math.scala 262:24:@34409.4]
  wire [31:0] x455_mul_1_io_a; // @[Math.scala 262:24:@34409.4]
  wire [31:0] x455_mul_1_io_b; // @[Math.scala 262:24:@34409.4]
  wire  x455_mul_1_io_flow; // @[Math.scala 262:24:@34409.4]
  wire [31:0] x455_mul_1_io_result; // @[Math.scala 262:24:@34409.4]
  wire [31:0] x456_1_io_b; // @[Math.scala 720:24:@34421.4]
  wire [31:0] x456_1_io_result; // @[Math.scala 720:24:@34421.4]
  wire  x459_x9_1_clock; // @[Math.scala 150:24:@34440.4]
  wire  x459_x9_1_reset; // @[Math.scala 150:24:@34440.4]
  wire [31:0] x459_x9_1_io_a; // @[Math.scala 150:24:@34440.4]
  wire [31:0] x459_x9_1_io_b; // @[Math.scala 150:24:@34440.4]
  wire  x459_x9_1_io_flow; // @[Math.scala 150:24:@34440.4]
  wire [31:0] x459_x9_1_io_result; // @[Math.scala 150:24:@34440.4]
  wire  x460_x10_1_clock; // @[Math.scala 150:24:@34450.4]
  wire  x460_x10_1_reset; // @[Math.scala 150:24:@34450.4]
  wire [31:0] x460_x10_1_io_a; // @[Math.scala 150:24:@34450.4]
  wire [31:0] x460_x10_1_io_b; // @[Math.scala 150:24:@34450.4]
  wire  x460_x10_1_io_flow; // @[Math.scala 150:24:@34450.4]
  wire [31:0] x460_x10_1_io_result; // @[Math.scala 150:24:@34450.4]
  wire  x461_sum_1_clock; // @[Math.scala 150:24:@34460.4]
  wire  x461_sum_1_reset; // @[Math.scala 150:24:@34460.4]
  wire [31:0] x461_sum_1_io_a; // @[Math.scala 150:24:@34460.4]
  wire [31:0] x461_sum_1_io_b; // @[Math.scala 150:24:@34460.4]
  wire  x461_sum_1_io_flow; // @[Math.scala 150:24:@34460.4]
  wire [31:0] x461_sum_1_io_result; // @[Math.scala 150:24:@34460.4]
  wire [31:0] x462_1_io_b; // @[Math.scala 720:24:@34470.4]
  wire [31:0] x462_1_io_result; // @[Math.scala 720:24:@34470.4]
  wire  x463_mul_1_clock; // @[Math.scala 262:24:@34481.4]
  wire [31:0] x463_mul_1_io_a; // @[Math.scala 262:24:@34481.4]
  wire [31:0] x463_mul_1_io_b; // @[Math.scala 262:24:@34481.4]
  wire  x463_mul_1_io_flow; // @[Math.scala 262:24:@34481.4]
  wire [31:0] x463_mul_1_io_result; // @[Math.scala 262:24:@34481.4]
  wire [31:0] x464_1_io_b; // @[Math.scala 720:24:@34491.4]
  wire [31:0] x464_1_io_result; // @[Math.scala 720:24:@34491.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@34506.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@34506.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@34506.4]
  wire [63:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@34506.4]
  wire [63:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@34506.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@34515.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@34515.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@34515.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@34515.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@34515.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@34524.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@34524.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@34524.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@34524.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@34524.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@34533.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@34533.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@34533.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@34533.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@34533.4]
  wire  b297; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 62:18:@31980.4]
  wire  b298; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 63:18:@31981.4]
  wire  _T_205; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 67:30:@31983.4]
  wire  _T_206; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 67:37:@31984.4]
  wire  _T_210; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:76:@31989.4]
  wire  _T_211; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:62:@31990.4]
  wire  _T_213; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:101:@31991.4]
  wire [63:0] x547_x299_D1_0_number; // @[package.scala 96:25:@32000.4 package.scala 96:25:@32001.4]
  wire [31:0] b295_number; // @[Math.scala 723:22:@31965.4 Math.scala 724:14:@31966.4]
  wire [31:0] _T_244; // @[Math.scala 406:49:@32166.4]
  wire [31:0] _T_246; // @[Math.scala 406:56:@32168.4]
  wire [31:0] _T_247; // @[Math.scala 406:56:@32169.4]
  wire [31:0] x523_number; // @[implicits.scala 133:21:@32170.4]
  wire [31:0] _T_257; // @[Math.scala 406:49:@32179.4]
  wire [31:0] _T_259; // @[Math.scala 406:56:@32181.4]
  wire [31:0] _T_260; // @[Math.scala 406:56:@32182.4]
  wire [31:0] b296_number; // @[Math.scala 723:22:@31977.4 Math.scala 724:14:@31978.4]
  wire [31:0] _T_269; // @[Math.scala 406:49:@32190.4]
  wire [31:0] _T_271; // @[Math.scala 406:56:@32192.4]
  wire [31:0] _T_272; // @[Math.scala 406:56:@32193.4]
  wire  _T_276; // @[FixedPoint.scala 50:25:@32199.4]
  wire [1:0] _T_280; // @[Bitwise.scala 72:12:@32201.4]
  wire [29:0] _T_281; // @[FixedPoint.scala 18:52:@32202.4]
  wire  _T_287; // @[Math.scala 451:55:@32204.4]
  wire [1:0] _T_288; // @[FixedPoint.scala 18:52:@32205.4]
  wire  _T_294; // @[Math.scala 451:110:@32207.4]
  wire  _T_295; // @[Math.scala 451:94:@32208.4]
  wire [31:0] _T_297; // @[Cat.scala 30:58:@32210.4]
  wire [31:0] x308_1_number; // @[Math.scala 454:20:@32211.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@32216.4]
  wire [40:0] _T_302; // @[Math.scala 461:32:@32216.4]
  wire [36:0] _GEN_1; // @[Math.scala 461:32:@32221.4]
  wire [36:0] _T_305; // @[Math.scala 461:32:@32221.4]
  wire  _T_311; // @[FixedPoint.scala 50:25:@32236.4]
  wire [1:0] _T_315; // @[Bitwise.scala 72:12:@32238.4]
  wire [29:0] _T_316; // @[FixedPoint.scala 18:52:@32239.4]
  wire  _T_322; // @[Math.scala 451:55:@32241.4]
  wire [1:0] _T_323; // @[FixedPoint.scala 18:52:@32242.4]
  wire  _T_329; // @[Math.scala 451:110:@32244.4]
  wire  _T_330; // @[Math.scala 451:94:@32245.4]
  wire [31:0] _T_332; // @[Cat.scala 30:58:@32247.4]
  wire  _T_360; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:101:@32324.4]
  wire  _T_364; // @[package.scala 96:25:@32332.4 package.scala 96:25:@32333.4]
  wire  _T_366; // @[implicits.scala 55:10:@32334.4]
  wire  _T_367; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:118:@32335.4]
  wire  _T_369; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:206:@32337.4]
  wire  _T_370; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:225:@32338.4]
  wire  x549_b297_D3; // @[package.scala 96:25:@32276.4 package.scala 96:25:@32277.4]
  wire  _T_371; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:251:@32339.4]
  wire  x551_b298_D3; // @[package.scala 96:25:@32294.4 package.scala 96:25:@32295.4]
  wire [31:0] x313_rdcol_number; // @[Math.scala 154:22:@32356.4 Math.scala 155:14:@32357.4]
  wire [31:0] _T_388; // @[Math.scala 406:49:@32365.4]
  wire [31:0] _T_390; // @[Math.scala 406:56:@32367.4]
  wire [31:0] _T_391; // @[Math.scala 406:56:@32368.4]
  wire  _T_395; // @[FixedPoint.scala 50:25:@32374.4]
  wire [1:0] _T_399; // @[Bitwise.scala 72:12:@32376.4]
  wire [29:0] _T_400; // @[FixedPoint.scala 18:52:@32377.4]
  wire  _T_406; // @[Math.scala 451:55:@32379.4]
  wire [1:0] _T_407; // @[FixedPoint.scala 18:52:@32380.4]
  wire  _T_413; // @[Math.scala 451:110:@32382.4]
  wire  _T_414; // @[Math.scala 451:94:@32383.4]
  wire [31:0] _T_416; // @[Cat.scala 30:58:@32385.4]
  wire  _T_436; // @[package.scala 96:25:@32434.4 package.scala 96:25:@32435.4]
  wire  _T_438; // @[implicits.scala 55:10:@32436.4]
  wire  _T_439; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:118:@32437.4]
  wire  _T_441; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:206:@32439.4]
  wire  _T_442; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:225:@32440.4]
  wire  _T_443; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:251:@32441.4]
  wire [31:0] x558_b295_D6_number; // @[package.scala 96:25:@32455.4 package.scala 96:25:@32456.4]
  wire [31:0] _T_453; // @[Math.scala 476:37:@32461.4]
  wire  x320; // @[Math.scala 476:44:@32463.4]
  wire [31:0] x559_x313_rdcol_D6_number; // @[package.scala 96:25:@32471.4 package.scala 96:25:@32472.4]
  wire [31:0] _T_464; // @[Math.scala 476:37:@32477.4]
  wire  x321; // @[Math.scala 476:44:@32479.4]
  wire  x560_x320_D1; // @[package.scala 96:25:@32487.4 package.scala 96:25:@32488.4]
  wire  x322; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 152:24:@32491.4]
  wire  _T_503; // @[package.scala 96:25:@32559.4 package.scala 96:25:@32560.4]
  wire  _T_505; // @[implicits.scala 55:10:@32561.4]
  wire  _T_506; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 171:146:@32562.4]
  wire  x565_x323_D2; // @[package.scala 96:25:@32538.4 package.scala 96:25:@32539.4]
  wire  _T_507; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 171:234:@32563.4]
  wire  x562_b297_D9; // @[package.scala 96:25:@32511.4 package.scala 96:25:@32512.4]
  wire  _T_508; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 171:242:@32564.4]
  wire  x564_b298_D9; // @[package.scala 96:25:@32529.4 package.scala 96:25:@32530.4]
  wire [31:0] x567_b296_D6_number; // @[package.scala 96:25:@32580.4 package.scala 96:25:@32581.4]
  wire [31:0] _T_521; // @[Math.scala 476:37:@32588.4]
  wire  x326; // @[Math.scala 476:44:@32590.4]
  wire  x327; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 187:59:@32593.4]
  wire  _T_548; // @[package.scala 96:25:@32634.4 package.scala 96:25:@32635.4]
  wire  _T_550; // @[implicits.scala 55:10:@32636.4]
  wire  _T_551; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:194:@32637.4]
  wire  x568_x328_D3; // @[package.scala 96:25:@32604.4 package.scala 96:25:@32605.4]
  wire  _T_552; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:282:@32638.4]
  wire  _T_553; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:290:@32639.4]
  wire [31:0] x331_rdcol_number; // @[Math.scala 154:22:@32658.4 Math.scala 155:14:@32659.4]
  wire [31:0] _T_568; // @[Math.scala 476:37:@32664.4]
  wire  x332; // @[Math.scala 476:44:@32666.4]
  wire  x333; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 208:59:@32669.4]
  wire [31:0] _T_584; // @[Math.scala 406:56:@32680.4]
  wire [31:0] _T_585; // @[Math.scala 406:56:@32681.4]
  wire  _T_589; // @[FixedPoint.scala 50:25:@32687.4]
  wire [1:0] _T_593; // @[Bitwise.scala 72:12:@32689.4]
  wire [29:0] _T_594; // @[FixedPoint.scala 18:52:@32690.4]
  wire  _T_600; // @[Math.scala 451:55:@32692.4]
  wire [1:0] _T_601; // @[FixedPoint.scala 18:52:@32693.4]
  wire  _T_607; // @[Math.scala 451:110:@32695.4]
  wire  _T_608; // @[Math.scala 451:94:@32696.4]
  wire [31:0] _T_610; // @[Cat.scala 30:58:@32698.4]
  wire  _T_639; // @[package.scala 96:25:@32757.4 package.scala 96:25:@32758.4]
  wire  _T_641; // @[implicits.scala 55:10:@32759.4]
  wire  _T_642; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:194:@32760.4]
  wire  x572_x334_D2; // @[package.scala 96:25:@32727.4 package.scala 96:25:@32728.4]
  wire  _T_643; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:282:@32761.4]
  wire  _T_644; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:290:@32762.4]
  wire [31:0] x340_rdcol_number; // @[Math.scala 154:22:@32781.4 Math.scala 155:14:@32782.4]
  wire [31:0] _T_659; // @[Math.scala 476:37:@32787.4]
  wire  x341; // @[Math.scala 476:44:@32789.4]
  wire  x342; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 237:59:@32792.4]
  wire [31:0] _T_675; // @[Math.scala 406:56:@32803.4]
  wire [31:0] _T_676; // @[Math.scala 406:56:@32804.4]
  wire  _T_680; // @[FixedPoint.scala 50:25:@32810.4]
  wire [1:0] _T_684; // @[Bitwise.scala 72:12:@32812.4]
  wire [29:0] _T_685; // @[FixedPoint.scala 18:52:@32813.4]
  wire  _T_691; // @[Math.scala 451:55:@32815.4]
  wire [1:0] _T_692; // @[FixedPoint.scala 18:52:@32816.4]
  wire  _T_698; // @[Math.scala 451:110:@32818.4]
  wire  _T_699; // @[Math.scala 451:94:@32819.4]
  wire [31:0] _T_701; // @[Cat.scala 30:58:@32821.4]
  wire  _T_727; // @[package.scala 96:25:@32871.4 package.scala 96:25:@32872.4]
  wire  _T_729; // @[implicits.scala 55:10:@32873.4]
  wire  _T_730; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 256:194:@32874.4]
  wire  x575_x343_D2; // @[package.scala 96:25:@32841.4 package.scala 96:25:@32842.4]
  wire  _T_731; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 256:282:@32875.4]
  wire  _T_732; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 256:290:@32876.4]
  wire [31:0] x349_rdrow_number; // @[Math.scala 195:22:@32895.4 Math.scala 196:14:@32896.4]
  wire [31:0] _T_749; // @[Math.scala 406:49:@32902.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@32904.4]
  wire [31:0] _T_752; // @[Math.scala 406:56:@32905.4]
  wire [31:0] x532_number; // @[implicits.scala 133:21:@32906.4]
  wire  x351; // @[Math.scala 476:44:@32914.4]
  wire  x352; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 266:24:@32917.4]
  wire [31:0] _T_773; // @[Math.scala 406:49:@32926.4]
  wire [31:0] _T_775; // @[Math.scala 406:56:@32928.4]
  wire [31:0] _T_776; // @[Math.scala 406:56:@32929.4]
  wire  _T_780; // @[FixedPoint.scala 50:25:@32935.4]
  wire [1:0] _T_784; // @[Bitwise.scala 72:12:@32937.4]
  wire [29:0] _T_785; // @[FixedPoint.scala 18:52:@32938.4]
  wire  _T_791; // @[Math.scala 451:55:@32940.4]
  wire [1:0] _T_792; // @[FixedPoint.scala 18:52:@32941.4]
  wire  _T_798; // @[Math.scala 451:110:@32943.4]
  wire  _T_799; // @[Math.scala 451:94:@32944.4]
  wire [31:0] _T_801; // @[Cat.scala 30:58:@32946.4]
  wire [31:0] x355_1_number; // @[Math.scala 454:20:@32947.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@32952.4]
  wire [40:0] _T_806; // @[Math.scala 461:32:@32952.4]
  wire [36:0] _GEN_3; // @[Math.scala 461:32:@32957.4]
  wire [36:0] _T_809; // @[Math.scala 461:32:@32957.4]
  wire  _T_836; // @[package.scala 96:25:@33016.4 package.scala 96:25:@33017.4]
  wire  _T_838; // @[implicits.scala 55:10:@33018.4]
  wire  _T_839; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:194:@33019.4]
  wire  x580_x353_D2; // @[package.scala 96:25:@33004.4 package.scala 96:25:@33005.4]
  wire  _T_840; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:282:@33020.4]
  wire  _T_841; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:290:@33021.4]
  wire  x581_x326_D1; // @[package.scala 96:25:@33037.4 package.scala 96:25:@33038.4]
  wire  x360; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 303:59:@33041.4]
  wire  _T_873; // @[package.scala 96:25:@33085.4 package.scala 96:25:@33086.4]
  wire  _T_875; // @[implicits.scala 55:10:@33087.4]
  wire  _T_876; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:194:@33088.4]
  wire  x583_x361_D2; // @[package.scala 96:25:@33073.4 package.scala 96:25:@33074.4]
  wire  _T_877; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:282:@33089.4]
  wire  _T_878; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:290:@33090.4]
  wire  x365; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 322:59:@33101.4]
  wire  _T_905; // @[package.scala 96:25:@33143.4 package.scala 96:25:@33144.4]
  wire  _T_907; // @[implicits.scala 55:10:@33145.4]
  wire  _T_908; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:194:@33146.4]
  wire  x585_x366_D2; // @[package.scala 96:25:@33131.4 package.scala 96:25:@33132.4]
  wire  _T_909; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:282:@33147.4]
  wire  _T_910; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:290:@33148.4]
  wire  x370; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 339:59:@33159.4]
  wire  _T_937; // @[package.scala 96:25:@33201.4 package.scala 96:25:@33202.4]
  wire  _T_939; // @[implicits.scala 55:10:@33203.4]
  wire  _T_940; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:194:@33204.4]
  wire  x587_x371_D2; // @[package.scala 96:25:@33189.4 package.scala 96:25:@33190.4]
  wire  _T_941; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:282:@33205.4]
  wire  _T_942; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:290:@33206.4]
  wire [31:0] x375_rdrow_number; // @[Math.scala 195:22:@33225.4 Math.scala 196:14:@33226.4]
  wire [31:0] _T_959; // @[Math.scala 406:49:@33232.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@33234.4]
  wire [31:0] _T_962; // @[Math.scala 406:56:@33235.4]
  wire [31:0] x537_number; // @[implicits.scala 133:21:@33236.4]
  wire  x377; // @[Math.scala 476:44:@33244.4]
  wire  x378; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 362:24:@33247.4]
  wire [31:0] _T_983; // @[Math.scala 406:49:@33256.4]
  wire [31:0] _T_985; // @[Math.scala 406:56:@33258.4]
  wire [31:0] _T_986; // @[Math.scala 406:56:@33259.4]
  wire  _T_990; // @[FixedPoint.scala 50:25:@33265.4]
  wire [1:0] _T_994; // @[Bitwise.scala 72:12:@33267.4]
  wire [29:0] _T_995; // @[FixedPoint.scala 18:52:@33268.4]
  wire  _T_1001; // @[Math.scala 451:55:@33270.4]
  wire [1:0] _T_1002; // @[FixedPoint.scala 18:52:@33271.4]
  wire  _T_1008; // @[Math.scala 451:110:@33273.4]
  wire  _T_1009; // @[Math.scala 451:94:@33274.4]
  wire [31:0] _T_1011; // @[Cat.scala 30:58:@33276.4]
  wire [31:0] x381_1_number; // @[Math.scala 454:20:@33277.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@33282.4]
  wire [40:0] _T_1016; // @[Math.scala 461:32:@33282.4]
  wire [36:0] _GEN_5; // @[Math.scala 461:32:@33287.4]
  wire [36:0] _T_1019; // @[Math.scala 461:32:@33287.4]
  wire  _T_1043; // @[package.scala 96:25:@33337.4 package.scala 96:25:@33338.4]
  wire  _T_1045; // @[implicits.scala 55:10:@33339.4]
  wire  _T_1046; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 385:194:@33340.4]
  wire  x588_x379_D2; // @[package.scala 96:25:@33316.4 package.scala 96:25:@33317.4]
  wire  _T_1047; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 385:282:@33341.4]
  wire  _T_1048; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 385:290:@33342.4]
  wire  x386; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 389:24:@33353.4]
  wire  _T_1072; // @[package.scala 96:25:@33386.4 package.scala 96:25:@33387.4]
  wire  _T_1074; // @[implicits.scala 55:10:@33388.4]
  wire  _T_1075; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:194:@33389.4]
  wire  x590_x387_D2; // @[package.scala 96:25:@33374.4 package.scala 96:25:@33375.4]
  wire  _T_1076; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:282:@33390.4]
  wire  _T_1077; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:290:@33391.4]
  wire  x391; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 404:24:@33402.4]
  wire  _T_1101; // @[package.scala 96:25:@33435.4 package.scala 96:25:@33436.4]
  wire  _T_1103; // @[implicits.scala 55:10:@33437.4]
  wire  _T_1104; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:194:@33438.4]
  wire  x591_x392_D2; // @[package.scala 96:25:@33423.4 package.scala 96:25:@33424.4]
  wire  _T_1105; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:282:@33439.4]
  wire  _T_1106; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:290:@33440.4]
  wire  x396; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 425:59:@33451.4]
  wire  _T_1132; // @[package.scala 96:25:@33486.4 package.scala 96:25:@33487.4]
  wire  _T_1134; // @[implicits.scala 55:10:@33488.4]
  wire  _T_1135; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 438:194:@33489.4]
  wire  x592_x397_D2; // @[package.scala 96:25:@33474.4 package.scala 96:25:@33475.4]
  wire  _T_1136; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 438:282:@33490.4]
  wire  _T_1137; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 438:290:@33491.4]
  wire [31:0] x329_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 196:29:@32625.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:407:@32646.4]
  wire [32:0] _GEN_6; // @[Math.scala 461:32:@33503.4]
  wire [31:0] x358_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 287:29:@33007.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:407:@33028.4]
  wire [32:0] _GEN_7; // @[Math.scala 461:32:@33515.4]
  wire [31:0] x363_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 314:29:@33076.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:407:@33097.4]
  wire [33:0] _GEN_8; // @[Math.scala 461:32:@33527.4]
  wire [31:0] x368_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 331:29:@33134.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:407:@33155.4]
  wire [32:0] _GEN_9; // @[Math.scala 461:32:@33539.4]
  wire [31:0] x389_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 396:29:@33377.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:407:@33398.4]
  wire [32:0] _GEN_10; // @[Math.scala 461:32:@33551.4]
  wire [31:0] x338_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 225:29:@32748.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:407:@32769.4]
  wire [32:0] _GEN_11; // @[Math.scala 461:32:@33709.4]
  wire [32:0] _GEN_12; // @[Math.scala 461:32:@33721.4]
  wire [33:0] _GEN_13; // @[Math.scala 461:32:@33733.4]
  wire [31:0] x373_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 348:29:@33192.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:407:@33213.4]
  wire [32:0] _GEN_14; // @[Math.scala 461:32:@33745.4]
  wire [31:0] x394_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 411:29:@33426.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:407:@33447.4]
  wire [32:0] _GEN_15; // @[Math.scala 461:32:@33757.4]
  wire  _T_1311; // @[package.scala 96:25:@33975.4 package.scala 96:25:@33976.4]
  wire  _T_1313; // @[implicits.scala 55:10:@33977.4]
  wire  _T_1314; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:167:@33978.4]
  wire  _T_1316; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:256:@33980.4]
  wire  _T_1317; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:275:@33981.4]
  wire  x601_b297_D23; // @[package.scala 96:25:@33919.4 package.scala 96:25:@33920.4]
  wire  _T_1318; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:301:@33982.4]
  wire  x603_b298_D23; // @[package.scala 96:25:@33937.4 package.scala 96:25:@33938.4]
  wire  _T_1334; // @[package.scala 96:25:@34025.4 package.scala 96:25:@34026.4]
  wire  _T_1336; // @[implicits.scala 55:10:@34027.4]
  wire  _T_1337; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:167:@34028.4]
  wire  _T_1339; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:256:@34030.4]
  wire  _T_1340; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:275:@34031.4]
  wire  _T_1341; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:301:@34032.4]
  wire  _T_1372; // @[package.scala 96:25:@34103.4 package.scala 96:25:@34104.4]
  wire  _T_1374; // @[implicits.scala 55:10:@34105.4]
  wire  _T_1375; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 573:195:@34106.4]
  wire  x614_x323_D17; // @[package.scala 96:25:@34082.4 package.scala 96:25:@34083.4]
  wire  _T_1376; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 573:284:@34107.4]
  wire  x611_b297_D24; // @[package.scala 96:25:@34055.4 package.scala 96:25:@34056.4]
  wire  _T_1377; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 573:292:@34108.4]
  wire  x613_b298_D24; // @[package.scala 96:25:@34073.4 package.scala 96:25:@34074.4]
  wire  _T_1400; // @[package.scala 96:25:@34154.4 package.scala 96:25:@34155.4]
  wire  _T_1402; // @[implicits.scala 55:10:@34156.4]
  wire  _T_1403; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:195:@34157.4]
  wire  x616_x328_D18; // @[package.scala 96:25:@34124.4 package.scala 96:25:@34125.4]
  wire  _T_1404; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:284:@34158.4]
  wire  _T_1405; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:292:@34159.4]
  wire  _T_1428; // @[package.scala 96:25:@34205.4 package.scala 96:25:@34206.4]
  wire  _T_1430; // @[implicits.scala 55:10:@34207.4]
  wire  _T_1431; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:195:@34208.4]
  wire  x619_x334_D17; // @[package.scala 96:25:@34175.4 package.scala 96:25:@34176.4]
  wire  _T_1432; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:284:@34209.4]
  wire  _T_1433; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:292:@34210.4]
  wire  _T_1456; // @[package.scala 96:25:@34256.4 package.scala 96:25:@34257.4]
  wire  _T_1458; // @[implicits.scala 55:10:@34258.4]
  wire  _T_1459; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:195:@34259.4]
  wire  x624_x353_D17; // @[package.scala 96:25:@34244.4 package.scala 96:25:@34245.4]
  wire  _T_1460; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:284:@34260.4]
  wire  _T_1461; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:292:@34261.4]
  wire  _T_1481; // @[package.scala 96:25:@34298.4 package.scala 96:25:@34299.4]
  wire  _T_1483; // @[implicits.scala 55:10:@34300.4]
  wire  _T_1484; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:195:@34301.4]
  wire  x625_x361_D17; // @[package.scala 96:25:@34277.4 package.scala 96:25:@34278.4]
  wire  _T_1485; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:284:@34302.4]
  wire  _T_1486; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:292:@34303.4]
  wire  _T_1506; // @[package.scala 96:25:@34340.4 package.scala 96:25:@34341.4]
  wire  _T_1508; // @[implicits.scala 55:10:@34342.4]
  wire  _T_1509; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 634:195:@34343.4]
  wire  x627_x366_D17; // @[package.scala 96:25:@34319.4 package.scala 96:25:@34320.4]
  wire  _T_1510; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 634:284:@34344.4]
  wire  _T_1511; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 634:292:@34345.4]
  wire [31:0] x439_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 582:29:@34145.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:339:@34166.4]
  wire [32:0] _GEN_16; // @[Math.scala 461:32:@34359.4]
  wire [32:0] _T_1518; // @[Math.scala 461:32:@34359.4]
  wire [31:0] x443_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 608:29:@34247.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:339:@34268.4]
  wire [33:0] _GEN_17; // @[Math.scala 461:32:@34364.4]
  wire [33:0] _T_1521; // @[Math.scala 461:32:@34364.4]
  wire [31:0] x441_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 595:29:@34196.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:339:@34217.4]
  wire [32:0] _GEN_18; // @[Math.scala 461:32:@34431.4]
  wire [32:0] _T_1548; // @[Math.scala 461:32:@34431.4]
  wire [31:0] x445_rd_0_number; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 619:29:@34289.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:339:@34310.4]
  wire [33:0] _GEN_19; // @[Math.scala 461:32:@34436.4]
  wire [33:0] _T_1551; // @[Math.scala 461:32:@34436.4]
  wire [31:0] x456_number; // @[Math.scala 723:22:@34426.4 Math.scala 724:14:@34427.4]
  wire [31:0] x464_number; // @[Math.scala 723:22:@34496.4 Math.scala 724:14:@34497.4]
  wire  _T_1595; // @[package.scala 96:25:@34538.4 package.scala 96:25:@34539.4]
  wire  _T_1597; // @[implicits.scala 55:10:@34540.4]
  wire  x630_b297_D37; // @[package.scala 96:25:@34529.4 package.scala 96:25:@34530.4]
  wire  _T_1598; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 688:117:@34541.4]
  wire  x629_b298_D37; // @[package.scala 96:25:@34520.4 package.scala 96:25:@34521.4]
  wire  _T_1599; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 688:123:@34542.4]
  wire [31:0] x550_x311_sum_D1_number; // @[package.scala 96:25:@32285.4 package.scala 96:25:@32286.4]
  wire [31:0] x552_x525_D3_number; // @[package.scala 96:25:@32303.4 package.scala 96:25:@32304.4]
  wire [31:0] x553_x524_D3_number; // @[package.scala 96:25:@32312.4 package.scala 96:25:@32313.4]
  wire [31:0] x555_x529_D2_number; // @[package.scala 96:25:@32405.4 package.scala 96:25:@32406.4]
  wire [31:0] x556_x317_sum_D1_number; // @[package.scala 96:25:@32414.4 package.scala 96:25:@32415.4]
  wire [31:0] x561_x529_D8_number; // @[package.scala 96:25:@32502.4 package.scala 96:25:@32503.4]
  wire [31:0] x563_x317_sum_D7_number; // @[package.scala 96:25:@32520.4 package.scala 96:25:@32521.4]
  wire [31:0] x566_x524_D9_number; // @[package.scala 96:25:@32547.4 package.scala 96:25:@32548.4]
  wire [31:0] x569_x311_sum_D7_number; // @[package.scala 96:25:@32613.4 package.scala 96:25:@32614.4]
  wire [31:0] x570_x525_D9_number; // @[package.scala 96:25:@32622.4 package.scala 96:25:@32623.4]
  wire [31:0] x573_x530_D2_number; // @[package.scala 96:25:@32736.4 package.scala 96:25:@32737.4]
  wire [31:0] x574_x337_sum_D1_number; // @[package.scala 96:25:@32745.4 package.scala 96:25:@32746.4]
  wire [31:0] x576_x531_D2_number; // @[package.scala 96:25:@32850.4 package.scala 96:25:@32851.4]
  wire [31:0] x577_x346_sum_D1_number; // @[package.scala 96:25:@32859.4 package.scala 96:25:@32860.4]
  wire [31:0] x357_sum_number; // @[Math.scala 154:22:@32986.4 Math.scala 155:14:@32987.4]
  wire [31:0] x579_x533_D2_number; // @[package.scala 96:25:@32995.4 package.scala 96:25:@32996.4]
  wire [31:0] x362_sum_number; // @[Math.scala 154:22:@33064.4 Math.scala 155:14:@33065.4]
  wire [31:0] x367_sum_number; // @[Math.scala 154:22:@33122.4 Math.scala 155:14:@33123.4]
  wire [31:0] x372_sum_number; // @[Math.scala 154:22:@33180.4 Math.scala 155:14:@33181.4]
  wire [31:0] x383_sum_number; // @[Math.scala 154:22:@33307.4 Math.scala 155:14:@33308.4]
  wire [31:0] x589_x538_D2_number; // @[package.scala 96:25:@33325.4 package.scala 96:25:@33326.4]
  wire [31:0] x388_sum_number; // @[Math.scala 154:22:@33365.4 Math.scala 155:14:@33366.4]
  wire [31:0] x393_sum_number; // @[Math.scala 154:22:@33414.4 Math.scala 155:14:@33415.4]
  wire [31:0] x398_sum_number; // @[Math.scala 154:22:@33465.4 Math.scala 155:14:@33466.4]
  wire [32:0] _T_1144; // @[package.scala 96:25:@33509.4 package.scala 96:25:@33510.4]
  wire [32:0] _T_1149; // @[package.scala 96:25:@33521.4 package.scala 96:25:@33522.4]
  wire [33:0] _T_1154; // @[package.scala 96:25:@33533.4 package.scala 96:25:@33534.4]
  wire [32:0] _T_1159; // @[package.scala 96:25:@33545.4 package.scala 96:25:@33546.4]
  wire [32:0] _T_1164; // @[package.scala 96:25:@33557.4 package.scala 96:25:@33558.4]
  wire [32:0] _T_1218; // @[package.scala 96:25:@33715.4 package.scala 96:25:@33716.4]
  wire [32:0] _T_1223; // @[package.scala 96:25:@33727.4 package.scala 96:25:@33728.4]
  wire [33:0] _T_1228; // @[package.scala 96:25:@33739.4 package.scala 96:25:@33740.4]
  wire [32:0] _T_1233; // @[package.scala 96:25:@33751.4 package.scala 96:25:@33752.4]
  wire [32:0] _T_1238; // @[package.scala 96:25:@33763.4 package.scala 96:25:@33764.4]
  wire [31:0] x602_x311_sum_D21_number; // @[package.scala 96:25:@33928.4 package.scala 96:25:@33929.4]
  wire [31:0] x604_x525_D23_number; // @[package.scala 96:25:@33946.4 package.scala 96:25:@33947.4]
  wire [31:0] x605_x524_D23_number; // @[package.scala 96:25:@33955.4 package.scala 96:25:@33956.4]
  wire [31:0] x608_x529_D22_number; // @[package.scala 96:25:@34005.4 package.scala 96:25:@34006.4]
  wire [31:0] x609_x317_sum_D21_number; // @[package.scala 96:25:@34014.4 package.scala 96:25:@34015.4]
  wire [31:0] x610_x529_D23_number; // @[package.scala 96:25:@34046.4 package.scala 96:25:@34047.4]
  wire [31:0] x612_x317_sum_D22_number; // @[package.scala 96:25:@34064.4 package.scala 96:25:@34065.4]
  wire [31:0] x615_x524_D24_number; // @[package.scala 96:25:@34091.4 package.scala 96:25:@34092.4]
  wire [31:0] x617_x311_sum_D22_number; // @[package.scala 96:25:@34133.4 package.scala 96:25:@34134.4]
  wire [31:0] x618_x525_D24_number; // @[package.scala 96:25:@34142.4 package.scala 96:25:@34143.4]
  wire [31:0] x620_x530_D17_number; // @[package.scala 96:25:@34184.4 package.scala 96:25:@34185.4]
  wire [31:0] x621_x337_sum_D16_number; // @[package.scala 96:25:@34193.4 package.scala 96:25:@34194.4]
  wire [31:0] x622_x533_D17_number; // @[package.scala 96:25:@34226.4 package.scala 96:25:@34227.4]
  wire [31:0] x623_x357_sum_D15_number; // @[package.scala 96:25:@34235.4 package.scala 96:25:@34236.4]
  wire [31:0] x626_x362_sum_D15_number; // @[package.scala 96:25:@34286.4 package.scala 96:25:@34287.4]
  wire [31:0] x628_x367_sum_D15_number; // @[package.scala 96:25:@34328.4 package.scala 96:25:@34329.4]
  _ _ ( // @[Math.scala 720:24:@31960.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@31972.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@31995.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x301_lb_0 x301_lb_0 ( // @[m_x301_lb_0.scala 39:17:@32005.4]
    .clock(x301_lb_0_clock),
    .reset(x301_lb_0_reset),
    .io_rPort_11_banks_1(x301_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x301_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x301_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x301_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x301_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x301_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x301_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x301_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x301_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x301_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x301_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x301_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x301_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x301_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x301_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x301_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x301_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x301_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x301_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x301_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x301_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x301_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x301_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x301_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x301_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x301_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x301_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x301_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x301_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x301_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x301_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x301_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x301_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x301_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x301_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x301_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x301_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x301_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x301_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x301_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x301_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x301_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x301_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x301_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x301_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x301_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x301_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x301_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x301_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x301_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x301_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x301_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x301_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x301_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x301_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x301_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x301_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x301_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x301_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x301_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x301_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x301_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x301_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x301_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x301_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x301_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x301_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x301_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x301_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x301_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x301_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x301_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x301_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x301_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x301_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x301_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x301_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x301_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x301_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x301_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x301_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x301_lb_0_io_wPort_0_en_0)
  );
  x302_lb2_0 x302_lb2_0 ( // @[m_x302_lb2_0.scala 33:17:@32098.4]
    .clock(x302_lb2_0_clock),
    .reset(x302_lb2_0_reset),
    .io_rPort_5_banks_1(x302_lb2_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x302_lb2_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x302_lb2_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x302_lb2_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x302_lb2_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x302_lb2_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x302_lb2_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x302_lb2_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x302_lb2_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x302_lb2_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x302_lb2_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x302_lb2_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x302_lb2_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x302_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x302_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x302_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x302_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x302_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x302_lb2_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x302_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x302_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x302_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x302_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x302_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x302_lb2_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x302_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x302_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x302_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x302_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x302_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x302_lb2_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x302_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x302_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x302_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x302_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x302_lb2_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x302_lb2_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x302_lb2_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x302_lb2_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x302_lb2_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x302_lb2_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x302_lb2_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x302_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x302_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x302_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x302_lb2_0_io_wPort_0_en_0)
  );
  x520_sub x528_sub_1 ( // @[Math.scala 191:24:@32225.4]
    .clock(x528_sub_1_clock),
    .reset(x528_sub_1_reset),
    .io_a(x528_sub_1_io_a),
    .io_b(x528_sub_1_io_b),
    .io_flow(x528_sub_1_io_flow),
    .io_result(x528_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@32252.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x280_sum x311_sum_1 ( // @[Math.scala 150:24:@32261.4]
    .clock(x311_sum_1_clock),
    .reset(x311_sum_1_reset),
    .io_a(x311_sum_1_io_a),
    .io_b(x311_sum_1_io_b),
    .io_flow(x311_sum_1_io_flow),
    .io_result(x311_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@32271.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_3 ( // @[package.scala 93:22:@32280.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@32289.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_233 RetimeWrapper_5 ( // @[package.scala 93:22:@32298.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_233 RetimeWrapper_6 ( // @[package.scala 93:22:@32307.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_235 RetimeWrapper_7 ( // @[package.scala 93:22:@32316.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_8 ( // @[package.scala 93:22:@32327.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x280_sum x313_rdcol_1 ( // @[Math.scala 150:24:@32350.4]
    .clock(x313_rdcol_1_clock),
    .reset(x313_rdcol_1_reset),
    .io_a(x313_rdcol_1_io_a),
    .io_b(x313_rdcol_1_io_b),
    .io_flow(x313_rdcol_1_io_flow),
    .io_result(x313_rdcol_1_io_result)
  );
  x280_sum x317_sum_1 ( // @[Math.scala 150:24:@32390.4]
    .clock(x317_sum_1_clock),
    .reset(x317_sum_1_reset),
    .io_a(x317_sum_1_io_a),
    .io_b(x317_sum_1_io_b),
    .io_flow(x317_sum_1_io_flow),
    .io_result(x317_sum_1_io_result)
  );
  RetimeWrapper_235 RetimeWrapper_9 ( // @[package.scala 93:22:@32400.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_10 ( // @[package.scala 93:22:@32409.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_235 RetimeWrapper_11 ( // @[package.scala 93:22:@32418.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_12 ( // @[package.scala 93:22:@32429.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_13 ( // @[package.scala 93:22:@32450.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_14 ( // @[package.scala 93:22:@32466.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@32482.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_16 ( // @[package.scala 93:22:@32497.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_17 ( // @[package.scala 93:22:@32506.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_18 ( // @[package.scala 93:22:@32515.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_19 ( // @[package.scala 93:22:@32524.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@32533.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_251 RetimeWrapper_21 ( // @[package.scala 93:22:@32542.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_22 ( // @[package.scala 93:22:@32554.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_23 ( // @[package.scala 93:22:@32575.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_24 ( // @[package.scala 93:22:@32599.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_25 ( // @[package.scala 93:22:@32608.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_251 RetimeWrapper_26 ( // @[package.scala 93:22:@32617.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_27 ( // @[package.scala 93:22:@32629.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x280_sum x331_rdcol_1 ( // @[Math.scala 150:24:@32652.4]
    .clock(x331_rdcol_1_clock),
    .reset(x331_rdcol_1_reset),
    .io_a(x331_rdcol_1_io_a),
    .io_b(x331_rdcol_1_io_b),
    .io_flow(x331_rdcol_1_io_flow),
    .io_result(x331_rdcol_1_io_result)
  );
  RetimeWrapper_243 RetimeWrapper_28 ( // @[package.scala 93:22:@32703.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x280_sum x337_sum_1 ( // @[Math.scala 150:24:@32712.4]
    .clock(x337_sum_1_clock),
    .reset(x337_sum_1_reset),
    .io_a(x337_sum_1_io_a),
    .io_b(x337_sum_1_io_b),
    .io_flow(x337_sum_1_io_flow),
    .io_result(x337_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@32722.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_235 RetimeWrapper_30 ( // @[package.scala 93:22:@32731.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_31 ( // @[package.scala 93:22:@32740.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_32 ( // @[package.scala 93:22:@32752.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x280_sum x340_rdcol_1 ( // @[Math.scala 150:24:@32775.4]
    .clock(x340_rdcol_1_clock),
    .reset(x340_rdcol_1_reset),
    .io_a(x340_rdcol_1_io_a),
    .io_b(x340_rdcol_1_io_b),
    .io_flow(x340_rdcol_1_io_flow),
    .io_result(x340_rdcol_1_io_result)
  );
  x280_sum x346_sum_1 ( // @[Math.scala 150:24:@32826.4]
    .clock(x346_sum_1_clock),
    .reset(x346_sum_1_reset),
    .io_a(x346_sum_1_io_a),
    .io_b(x346_sum_1_io_b),
    .io_flow(x346_sum_1_io_flow),
    .io_result(x346_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@32836.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_235 RetimeWrapper_34 ( // @[package.scala 93:22:@32845.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_35 ( // @[package.scala 93:22:@32854.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_36 ( // @[package.scala 93:22:@32866.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x520_sub x349_rdrow_1 ( // @[Math.scala 191:24:@32889.4]
    .clock(x349_rdrow_1_clock),
    .reset(x349_rdrow_1_reset),
    .io_a(x349_rdrow_1_io_a),
    .io_b(x349_rdrow_1_io_b),
    .io_flow(x349_rdrow_1_io_flow),
    .io_result(x349_rdrow_1_io_result)
  );
  x520_sub x536_sub_1 ( // @[Math.scala 191:24:@32961.4]
    .clock(x536_sub_1_clock),
    .reset(x536_sub_1_reset),
    .io_a(x536_sub_1_io_a),
    .io_b(x536_sub_1_io_b),
    .io_flow(x536_sub_1_io_flow),
    .io_result(x536_sub_1_io_result)
  );
  RetimeWrapper_248 RetimeWrapper_37 ( // @[package.scala 93:22:@32971.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x280_sum x357_sum_1 ( // @[Math.scala 150:24:@32980.4]
    .clock(x357_sum_1_clock),
    .reset(x357_sum_1_reset),
    .io_a(x357_sum_1_io_a),
    .io_b(x357_sum_1_io_b),
    .io_flow(x357_sum_1_io_flow),
    .io_result(x357_sum_1_io_result)
  );
  RetimeWrapper_235 RetimeWrapper_38 ( // @[package.scala 93:22:@32990.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@32999.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_40 ( // @[package.scala 93:22:@33011.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@33032.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_42 ( // @[package.scala 93:22:@33047.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  x280_sum x362_sum_1 ( // @[Math.scala 150:24:@33058.4]
    .clock(x362_sum_1_clock),
    .reset(x362_sum_1_reset),
    .io_a(x362_sum_1_io_a),
    .io_b(x362_sum_1_io_b),
    .io_flow(x362_sum_1_io_flow),
    .io_result(x362_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@33068.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_44 ( // @[package.scala 93:22:@33080.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_45 ( // @[package.scala 93:22:@33107.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x280_sum x367_sum_1 ( // @[Math.scala 150:24:@33116.4]
    .clock(x367_sum_1_clock),
    .reset(x367_sum_1_reset),
    .io_a(x367_sum_1_io_a),
    .io_b(x367_sum_1_io_b),
    .io_flow(x367_sum_1_io_flow),
    .io_result(x367_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@33126.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_47 ( // @[package.scala 93:22:@33138.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_48 ( // @[package.scala 93:22:@33165.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x280_sum x372_sum_1 ( // @[Math.scala 150:24:@33174.4]
    .clock(x372_sum_1_clock),
    .reset(x372_sum_1_reset),
    .io_a(x372_sum_1_io_a),
    .io_b(x372_sum_1_io_b),
    .io_flow(x372_sum_1_io_flow),
    .io_result(x372_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@33184.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_50 ( // @[package.scala 93:22:@33196.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x520_sub x375_rdrow_1 ( // @[Math.scala 191:24:@33219.4]
    .clock(x375_rdrow_1_clock),
    .reset(x375_rdrow_1_reset),
    .io_a(x375_rdrow_1_io_a),
    .io_b(x375_rdrow_1_io_b),
    .io_flow(x375_rdrow_1_io_flow),
    .io_result(x375_rdrow_1_io_result)
  );
  x520_sub x541_sub_1 ( // @[Math.scala 191:24:@33291.4]
    .clock(x541_sub_1_clock),
    .reset(x541_sub_1_reset),
    .io_a(x541_sub_1_io_a),
    .io_b(x541_sub_1_io_b),
    .io_flow(x541_sub_1_io_flow),
    .io_result(x541_sub_1_io_result)
  );
  x280_sum x383_sum_1 ( // @[Math.scala 150:24:@33301.4]
    .clock(x383_sum_1_clock),
    .reset(x383_sum_1_reset),
    .io_a(x383_sum_1_io_a),
    .io_b(x383_sum_1_io_b),
    .io_flow(x383_sum_1_io_flow),
    .io_result(x383_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@33311.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_235 RetimeWrapper_52 ( // @[package.scala 93:22:@33320.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_53 ( // @[package.scala 93:22:@33332.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x280_sum x388_sum_1 ( // @[Math.scala 150:24:@33359.4]
    .clock(x388_sum_1_clock),
    .reset(x388_sum_1_reset),
    .io_a(x388_sum_1_io_a),
    .io_b(x388_sum_1_io_b),
    .io_flow(x388_sum_1_io_flow),
    .io_result(x388_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@33369.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_55 ( // @[package.scala 93:22:@33381.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x280_sum x393_sum_1 ( // @[Math.scala 150:24:@33408.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@33418.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_57 ( // @[package.scala 93:22:@33430.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x280_sum x398_sum_1 ( // @[Math.scala 150:24:@33459.4]
    .clock(x398_sum_1_clock),
    .reset(x398_sum_1_reset),
    .io_a(x398_sum_1_io_a),
    .io_b(x398_sum_1_io_b),
    .io_flow(x398_sum_1_io_flow),
    .io_result(x398_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@33469.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_247 RetimeWrapper_59 ( // @[package.scala 93:22:@33481.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_60 ( // @[package.scala 93:22:@33504.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_61 ( // @[package.scala 93:22:@33516.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_62 ( // @[package.scala 93:22:@33528.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_63 ( // @[package.scala 93:22:@33540.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_64 ( // @[package.scala 93:22:@33552.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_65 ( // @[package.scala 93:22:@33562.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x406_x7 x406_x7_1 ( // @[Math.scala 150:24:@33571.4]
    .clock(x406_x7_1_clock),
    .reset(x406_x7_1_reset),
    .io_a(x406_x7_1_io_a),
    .io_b(x406_x7_1_io_b),
    .io_flow(x406_x7_1_io_flow),
    .io_result(x406_x7_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_66 ( // @[package.scala 93:22:@33581.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x406_x7 x407_x8_1 ( // @[Math.scala 150:24:@33590.4]
    .clock(x407_x8_1_clock),
    .reset(x407_x8_1_reset),
    .io_a(x407_x8_1_io_a),
    .io_b(x407_x8_1_io_b),
    .io_flow(x407_x8_1_io_flow),
    .io_result(x407_x8_1_io_result)
  );
  x406_x7 x408_x7_1 ( // @[Math.scala 150:24:@33600.4]
    .clock(x408_x7_1_clock),
    .reset(x408_x7_1_reset),
    .io_a(x408_x7_1_io_a),
    .io_b(x408_x7_1_io_b),
    .io_flow(x408_x7_1_io_flow),
    .io_result(x408_x7_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_67 ( // @[package.scala 93:22:@33610.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x406_x7 x409_x8_1 ( // @[Math.scala 150:24:@33619.4]
    .clock(x409_x8_1_clock),
    .reset(x409_x8_1_reset),
    .io_a(x409_x8_1_io_a),
    .io_b(x409_x8_1_io_b),
    .io_flow(x409_x8_1_io_flow),
    .io_result(x409_x8_1_io_result)
  );
  x406_x7 x410_x7_1 ( // @[Math.scala 150:24:@33629.4]
    .clock(x410_x7_1_clock),
    .reset(x410_x7_1_reset),
    .io_a(x410_x7_1_io_a),
    .io_b(x410_x7_1_io_b),
    .io_flow(x410_x7_1_io_flow),
    .io_result(x410_x7_1_io_result)
  );
  x406_x7 x411_x8_1 ( // @[Math.scala 150:24:@33639.4]
    .clock(x411_x8_1_clock),
    .reset(x411_x8_1_reset),
    .io_a(x411_x8_1_io_a),
    .io_b(x411_x8_1_io_b),
    .io_flow(x411_x8_1_io_flow),
    .io_result(x411_x8_1_io_result)
  );
  x406_x7 x412_x7_1 ( // @[Math.scala 150:24:@33649.4]
    .clock(x412_x7_1_clock),
    .reset(x412_x7_1_reset),
    .io_a(x412_x7_1_io_a),
    .io_b(x412_x7_1_io_b),
    .io_flow(x412_x7_1_io_flow),
    .io_result(x412_x7_1_io_result)
  );
  RetimeWrapper_321 RetimeWrapper_68 ( // @[package.scala 93:22:@33659.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  x406_x7 x413_sum_1 ( // @[Math.scala 150:24:@33668.4]
    .clock(x413_sum_1_clock),
    .reset(x413_sum_1_reset),
    .io_a(x413_sum_1_io_a),
    .io_b(x413_sum_1_io_b),
    .io_flow(x413_sum_1_io_flow),
    .io_result(x413_sum_1_io_result)
  );
  x414 x414_1 ( // @[Math.scala 720:24:@33678.4]
    .io_b(x414_1_io_b),
    .io_result(x414_1_io_result)
  );
  x415_mul x415_mul_1 ( // @[Math.scala 262:24:@33689.4]
    .clock(x415_mul_1_clock),
    .io_a(x415_mul_1_io_a),
    .io_b(x415_mul_1_io_b),
    .io_flow(x415_mul_1_io_flow),
    .io_result(x415_mul_1_io_result)
  );
  x416 x416_1 ( // @[Math.scala 720:24:@33699.4]
    .io_b(x416_1_io_b),
    .io_result(x416_1_io_result)
  );
  RetimeWrapper_306 RetimeWrapper_69 ( // @[package.scala 93:22:@33710.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_70 ( // @[package.scala 93:22:@33722.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_308 RetimeWrapper_71 ( // @[package.scala 93:22:@33734.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_72 ( // @[package.scala 93:22:@33746.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_306 RetimeWrapper_73 ( // @[package.scala 93:22:@33758.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_74 ( // @[package.scala 93:22:@33768.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x406_x7 x422_x7_1 ( // @[Math.scala 150:24:@33777.4]
    .clock(x422_x7_1_clock),
    .reset(x422_x7_1_reset),
    .io_a(x422_x7_1_io_a),
    .io_b(x422_x7_1_io_b),
    .io_flow(x422_x7_1_io_flow),
    .io_result(x422_x7_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_75 ( // @[package.scala 93:22:@33787.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  x406_x7 x423_x8_1 ( // @[Math.scala 150:24:@33796.4]
    .clock(x423_x8_1_clock),
    .reset(x423_x8_1_reset),
    .io_a(x423_x8_1_io_a),
    .io_b(x423_x8_1_io_b),
    .io_flow(x423_x8_1_io_flow),
    .io_result(x423_x8_1_io_result)
  );
  x406_x7 x424_x7_1 ( // @[Math.scala 150:24:@33806.4]
    .clock(x424_x7_1_clock),
    .reset(x424_x7_1_reset),
    .io_a(x424_x7_1_io_a),
    .io_b(x424_x7_1_io_b),
    .io_flow(x424_x7_1_io_flow),
    .io_result(x424_x7_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_76 ( // @[package.scala 93:22:@33816.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x406_x7 x425_x8_1 ( // @[Math.scala 150:24:@33825.4]
    .clock(x425_x8_1_clock),
    .reset(x425_x8_1_reset),
    .io_a(x425_x8_1_io_a),
    .io_b(x425_x8_1_io_b),
    .io_flow(x425_x8_1_io_flow),
    .io_result(x425_x8_1_io_result)
  );
  x406_x7 x426_x7_1 ( // @[Math.scala 150:24:@33835.4]
    .clock(x426_x7_1_clock),
    .reset(x426_x7_1_reset),
    .io_a(x426_x7_1_io_a),
    .io_b(x426_x7_1_io_b),
    .io_flow(x426_x7_1_io_flow),
    .io_result(x426_x7_1_io_result)
  );
  x406_x7 x427_x8_1 ( // @[Math.scala 150:24:@33845.4]
    .clock(x427_x8_1_clock),
    .reset(x427_x8_1_reset),
    .io_a(x427_x8_1_io_a),
    .io_b(x427_x8_1_io_b),
    .io_flow(x427_x8_1_io_flow),
    .io_result(x427_x8_1_io_result)
  );
  x406_x7 x428_x7_1 ( // @[Math.scala 150:24:@33855.4]
    .clock(x428_x7_1_clock),
    .reset(x428_x7_1_reset),
    .io_a(x428_x7_1_io_a),
    .io_b(x428_x7_1_io_b),
    .io_flow(x428_x7_1_io_flow),
    .io_result(x428_x7_1_io_result)
  );
  RetimeWrapper_321 RetimeWrapper_77 ( // @[package.scala 93:22:@33865.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x406_x7 x429_sum_1 ( // @[Math.scala 150:24:@33874.4]
    .clock(x429_sum_1_clock),
    .reset(x429_sum_1_reset),
    .io_a(x429_sum_1_io_a),
    .io_b(x429_sum_1_io_b),
    .io_flow(x429_sum_1_io_flow),
    .io_result(x429_sum_1_io_result)
  );
  x414 x430_1 ( // @[Math.scala 720:24:@33884.4]
    .io_b(x430_1_io_b),
    .io_result(x430_1_io_result)
  );
  x415_mul x431_mul_1 ( // @[Math.scala 262:24:@33895.4]
    .clock(x431_mul_1_clock),
    .io_a(x431_mul_1_io_a),
    .io_b(x431_mul_1_io_b),
    .io_flow(x431_mul_1_io_flow),
    .io_result(x431_mul_1_io_result)
  );
  x416 x432_1 ( // @[Math.scala 720:24:@33905.4]
    .io_b(x432_1_io_b),
    .io_result(x432_1_io_result)
  );
  RetimeWrapper_340 RetimeWrapper_78 ( // @[package.scala 93:22:@33914.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_341 RetimeWrapper_79 ( // @[package.scala 93:22:@33923.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_340 RetimeWrapper_80 ( // @[package.scala 93:22:@33932.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_343 RetimeWrapper_81 ( // @[package.scala 93:22:@33941.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_343 RetimeWrapper_82 ( // @[package.scala 93:22:@33950.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_83 ( // @[package.scala 93:22:@33959.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_340 RetimeWrapper_84 ( // @[package.scala 93:22:@33970.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_85 ( // @[package.scala 93:22:@33991.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_348 RetimeWrapper_86 ( // @[package.scala 93:22:@34000.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_341 RetimeWrapper_87 ( // @[package.scala 93:22:@34009.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_340 RetimeWrapper_88 ( // @[package.scala 93:22:@34020.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_343 RetimeWrapper_89 ( // @[package.scala 93:22:@34041.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_90 ( // @[package.scala 93:22:@34050.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_348 RetimeWrapper_91 ( // @[package.scala 93:22:@34059.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_92 ( // @[package.scala 93:22:@34068.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_93 ( // @[package.scala 93:22:@34077.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_356 RetimeWrapper_94 ( // @[package.scala 93:22:@34086.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_95 ( // @[package.scala 93:22:@34098.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_358 RetimeWrapper_96 ( // @[package.scala 93:22:@34119.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_348 RetimeWrapper_97 ( // @[package.scala 93:22:@34128.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_356 RetimeWrapper_98 ( // @[package.scala 93:22:@34137.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_99 ( // @[package.scala 93:22:@34149.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_100 ( // @[package.scala 93:22:@34170.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_363 RetimeWrapper_101 ( // @[package.scala 93:22:@34179.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_364 RetimeWrapper_102 ( // @[package.scala 93:22:@34188.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_103 ( // @[package.scala 93:22:@34200.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_363 RetimeWrapper_104 ( // @[package.scala 93:22:@34221.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_105 ( // @[package.scala 93:22:@34230.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_106 ( // @[package.scala 93:22:@34239.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_107 ( // @[package.scala 93:22:@34251.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_108 ( // @[package.scala 93:22:@34272.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_109 ( // @[package.scala 93:22:@34281.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_110 ( // @[package.scala 93:22:@34293.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_355 RetimeWrapper_111 ( // @[package.scala 93:22:@34314.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_112 ( // @[package.scala 93:22:@34323.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_352 RetimeWrapper_113 ( // @[package.scala 93:22:@34335.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  x406_x7 x451_x9_1 ( // @[Math.scala 150:24:@34368.4]
    .clock(x451_x9_1_clock),
    .reset(x451_x9_1_reset),
    .io_a(x451_x9_1_io_a),
    .io_b(x451_x9_1_io_b),
    .io_flow(x451_x9_1_io_flow),
    .io_result(x451_x9_1_io_result)
  );
  x406_x7 x452_x10_1 ( // @[Math.scala 150:24:@34378.4]
    .clock(x452_x10_1_clock),
    .reset(x452_x10_1_reset),
    .io_a(x452_x10_1_io_a),
    .io_b(x452_x10_1_io_b),
    .io_flow(x452_x10_1_io_flow),
    .io_result(x452_x10_1_io_result)
  );
  x406_x7 x453_sum_1 ( // @[Math.scala 150:24:@34388.4]
    .clock(x453_sum_1_clock),
    .reset(x453_sum_1_reset),
    .io_a(x453_sum_1_io_a),
    .io_b(x453_sum_1_io_b),
    .io_flow(x453_sum_1_io_flow),
    .io_result(x453_sum_1_io_result)
  );
  x414 x454_1 ( // @[Math.scala 720:24:@34398.4]
    .io_b(x454_1_io_b),
    .io_result(x454_1_io_result)
  );
  x415_mul x455_mul_1 ( // @[Math.scala 262:24:@34409.4]
    .clock(x455_mul_1_clock),
    .io_a(x455_mul_1_io_a),
    .io_b(x455_mul_1_io_b),
    .io_flow(x455_mul_1_io_flow),
    .io_result(x455_mul_1_io_result)
  );
  x416 x456_1 ( // @[Math.scala 720:24:@34421.4]
    .io_b(x456_1_io_b),
    .io_result(x456_1_io_result)
  );
  x406_x7 x459_x9_1 ( // @[Math.scala 150:24:@34440.4]
    .clock(x459_x9_1_clock),
    .reset(x459_x9_1_reset),
    .io_a(x459_x9_1_io_a),
    .io_b(x459_x9_1_io_b),
    .io_flow(x459_x9_1_io_flow),
    .io_result(x459_x9_1_io_result)
  );
  x406_x7 x460_x10_1 ( // @[Math.scala 150:24:@34450.4]
    .clock(x460_x10_1_clock),
    .reset(x460_x10_1_reset),
    .io_a(x460_x10_1_io_a),
    .io_b(x460_x10_1_io_b),
    .io_flow(x460_x10_1_io_flow),
    .io_result(x460_x10_1_io_result)
  );
  x406_x7 x461_sum_1 ( // @[Math.scala 150:24:@34460.4]
    .clock(x461_sum_1_clock),
    .reset(x461_sum_1_reset),
    .io_a(x461_sum_1_io_a),
    .io_b(x461_sum_1_io_b),
    .io_flow(x461_sum_1_io_flow),
    .io_result(x461_sum_1_io_result)
  );
  x414 x462_1 ( // @[Math.scala 720:24:@34470.4]
    .io_b(x462_1_io_b),
    .io_result(x462_1_io_result)
  );
  x415_mul x463_mul_1 ( // @[Math.scala 262:24:@34481.4]
    .clock(x463_mul_1_clock),
    .io_a(x463_mul_1_io_a),
    .io_b(x463_mul_1_io_b),
    .io_flow(x463_mul_1_io_flow),
    .io_result(x463_mul_1_io_result)
  );
  x416 x464_1 ( // @[Math.scala 720:24:@34491.4]
    .io_b(x464_1_io_b),
    .io_result(x464_1_io_result)
  );
  RetimeWrapper_382 RetimeWrapper_114 ( // @[package.scala 93:22:@34506.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_383 RetimeWrapper_115 ( // @[package.scala 93:22:@34515.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_383 RetimeWrapper_116 ( // @[package.scala 93:22:@34524.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_383 RetimeWrapper_117 ( // @[package.scala 93:22:@34533.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  assign b297 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 62:18:@31980.4]
  assign b298 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 63:18:@31981.4]
  assign _T_205 = b297 & b298; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 67:30:@31983.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 67:37:@31984.4]
  assign _T_210 = io_in_x266_TID == 8'h0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:76:@31989.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:62:@31990.4]
  assign _T_213 = io_in_x266_TDEST == 8'h0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:101:@31991.4]
  assign x547_x299_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@32000.4 package.scala 96:25:@32001.4]
  assign b295_number = __io_result; // @[Math.scala 723:22:@31965.4 Math.scala 724:14:@31966.4]
  assign _T_244 = $signed(b295_number); // @[Math.scala 406:49:@32166.4]
  assign _T_246 = $signed(_T_244) & $signed(32'sh3); // @[Math.scala 406:56:@32168.4]
  assign _T_247 = $signed(_T_246); // @[Math.scala 406:56:@32169.4]
  assign x523_number = $unsigned(_T_247); // @[implicits.scala 133:21:@32170.4]
  assign _T_257 = $signed(x523_number); // @[Math.scala 406:49:@32179.4]
  assign _T_259 = $signed(_T_257) & $signed(32'sh3); // @[Math.scala 406:56:@32181.4]
  assign _T_260 = $signed(_T_259); // @[Math.scala 406:56:@32182.4]
  assign b296_number = __1_io_result; // @[Math.scala 723:22:@31977.4 Math.scala 724:14:@31978.4]
  assign _T_269 = $signed(b296_number); // @[Math.scala 406:49:@32190.4]
  assign _T_271 = $signed(_T_269) & $signed(32'sh3); // @[Math.scala 406:56:@32192.4]
  assign _T_272 = $signed(_T_271); // @[Math.scala 406:56:@32193.4]
  assign _T_276 = x523_number[31]; // @[FixedPoint.scala 50:25:@32199.4]
  assign _T_280 = _T_276 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32201.4]
  assign _T_281 = x523_number[31:2]; // @[FixedPoint.scala 18:52:@32202.4]
  assign _T_287 = _T_281 == 30'h3fffffff; // @[Math.scala 451:55:@32204.4]
  assign _T_288 = x523_number[1:0]; // @[FixedPoint.scala 18:52:@32205.4]
  assign _T_294 = _T_288 != 2'h0; // @[Math.scala 451:110:@32207.4]
  assign _T_295 = _T_287 & _T_294; // @[Math.scala 451:94:@32208.4]
  assign _T_297 = {_T_280,_T_281}; // @[Cat.scala 30:58:@32210.4]
  assign x308_1_number = _T_295 ? 32'h0 : _T_297; // @[Math.scala 454:20:@32211.4]
  assign _GEN_0 = {{9'd0}, x308_1_number}; // @[Math.scala 461:32:@32216.4]
  assign _T_302 = _GEN_0 << 9; // @[Math.scala 461:32:@32216.4]
  assign _GEN_1 = {{5'd0}, x308_1_number}; // @[Math.scala 461:32:@32221.4]
  assign _T_305 = _GEN_1 << 5; // @[Math.scala 461:32:@32221.4]
  assign _T_311 = b296_number[31]; // @[FixedPoint.scala 50:25:@32236.4]
  assign _T_315 = _T_311 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32238.4]
  assign _T_316 = b296_number[31:2]; // @[FixedPoint.scala 18:52:@32239.4]
  assign _T_322 = _T_316 == 30'h3fffffff; // @[Math.scala 451:55:@32241.4]
  assign _T_323 = b296_number[1:0]; // @[FixedPoint.scala 18:52:@32242.4]
  assign _T_329 = _T_323 != 2'h0; // @[Math.scala 451:110:@32244.4]
  assign _T_330 = _T_322 & _T_329; // @[Math.scala 451:94:@32245.4]
  assign _T_332 = {_T_315,_T_316}; // @[Cat.scala 30:58:@32247.4]
  assign _T_360 = ~ io_sigsIn_break; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:101:@32324.4]
  assign _T_364 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@32332.4 package.scala 96:25:@32333.4]
  assign _T_366 = io_rr ? _T_364 : 1'h0; // @[implicits.scala 55:10:@32334.4]
  assign _T_367 = _T_360 & _T_366; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:118:@32335.4]
  assign _T_369 = _T_367 & _T_360; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:206:@32337.4]
  assign _T_370 = _T_369 & io_sigsIn_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:225:@32338.4]
  assign x549_b297_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@32276.4 package.scala 96:25:@32277.4]
  assign _T_371 = _T_370 & x549_b297_D3; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 118:251:@32339.4]
  assign x551_b298_D3 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@32294.4 package.scala 96:25:@32295.4]
  assign x313_rdcol_number = x313_rdcol_1_io_result; // @[Math.scala 154:22:@32356.4 Math.scala 155:14:@32357.4]
  assign _T_388 = $signed(x313_rdcol_number); // @[Math.scala 406:49:@32365.4]
  assign _T_390 = $signed(_T_388) & $signed(32'sh3); // @[Math.scala 406:56:@32367.4]
  assign _T_391 = $signed(_T_390); // @[Math.scala 406:56:@32368.4]
  assign _T_395 = x313_rdcol_number[31]; // @[FixedPoint.scala 50:25:@32374.4]
  assign _T_399 = _T_395 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32376.4]
  assign _T_400 = x313_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@32377.4]
  assign _T_406 = _T_400 == 30'h3fffffff; // @[Math.scala 451:55:@32379.4]
  assign _T_407 = x313_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@32380.4]
  assign _T_413 = _T_407 != 2'h0; // @[Math.scala 451:110:@32382.4]
  assign _T_414 = _T_406 & _T_413; // @[Math.scala 451:94:@32383.4]
  assign _T_416 = {_T_399,_T_400}; // @[Cat.scala 30:58:@32385.4]
  assign _T_436 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@32434.4 package.scala 96:25:@32435.4]
  assign _T_438 = io_rr ? _T_436 : 1'h0; // @[implicits.scala 55:10:@32436.4]
  assign _T_439 = _T_360 & _T_438; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:118:@32437.4]
  assign _T_441 = _T_439 & _T_360; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:206:@32439.4]
  assign _T_442 = _T_441 & io_sigsIn_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:225:@32440.4]
  assign _T_443 = _T_442 & x549_b297_D3; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 139:251:@32441.4]
  assign x558_b295_D6_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@32455.4 package.scala 96:25:@32456.4]
  assign _T_453 = $signed(x558_b295_D6_number); // @[Math.scala 476:37:@32461.4]
  assign x320 = $signed(_T_453) < $signed(32'sh0); // @[Math.scala 476:44:@32463.4]
  assign x559_x313_rdcol_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@32471.4 package.scala 96:25:@32472.4]
  assign _T_464 = $signed(x559_x313_rdcol_D6_number); // @[Math.scala 476:37:@32477.4]
  assign x321 = $signed(_T_464) < $signed(32'sh0); // @[Math.scala 476:44:@32479.4]
  assign x560_x320_D1 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@32487.4 package.scala 96:25:@32488.4]
  assign x322 = x560_x320_D1 | x321; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 152:24:@32491.4]
  assign _T_503 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@32559.4 package.scala 96:25:@32560.4]
  assign _T_505 = io_rr ? _T_503 : 1'h0; // @[implicits.scala 55:10:@32561.4]
  assign _T_506 = _T_360 & _T_505; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 171:146:@32562.4]
  assign x565_x323_D2 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@32538.4 package.scala 96:25:@32539.4]
  assign _T_507 = _T_506 & x565_x323_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 171:234:@32563.4]
  assign x562_b297_D9 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@32511.4 package.scala 96:25:@32512.4]
  assign _T_508 = _T_507 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 171:242:@32564.4]
  assign x564_b298_D9 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@32529.4 package.scala 96:25:@32530.4]
  assign x567_b296_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@32580.4 package.scala 96:25:@32581.4]
  assign _T_521 = $signed(x567_b296_D6_number); // @[Math.scala 476:37:@32588.4]
  assign x326 = $signed(_T_521) < $signed(32'sh0); // @[Math.scala 476:44:@32590.4]
  assign x327 = x320 | x326; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 187:59:@32593.4]
  assign _T_548 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@32634.4 package.scala 96:25:@32635.4]
  assign _T_550 = io_rr ? _T_548 : 1'h0; // @[implicits.scala 55:10:@32636.4]
  assign _T_551 = _T_360 & _T_550; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:194:@32637.4]
  assign x568_x328_D3 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@32604.4 package.scala 96:25:@32605.4]
  assign _T_552 = _T_551 & x568_x328_D3; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:282:@32638.4]
  assign _T_553 = _T_552 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:290:@32639.4]
  assign x331_rdcol_number = x331_rdcol_1_io_result; // @[Math.scala 154:22:@32658.4 Math.scala 155:14:@32659.4]
  assign _T_568 = $signed(x331_rdcol_number); // @[Math.scala 476:37:@32664.4]
  assign x332 = $signed(_T_568) < $signed(32'sh0); // @[Math.scala 476:44:@32666.4]
  assign x333 = x560_x320_D1 | x332; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 208:59:@32669.4]
  assign _T_584 = $signed(_T_568) & $signed(32'sh3); // @[Math.scala 406:56:@32680.4]
  assign _T_585 = $signed(_T_584); // @[Math.scala 406:56:@32681.4]
  assign _T_589 = x331_rdcol_number[31]; // @[FixedPoint.scala 50:25:@32687.4]
  assign _T_593 = _T_589 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32689.4]
  assign _T_594 = x331_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@32690.4]
  assign _T_600 = _T_594 == 30'h3fffffff; // @[Math.scala 451:55:@32692.4]
  assign _T_601 = x331_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@32693.4]
  assign _T_607 = _T_601 != 2'h0; // @[Math.scala 451:110:@32695.4]
  assign _T_608 = _T_600 & _T_607; // @[Math.scala 451:94:@32696.4]
  assign _T_610 = {_T_593,_T_594}; // @[Cat.scala 30:58:@32698.4]
  assign _T_639 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@32757.4 package.scala 96:25:@32758.4]
  assign _T_641 = io_rr ? _T_639 : 1'h0; // @[implicits.scala 55:10:@32759.4]
  assign _T_642 = _T_360 & _T_641; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:194:@32760.4]
  assign x572_x334_D2 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@32727.4 package.scala 96:25:@32728.4]
  assign _T_643 = _T_642 & x572_x334_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:282:@32761.4]
  assign _T_644 = _T_643 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:290:@32762.4]
  assign x340_rdcol_number = x340_rdcol_1_io_result; // @[Math.scala 154:22:@32781.4 Math.scala 155:14:@32782.4]
  assign _T_659 = $signed(x340_rdcol_number); // @[Math.scala 476:37:@32787.4]
  assign x341 = $signed(_T_659) < $signed(32'sh0); // @[Math.scala 476:44:@32789.4]
  assign x342 = x560_x320_D1 | x341; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 237:59:@32792.4]
  assign _T_675 = $signed(_T_659) & $signed(32'sh3); // @[Math.scala 406:56:@32803.4]
  assign _T_676 = $signed(_T_675); // @[Math.scala 406:56:@32804.4]
  assign _T_680 = x340_rdcol_number[31]; // @[FixedPoint.scala 50:25:@32810.4]
  assign _T_684 = _T_680 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32812.4]
  assign _T_685 = x340_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@32813.4]
  assign _T_691 = _T_685 == 30'h3fffffff; // @[Math.scala 451:55:@32815.4]
  assign _T_692 = x340_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@32816.4]
  assign _T_698 = _T_692 != 2'h0; // @[Math.scala 451:110:@32818.4]
  assign _T_699 = _T_691 & _T_698; // @[Math.scala 451:94:@32819.4]
  assign _T_701 = {_T_684,_T_685}; // @[Cat.scala 30:58:@32821.4]
  assign _T_727 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@32871.4 package.scala 96:25:@32872.4]
  assign _T_729 = io_rr ? _T_727 : 1'h0; // @[implicits.scala 55:10:@32873.4]
  assign _T_730 = _T_360 & _T_729; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 256:194:@32874.4]
  assign x575_x343_D2 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@32841.4 package.scala 96:25:@32842.4]
  assign _T_731 = _T_730 & x575_x343_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 256:282:@32875.4]
  assign _T_732 = _T_731 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 256:290:@32876.4]
  assign x349_rdrow_number = x349_rdrow_1_io_result; // @[Math.scala 195:22:@32895.4 Math.scala 196:14:@32896.4]
  assign _T_749 = $signed(x349_rdrow_number); // @[Math.scala 406:49:@32902.4]
  assign _T_751 = $signed(_T_749) & $signed(32'sh3); // @[Math.scala 406:56:@32904.4]
  assign _T_752 = $signed(_T_751); // @[Math.scala 406:56:@32905.4]
  assign x532_number = $unsigned(_T_752); // @[implicits.scala 133:21:@32906.4]
  assign x351 = $signed(_T_749) < $signed(32'sh0); // @[Math.scala 476:44:@32914.4]
  assign x352 = x351 | x321; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 266:24:@32917.4]
  assign _T_773 = $signed(x532_number); // @[Math.scala 406:49:@32926.4]
  assign _T_775 = $signed(_T_773) & $signed(32'sh3); // @[Math.scala 406:56:@32928.4]
  assign _T_776 = $signed(_T_775); // @[Math.scala 406:56:@32929.4]
  assign _T_780 = x532_number[31]; // @[FixedPoint.scala 50:25:@32935.4]
  assign _T_784 = _T_780 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32937.4]
  assign _T_785 = x532_number[31:2]; // @[FixedPoint.scala 18:52:@32938.4]
  assign _T_791 = _T_785 == 30'h3fffffff; // @[Math.scala 451:55:@32940.4]
  assign _T_792 = x532_number[1:0]; // @[FixedPoint.scala 18:52:@32941.4]
  assign _T_798 = _T_792 != 2'h0; // @[Math.scala 451:110:@32943.4]
  assign _T_799 = _T_791 & _T_798; // @[Math.scala 451:94:@32944.4]
  assign _T_801 = {_T_784,_T_785}; // @[Cat.scala 30:58:@32946.4]
  assign x355_1_number = _T_799 ? 32'h0 : _T_801; // @[Math.scala 454:20:@32947.4]
  assign _GEN_2 = {{9'd0}, x355_1_number}; // @[Math.scala 461:32:@32952.4]
  assign _T_806 = _GEN_2 << 9; // @[Math.scala 461:32:@32952.4]
  assign _GEN_3 = {{5'd0}, x355_1_number}; // @[Math.scala 461:32:@32957.4]
  assign _T_809 = _GEN_3 << 5; // @[Math.scala 461:32:@32957.4]
  assign _T_836 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@33016.4 package.scala 96:25:@33017.4]
  assign _T_838 = io_rr ? _T_836 : 1'h0; // @[implicits.scala 55:10:@33018.4]
  assign _T_839 = _T_360 & _T_838; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:194:@33019.4]
  assign x580_x353_D2 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@33004.4 package.scala 96:25:@33005.4]
  assign _T_840 = _T_839 & x580_x353_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:282:@33020.4]
  assign _T_841 = _T_840 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:290:@33021.4]
  assign x581_x326_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@33037.4 package.scala 96:25:@33038.4]
  assign x360 = x351 | x581_x326_D1; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 303:59:@33041.4]
  assign _T_873 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@33085.4 package.scala 96:25:@33086.4]
  assign _T_875 = io_rr ? _T_873 : 1'h0; // @[implicits.scala 55:10:@33087.4]
  assign _T_876 = _T_360 & _T_875; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:194:@33088.4]
  assign x583_x361_D2 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@33073.4 package.scala 96:25:@33074.4]
  assign _T_877 = _T_876 & x583_x361_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:282:@33089.4]
  assign _T_878 = _T_877 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:290:@33090.4]
  assign x365 = x351 | x332; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 322:59:@33101.4]
  assign _T_905 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@33143.4 package.scala 96:25:@33144.4]
  assign _T_907 = io_rr ? _T_905 : 1'h0; // @[implicits.scala 55:10:@33145.4]
  assign _T_908 = _T_360 & _T_907; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:194:@33146.4]
  assign x585_x366_D2 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@33131.4 package.scala 96:25:@33132.4]
  assign _T_909 = _T_908 & x585_x366_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:282:@33147.4]
  assign _T_910 = _T_909 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:290:@33148.4]
  assign x370 = x351 | x341; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 339:59:@33159.4]
  assign _T_937 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@33201.4 package.scala 96:25:@33202.4]
  assign _T_939 = io_rr ? _T_937 : 1'h0; // @[implicits.scala 55:10:@33203.4]
  assign _T_940 = _T_360 & _T_939; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:194:@33204.4]
  assign x587_x371_D2 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@33189.4 package.scala 96:25:@33190.4]
  assign _T_941 = _T_940 & x587_x371_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:282:@33205.4]
  assign _T_942 = _T_941 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:290:@33206.4]
  assign x375_rdrow_number = x375_rdrow_1_io_result; // @[Math.scala 195:22:@33225.4 Math.scala 196:14:@33226.4]
  assign _T_959 = $signed(x375_rdrow_number); // @[Math.scala 406:49:@33232.4]
  assign _T_961 = $signed(_T_959) & $signed(32'sh3); // @[Math.scala 406:56:@33234.4]
  assign _T_962 = $signed(_T_961); // @[Math.scala 406:56:@33235.4]
  assign x537_number = $unsigned(_T_962); // @[implicits.scala 133:21:@33236.4]
  assign x377 = $signed(_T_959) < $signed(32'sh0); // @[Math.scala 476:44:@33244.4]
  assign x378 = x377 | x321; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 362:24:@33247.4]
  assign _T_983 = $signed(x537_number); // @[Math.scala 406:49:@33256.4]
  assign _T_985 = $signed(_T_983) & $signed(32'sh3); // @[Math.scala 406:56:@33258.4]
  assign _T_986 = $signed(_T_985); // @[Math.scala 406:56:@33259.4]
  assign _T_990 = x537_number[31]; // @[FixedPoint.scala 50:25:@33265.4]
  assign _T_994 = _T_990 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33267.4]
  assign _T_995 = x537_number[31:2]; // @[FixedPoint.scala 18:52:@33268.4]
  assign _T_1001 = _T_995 == 30'h3fffffff; // @[Math.scala 451:55:@33270.4]
  assign _T_1002 = x537_number[1:0]; // @[FixedPoint.scala 18:52:@33271.4]
  assign _T_1008 = _T_1002 != 2'h0; // @[Math.scala 451:110:@33273.4]
  assign _T_1009 = _T_1001 & _T_1008; // @[Math.scala 451:94:@33274.4]
  assign _T_1011 = {_T_994,_T_995}; // @[Cat.scala 30:58:@33276.4]
  assign x381_1_number = _T_1009 ? 32'h0 : _T_1011; // @[Math.scala 454:20:@33277.4]
  assign _GEN_4 = {{9'd0}, x381_1_number}; // @[Math.scala 461:32:@33282.4]
  assign _T_1016 = _GEN_4 << 9; // @[Math.scala 461:32:@33282.4]
  assign _GEN_5 = {{5'd0}, x381_1_number}; // @[Math.scala 461:32:@33287.4]
  assign _T_1019 = _GEN_5 << 5; // @[Math.scala 461:32:@33287.4]
  assign _T_1043 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@33337.4 package.scala 96:25:@33338.4]
  assign _T_1045 = io_rr ? _T_1043 : 1'h0; // @[implicits.scala 55:10:@33339.4]
  assign _T_1046 = _T_360 & _T_1045; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 385:194:@33340.4]
  assign x588_x379_D2 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@33316.4 package.scala 96:25:@33317.4]
  assign _T_1047 = _T_1046 & x588_x379_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 385:282:@33341.4]
  assign _T_1048 = _T_1047 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 385:290:@33342.4]
  assign x386 = x377 | x581_x326_D1; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 389:24:@33353.4]
  assign _T_1072 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@33386.4 package.scala 96:25:@33387.4]
  assign _T_1074 = io_rr ? _T_1072 : 1'h0; // @[implicits.scala 55:10:@33388.4]
  assign _T_1075 = _T_360 & _T_1074; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:194:@33389.4]
  assign x590_x387_D2 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@33374.4 package.scala 96:25:@33375.4]
  assign _T_1076 = _T_1075 & x590_x387_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:282:@33390.4]
  assign _T_1077 = _T_1076 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:290:@33391.4]
  assign x391 = x377 | x332; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 404:24:@33402.4]
  assign _T_1101 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@33435.4 package.scala 96:25:@33436.4]
  assign _T_1103 = io_rr ? _T_1101 : 1'h0; // @[implicits.scala 55:10:@33437.4]
  assign _T_1104 = _T_360 & _T_1103; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:194:@33438.4]
  assign x591_x392_D2 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@33423.4 package.scala 96:25:@33424.4]
  assign _T_1105 = _T_1104 & x591_x392_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:282:@33439.4]
  assign _T_1106 = _T_1105 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:290:@33440.4]
  assign x396 = x377 | x341; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 425:59:@33451.4]
  assign _T_1132 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@33486.4 package.scala 96:25:@33487.4]
  assign _T_1134 = io_rr ? _T_1132 : 1'h0; // @[implicits.scala 55:10:@33488.4]
  assign _T_1135 = _T_360 & _T_1134; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 438:194:@33489.4]
  assign x592_x397_D2 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@33474.4 package.scala 96:25:@33475.4]
  assign _T_1136 = _T_1135 & x592_x397_D2; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 438:282:@33490.4]
  assign _T_1137 = _T_1136 & x562_b297_D9; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 438:290:@33491.4]
  assign x329_rd_0_number = x301_lb_0_io_rPort_3_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 196:29:@32625.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 200:407:@32646.4]
  assign _GEN_6 = {{1'd0}, x329_rd_0_number}; // @[Math.scala 461:32:@33503.4]
  assign x358_rd_0_number = x301_lb_0_io_rPort_11_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 287:29:@33007.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 291:407:@33028.4]
  assign _GEN_7 = {{1'd0}, x358_rd_0_number}; // @[Math.scala 461:32:@33515.4]
  assign x363_rd_0_number = x301_lb_0_io_rPort_8_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 314:29:@33076.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 318:407:@33097.4]
  assign _GEN_8 = {{2'd0}, x363_rd_0_number}; // @[Math.scala 461:32:@33527.4]
  assign x368_rd_0_number = x301_lb_0_io_rPort_9_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 331:29:@33134.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 335:407:@33155.4]
  assign _GEN_9 = {{1'd0}, x368_rd_0_number}; // @[Math.scala 461:32:@33539.4]
  assign x389_rd_0_number = x301_lb_0_io_rPort_2_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 396:29:@33377.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 400:407:@33398.4]
  assign _GEN_10 = {{1'd0}, x389_rd_0_number}; // @[Math.scala 461:32:@33551.4]
  assign x338_rd_0_number = x301_lb_0_io_rPort_7_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 225:29:@32748.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 229:407:@32769.4]
  assign _GEN_11 = {{1'd0}, x338_rd_0_number}; // @[Math.scala 461:32:@33709.4]
  assign _GEN_12 = {{1'd0}, x363_rd_0_number}; // @[Math.scala 461:32:@33721.4]
  assign _GEN_13 = {{2'd0}, x368_rd_0_number}; // @[Math.scala 461:32:@33733.4]
  assign x373_rd_0_number = x301_lb_0_io_rPort_10_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 348:29:@33192.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 352:407:@33213.4]
  assign _GEN_14 = {{1'd0}, x373_rd_0_number}; // @[Math.scala 461:32:@33745.4]
  assign x394_rd_0_number = x301_lb_0_io_rPort_6_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 411:29:@33426.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 415:407:@33447.4]
  assign _GEN_15 = {{1'd0}, x394_rd_0_number}; // @[Math.scala 461:32:@33757.4]
  assign _T_1311 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@33975.4 package.scala 96:25:@33976.4]
  assign _T_1313 = io_rr ? _T_1311 : 1'h0; // @[implicits.scala 55:10:@33977.4]
  assign _T_1314 = _T_360 & _T_1313; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:167:@33978.4]
  assign _T_1316 = _T_1314 & _T_360; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:256:@33980.4]
  assign _T_1317 = _T_1316 & io_sigsIn_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:275:@33981.4]
  assign x601_b297_D23 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@33919.4 package.scala 96:25:@33920.4]
  assign _T_1318 = _T_1317 & x601_b297_D23; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 544:301:@33982.4]
  assign x603_b298_D23 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@33937.4 package.scala 96:25:@33938.4]
  assign _T_1334 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@34025.4 package.scala 96:25:@34026.4]
  assign _T_1336 = io_rr ? _T_1334 : 1'h0; // @[implicits.scala 55:10:@34027.4]
  assign _T_1337 = _T_360 & _T_1336; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:167:@34028.4]
  assign _T_1339 = _T_1337 & _T_360; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:256:@34030.4]
  assign _T_1340 = _T_1339 & io_sigsIn_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:275:@34031.4]
  assign _T_1341 = _T_1340 & x601_b297_D23; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 555:301:@34032.4]
  assign _T_1372 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@34103.4 package.scala 96:25:@34104.4]
  assign _T_1374 = io_rr ? _T_1372 : 1'h0; // @[implicits.scala 55:10:@34105.4]
  assign _T_1375 = _T_360 & _T_1374; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 573:195:@34106.4]
  assign x614_x323_D17 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@34082.4 package.scala 96:25:@34083.4]
  assign _T_1376 = _T_1375 & x614_x323_D17; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 573:284:@34107.4]
  assign x611_b297_D24 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@34055.4 package.scala 96:25:@34056.4]
  assign _T_1377 = _T_1376 & x611_b297_D24; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 573:292:@34108.4]
  assign x613_b298_D24 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@34073.4 package.scala 96:25:@34074.4]
  assign _T_1400 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@34154.4 package.scala 96:25:@34155.4]
  assign _T_1402 = io_rr ? _T_1400 : 1'h0; // @[implicits.scala 55:10:@34156.4]
  assign _T_1403 = _T_360 & _T_1402; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:195:@34157.4]
  assign x616_x328_D18 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@34124.4 package.scala 96:25:@34125.4]
  assign _T_1404 = _T_1403 & x616_x328_D18; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:284:@34158.4]
  assign _T_1405 = _T_1404 & x611_b297_D24; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:292:@34159.4]
  assign _T_1428 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@34205.4 package.scala 96:25:@34206.4]
  assign _T_1430 = io_rr ? _T_1428 : 1'h0; // @[implicits.scala 55:10:@34207.4]
  assign _T_1431 = _T_360 & _T_1430; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:195:@34208.4]
  assign x619_x334_D17 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@34175.4 package.scala 96:25:@34176.4]
  assign _T_1432 = _T_1431 & x619_x334_D17; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:284:@34209.4]
  assign _T_1433 = _T_1432 & x611_b297_D24; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:292:@34210.4]
  assign _T_1456 = RetimeWrapper_107_io_out; // @[package.scala 96:25:@34256.4 package.scala 96:25:@34257.4]
  assign _T_1458 = io_rr ? _T_1456 : 1'h0; // @[implicits.scala 55:10:@34258.4]
  assign _T_1459 = _T_360 & _T_1458; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:195:@34259.4]
  assign x624_x353_D17 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@34244.4 package.scala 96:25:@34245.4]
  assign _T_1460 = _T_1459 & x624_x353_D17; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:284:@34260.4]
  assign _T_1461 = _T_1460 & x611_b297_D24; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:292:@34261.4]
  assign _T_1481 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@34298.4 package.scala 96:25:@34299.4]
  assign _T_1483 = io_rr ? _T_1481 : 1'h0; // @[implicits.scala 55:10:@34300.4]
  assign _T_1484 = _T_360 & _T_1483; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:195:@34301.4]
  assign x625_x361_D17 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@34277.4 package.scala 96:25:@34278.4]
  assign _T_1485 = _T_1484 & x625_x361_D17; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:284:@34302.4]
  assign _T_1486 = _T_1485 & x611_b297_D24; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:292:@34303.4]
  assign _T_1506 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@34340.4 package.scala 96:25:@34341.4]
  assign _T_1508 = io_rr ? _T_1506 : 1'h0; // @[implicits.scala 55:10:@34342.4]
  assign _T_1509 = _T_360 & _T_1508; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 634:195:@34343.4]
  assign x627_x366_D17 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@34319.4 package.scala 96:25:@34320.4]
  assign _T_1510 = _T_1509 & x627_x366_D17; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 634:284:@34344.4]
  assign _T_1511 = _T_1510 & x611_b297_D24; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 634:292:@34345.4]
  assign x439_rd_0_number = x302_lb2_0_io_rPort_1_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 582:29:@34145.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 586:339:@34166.4]
  assign _GEN_16 = {{1'd0}, x439_rd_0_number}; // @[Math.scala 461:32:@34359.4]
  assign _T_1518 = _GEN_16 << 1; // @[Math.scala 461:32:@34359.4]
  assign x443_rd_0_number = x302_lb2_0_io_rPort_0_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 608:29:@34247.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 612:339:@34268.4]
  assign _GEN_17 = {{2'd0}, x443_rd_0_number}; // @[Math.scala 461:32:@34364.4]
  assign _T_1521 = _GEN_17 << 2; // @[Math.scala 461:32:@34364.4]
  assign x441_rd_0_number = x302_lb2_0_io_rPort_3_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 595:29:@34196.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 599:339:@34217.4]
  assign _GEN_18 = {{1'd0}, x441_rd_0_number}; // @[Math.scala 461:32:@34431.4]
  assign _T_1548 = _GEN_18 << 1; // @[Math.scala 461:32:@34431.4]
  assign x445_rd_0_number = x302_lb2_0_io_rPort_2_output_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 619:29:@34289.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 623:339:@34310.4]
  assign _GEN_19 = {{2'd0}, x445_rd_0_number}; // @[Math.scala 461:32:@34436.4]
  assign _T_1551 = _GEN_19 << 2; // @[Math.scala 461:32:@34436.4]
  assign x456_number = x456_1_io_result; // @[Math.scala 723:22:@34426.4 Math.scala 724:14:@34427.4]
  assign x464_number = x464_1_io_result; // @[Math.scala 723:22:@34496.4 Math.scala 724:14:@34497.4]
  assign _T_1595 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@34538.4 package.scala 96:25:@34539.4]
  assign _T_1597 = io_rr ? _T_1595 : 1'h0; // @[implicits.scala 55:10:@34540.4]
  assign x630_b297_D37 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@34529.4 package.scala 96:25:@34530.4]
  assign _T_1598 = _T_1597 & x630_b297_D37; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 688:117:@34541.4]
  assign x629_b298_D37 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@34520.4 package.scala 96:25:@34521.4]
  assign _T_1599 = _T_1598 & x629_b298_D37; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 688:123:@34542.4]
  assign x550_x311_sum_D1_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32285.4 package.scala 96:25:@32286.4]
  assign x552_x525_D3_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@32303.4 package.scala 96:25:@32304.4]
  assign x553_x524_D3_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@32312.4 package.scala 96:25:@32313.4]
  assign x555_x529_D2_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@32405.4 package.scala 96:25:@32406.4]
  assign x556_x317_sum_D1_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@32414.4 package.scala 96:25:@32415.4]
  assign x561_x529_D8_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@32502.4 package.scala 96:25:@32503.4]
  assign x563_x317_sum_D7_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@32520.4 package.scala 96:25:@32521.4]
  assign x566_x524_D9_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@32547.4 package.scala 96:25:@32548.4]
  assign x569_x311_sum_D7_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@32613.4 package.scala 96:25:@32614.4]
  assign x570_x525_D9_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@32622.4 package.scala 96:25:@32623.4]
  assign x573_x530_D2_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@32736.4 package.scala 96:25:@32737.4]
  assign x574_x337_sum_D1_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@32745.4 package.scala 96:25:@32746.4]
  assign x576_x531_D2_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@32850.4 package.scala 96:25:@32851.4]
  assign x577_x346_sum_D1_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@32859.4 package.scala 96:25:@32860.4]
  assign x357_sum_number = x357_sum_1_io_result; // @[Math.scala 154:22:@32986.4 Math.scala 155:14:@32987.4]
  assign x579_x533_D2_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@32995.4 package.scala 96:25:@32996.4]
  assign x362_sum_number = x362_sum_1_io_result; // @[Math.scala 154:22:@33064.4 Math.scala 155:14:@33065.4]
  assign x367_sum_number = x367_sum_1_io_result; // @[Math.scala 154:22:@33122.4 Math.scala 155:14:@33123.4]
  assign x372_sum_number = x372_sum_1_io_result; // @[Math.scala 154:22:@33180.4 Math.scala 155:14:@33181.4]
  assign x383_sum_number = x383_sum_1_io_result; // @[Math.scala 154:22:@33307.4 Math.scala 155:14:@33308.4]
  assign x589_x538_D2_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@33325.4 package.scala 96:25:@33326.4]
  assign x388_sum_number = x388_sum_1_io_result; // @[Math.scala 154:22:@33365.4 Math.scala 155:14:@33366.4]
  assign x393_sum_number = x393_sum_1_io_result; // @[Math.scala 154:22:@33414.4 Math.scala 155:14:@33415.4]
  assign x398_sum_number = x398_sum_1_io_result; // @[Math.scala 154:22:@33465.4 Math.scala 155:14:@33466.4]
  assign _T_1144 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@33509.4 package.scala 96:25:@33510.4]
  assign _T_1149 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@33521.4 package.scala 96:25:@33522.4]
  assign _T_1154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@33533.4 package.scala 96:25:@33534.4]
  assign _T_1159 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@33545.4 package.scala 96:25:@33546.4]
  assign _T_1164 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@33557.4 package.scala 96:25:@33558.4]
  assign _T_1218 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@33715.4 package.scala 96:25:@33716.4]
  assign _T_1223 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@33727.4 package.scala 96:25:@33728.4]
  assign _T_1228 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@33739.4 package.scala 96:25:@33740.4]
  assign _T_1233 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@33751.4 package.scala 96:25:@33752.4]
  assign _T_1238 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@33763.4 package.scala 96:25:@33764.4]
  assign x602_x311_sum_D21_number = RetimeWrapper_79_io_out; // @[package.scala 96:25:@33928.4 package.scala 96:25:@33929.4]
  assign x604_x525_D23_number = RetimeWrapper_81_io_out; // @[package.scala 96:25:@33946.4 package.scala 96:25:@33947.4]
  assign x605_x524_D23_number = RetimeWrapper_82_io_out; // @[package.scala 96:25:@33955.4 package.scala 96:25:@33956.4]
  assign x608_x529_D22_number = RetimeWrapper_86_io_out; // @[package.scala 96:25:@34005.4 package.scala 96:25:@34006.4]
  assign x609_x317_sum_D21_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@34014.4 package.scala 96:25:@34015.4]
  assign x610_x529_D23_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@34046.4 package.scala 96:25:@34047.4]
  assign x612_x317_sum_D22_number = RetimeWrapper_91_io_out; // @[package.scala 96:25:@34064.4 package.scala 96:25:@34065.4]
  assign x615_x524_D24_number = RetimeWrapper_94_io_out; // @[package.scala 96:25:@34091.4 package.scala 96:25:@34092.4]
  assign x617_x311_sum_D22_number = RetimeWrapper_97_io_out; // @[package.scala 96:25:@34133.4 package.scala 96:25:@34134.4]
  assign x618_x525_D24_number = RetimeWrapper_98_io_out; // @[package.scala 96:25:@34142.4 package.scala 96:25:@34143.4]
  assign x620_x530_D17_number = RetimeWrapper_101_io_out; // @[package.scala 96:25:@34184.4 package.scala 96:25:@34185.4]
  assign x621_x337_sum_D16_number = RetimeWrapper_102_io_out; // @[package.scala 96:25:@34193.4 package.scala 96:25:@34194.4]
  assign x622_x533_D17_number = RetimeWrapper_104_io_out; // @[package.scala 96:25:@34226.4 package.scala 96:25:@34227.4]
  assign x623_x357_sum_D15_number = RetimeWrapper_105_io_out; // @[package.scala 96:25:@34235.4 package.scala 96:25:@34236.4]
  assign x626_x362_sum_D15_number = RetimeWrapper_109_io_out; // @[package.scala 96:25:@34286.4 package.scala 96:25:@34287.4]
  assign x628_x367_sum_D15_number = RetimeWrapper_112_io_out; // @[package.scala 96:25:@34328.4 package.scala 96:25:@34329.4]
  assign io_in_x266_TREADY = _T_211 & _T_213; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 67:22:@31985.4 sm_x469_inr_Foreach_SAMPLER_BOX.scala 69:22:@31993.4]
  assign io_in_x267_TVALID = _T_1599 & io_sigsIn_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 688:22:@34544.4]
  assign io_in_x267_TDATA = {{192'd0}, RetimeWrapper_114_io_out}; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 689:24:@34545.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@31963.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@31975.4]
  assign RetimeWrapper_clock = clock; // @[:@31996.4]
  assign RetimeWrapper_reset = reset; // @[:@31997.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31999.4]
  assign RetimeWrapper_io_in = io_in_x266_TDATA[63:0]; // @[package.scala 94:16:@31998.4]
  assign x301_lb_0_clock = clock; // @[:@32006.4]
  assign x301_lb_0_reset = reset; // @[:@32007.4]
  assign x301_lb_0_io_rPort_11_banks_1 = x561_x529_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@33024.4]
  assign x301_lb_0_io_rPort_11_banks_0 = x579_x533_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33023.4]
  assign x301_lb_0_io_rPort_11_ofs_0 = x357_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33025.4]
  assign x301_lb_0_io_rPort_11_en_0 = _T_841 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33027.4]
  assign x301_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33026.4]
  assign x301_lb_0_io_rPort_10_banks_1 = x576_x531_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33209.4]
  assign x301_lb_0_io_rPort_10_banks_0 = x579_x533_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33208.4]
  assign x301_lb_0_io_rPort_10_ofs_0 = x372_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33210.4]
  assign x301_lb_0_io_rPort_10_en_0 = _T_942 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33212.4]
  assign x301_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33211.4]
  assign x301_lb_0_io_rPort_9_banks_1 = x573_x530_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33151.4]
  assign x301_lb_0_io_rPort_9_banks_0 = x579_x533_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33150.4]
  assign x301_lb_0_io_rPort_9_ofs_0 = x367_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33152.4]
  assign x301_lb_0_io_rPort_9_en_0 = _T_910 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33154.4]
  assign x301_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33153.4]
  assign x301_lb_0_io_rPort_8_banks_1 = x570_x525_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@33093.4]
  assign x301_lb_0_io_rPort_8_banks_0 = x579_x533_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33092.4]
  assign x301_lb_0_io_rPort_8_ofs_0 = x362_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33094.4]
  assign x301_lb_0_io_rPort_8_en_0 = _T_878 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33096.4]
  assign x301_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33095.4]
  assign x301_lb_0_io_rPort_7_banks_1 = x573_x530_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@32765.4]
  assign x301_lb_0_io_rPort_7_banks_0 = x566_x524_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@32764.4]
  assign x301_lb_0_io_rPort_7_ofs_0 = x574_x337_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@32766.4]
  assign x301_lb_0_io_rPort_7_en_0 = _T_644 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@32768.4]
  assign x301_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32767.4]
  assign x301_lb_0_io_rPort_6_banks_1 = x573_x530_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33443.4]
  assign x301_lb_0_io_rPort_6_banks_0 = x589_x538_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33442.4]
  assign x301_lb_0_io_rPort_6_ofs_0 = x393_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33444.4]
  assign x301_lb_0_io_rPort_6_en_0 = _T_1106 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33446.4]
  assign x301_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33445.4]
  assign x301_lb_0_io_rPort_5_banks_1 = x576_x531_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33494.4]
  assign x301_lb_0_io_rPort_5_banks_0 = x589_x538_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33493.4]
  assign x301_lb_0_io_rPort_5_ofs_0 = x398_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33495.4]
  assign x301_lb_0_io_rPort_5_en_0 = _T_1137 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33497.4]
  assign x301_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33496.4]
  assign x301_lb_0_io_rPort_4_banks_1 = x561_x529_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@32567.4]
  assign x301_lb_0_io_rPort_4_banks_0 = x566_x524_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@32566.4]
  assign x301_lb_0_io_rPort_4_ofs_0 = x563_x317_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@32568.4]
  assign x301_lb_0_io_rPort_4_en_0 = _T_508 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@32570.4]
  assign x301_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32569.4]
  assign x301_lb_0_io_rPort_3_banks_1 = x570_x525_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@32642.4]
  assign x301_lb_0_io_rPort_3_banks_0 = x566_x524_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@32641.4]
  assign x301_lb_0_io_rPort_3_ofs_0 = x569_x311_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@32643.4]
  assign x301_lb_0_io_rPort_3_en_0 = _T_553 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@32645.4]
  assign x301_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32644.4]
  assign x301_lb_0_io_rPort_2_banks_1 = x570_x525_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@33394.4]
  assign x301_lb_0_io_rPort_2_banks_0 = x589_x538_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33393.4]
  assign x301_lb_0_io_rPort_2_ofs_0 = x388_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33395.4]
  assign x301_lb_0_io_rPort_2_en_0 = _T_1077 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33397.4]
  assign x301_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33396.4]
  assign x301_lb_0_io_rPort_1_banks_1 = x561_x529_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@33345.4]
  assign x301_lb_0_io_rPort_1_banks_0 = x589_x538_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@33344.4]
  assign x301_lb_0_io_rPort_1_ofs_0 = x383_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@33346.4]
  assign x301_lb_0_io_rPort_1_en_0 = _T_1048 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@33348.4]
  assign x301_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33347.4]
  assign x301_lb_0_io_rPort_0_banks_1 = x576_x531_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@32879.4]
  assign x301_lb_0_io_rPort_0_banks_0 = x566_x524_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@32878.4]
  assign x301_lb_0_io_rPort_0_ofs_0 = x577_x346_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@32880.4]
  assign x301_lb_0_io_rPort_0_en_0 = _T_732 & x564_b298_D9; // @[MemInterfaceType.scala 110:79:@32882.4]
  assign x301_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32881.4]
  assign x301_lb_0_io_wPort_1_banks_1 = x555_x529_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@32444.4]
  assign x301_lb_0_io_wPort_1_banks_0 = x553_x524_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@32443.4]
  assign x301_lb_0_io_wPort_1_ofs_0 = x556_x317_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@32445.4]
  assign x301_lb_0_io_wPort_1_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@32446.4]
  assign x301_lb_0_io_wPort_1_en_0 = _T_443 & x551_b298_D3; // @[MemInterfaceType.scala 93:57:@32448.4]
  assign x301_lb_0_io_wPort_0_banks_1 = x552_x525_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@32342.4]
  assign x301_lb_0_io_wPort_0_banks_0 = x553_x524_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@32341.4]
  assign x301_lb_0_io_wPort_0_ofs_0 = x550_x311_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@32343.4]
  assign x301_lb_0_io_wPort_0_data_0 = RetimeWrapper_7_io_out; // @[MemInterfaceType.scala 90:56:@32344.4]
  assign x301_lb_0_io_wPort_0_en_0 = _T_371 & x551_b298_D3; // @[MemInterfaceType.scala 93:57:@32346.4]
  assign x302_lb2_0_clock = clock; // @[:@32099.4]
  assign x302_lb2_0_reset = reset; // @[:@32100.4]
  assign x302_lb2_0_io_rPort_5_banks_1 = x610_x529_D23_number[2:0]; // @[MemInterfaceType.scala 106:58:@34111.4]
  assign x302_lb2_0_io_rPort_5_banks_0 = x615_x524_D24_number[2:0]; // @[MemInterfaceType.scala 106:58:@34110.4]
  assign x302_lb2_0_io_rPort_5_ofs_0 = x612_x317_sum_D22_number[8:0]; // @[MemInterfaceType.scala 107:54:@34112.4]
  assign x302_lb2_0_io_rPort_5_en_0 = _T_1377 & x613_b298_D24; // @[MemInterfaceType.scala 110:79:@34114.4]
  assign x302_lb2_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34113.4]
  assign x302_lb2_0_io_rPort_4_banks_1 = x620_x530_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@34348.4]
  assign x302_lb2_0_io_rPort_4_banks_0 = x622_x533_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@34347.4]
  assign x302_lb2_0_io_rPort_4_ofs_0 = x628_x367_sum_D15_number[8:0]; // @[MemInterfaceType.scala 107:54:@34349.4]
  assign x302_lb2_0_io_rPort_4_en_0 = _T_1511 & x613_b298_D24; // @[MemInterfaceType.scala 110:79:@34351.4]
  assign x302_lb2_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34350.4]
  assign x302_lb2_0_io_rPort_3_banks_1 = x620_x530_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@34213.4]
  assign x302_lb2_0_io_rPort_3_banks_0 = x615_x524_D24_number[2:0]; // @[MemInterfaceType.scala 106:58:@34212.4]
  assign x302_lb2_0_io_rPort_3_ofs_0 = x621_x337_sum_D16_number[8:0]; // @[MemInterfaceType.scala 107:54:@34214.4]
  assign x302_lb2_0_io_rPort_3_en_0 = _T_1433 & x613_b298_D24; // @[MemInterfaceType.scala 110:79:@34216.4]
  assign x302_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34215.4]
  assign x302_lb2_0_io_rPort_2_banks_1 = x618_x525_D24_number[2:0]; // @[MemInterfaceType.scala 106:58:@34306.4]
  assign x302_lb2_0_io_rPort_2_banks_0 = x622_x533_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@34305.4]
  assign x302_lb2_0_io_rPort_2_ofs_0 = x626_x362_sum_D15_number[8:0]; // @[MemInterfaceType.scala 107:54:@34307.4]
  assign x302_lb2_0_io_rPort_2_en_0 = _T_1486 & x613_b298_D24; // @[MemInterfaceType.scala 110:79:@34309.4]
  assign x302_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34308.4]
  assign x302_lb2_0_io_rPort_1_banks_1 = x618_x525_D24_number[2:0]; // @[MemInterfaceType.scala 106:58:@34162.4]
  assign x302_lb2_0_io_rPort_1_banks_0 = x615_x524_D24_number[2:0]; // @[MemInterfaceType.scala 106:58:@34161.4]
  assign x302_lb2_0_io_rPort_1_ofs_0 = x617_x311_sum_D22_number[8:0]; // @[MemInterfaceType.scala 107:54:@34163.4]
  assign x302_lb2_0_io_rPort_1_en_0 = _T_1405 & x613_b298_D24; // @[MemInterfaceType.scala 110:79:@34165.4]
  assign x302_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34164.4]
  assign x302_lb2_0_io_rPort_0_banks_1 = x610_x529_D23_number[2:0]; // @[MemInterfaceType.scala 106:58:@34264.4]
  assign x302_lb2_0_io_rPort_0_banks_0 = x622_x533_D17_number[2:0]; // @[MemInterfaceType.scala 106:58:@34263.4]
  assign x302_lb2_0_io_rPort_0_ofs_0 = x623_x357_sum_D15_number[8:0]; // @[MemInterfaceType.scala 107:54:@34265.4]
  assign x302_lb2_0_io_rPort_0_en_0 = _T_1461 & x613_b298_D24; // @[MemInterfaceType.scala 110:79:@34267.4]
  assign x302_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34266.4]
  assign x302_lb2_0_io_wPort_1_banks_1 = x608_x529_D22_number[2:0]; // @[MemInterfaceType.scala 88:58:@34035.4]
  assign x302_lb2_0_io_wPort_1_banks_0 = x605_x524_D23_number[2:0]; // @[MemInterfaceType.scala 88:58:@34034.4]
  assign x302_lb2_0_io_wPort_1_ofs_0 = x609_x317_sum_D21_number[8:0]; // @[MemInterfaceType.scala 89:54:@34036.4]
  assign x302_lb2_0_io_wPort_1_data_0 = RetimeWrapper_85_io_out; // @[MemInterfaceType.scala 90:56:@34037.4]
  assign x302_lb2_0_io_wPort_1_en_0 = _T_1341 & x603_b298_D23; // @[MemInterfaceType.scala 93:57:@34039.4]
  assign x302_lb2_0_io_wPort_0_banks_1 = x604_x525_D23_number[2:0]; // @[MemInterfaceType.scala 88:58:@33985.4]
  assign x302_lb2_0_io_wPort_0_banks_0 = x605_x524_D23_number[2:0]; // @[MemInterfaceType.scala 88:58:@33984.4]
  assign x302_lb2_0_io_wPort_0_ofs_0 = x602_x311_sum_D21_number[8:0]; // @[MemInterfaceType.scala 89:54:@33986.4]
  assign x302_lb2_0_io_wPort_0_data_0 = RetimeWrapper_83_io_out; // @[MemInterfaceType.scala 90:56:@33987.4]
  assign x302_lb2_0_io_wPort_0_en_0 = _T_1318 & x603_b298_D23; // @[MemInterfaceType.scala 93:57:@33989.4]
  assign x528_sub_1_clock = clock; // @[:@32226.4]
  assign x528_sub_1_reset = reset; // @[:@32227.4]
  assign x528_sub_1_io_a = _T_302[31:0]; // @[Math.scala 192:17:@32228.4]
  assign x528_sub_1_io_b = _T_305[31:0]; // @[Math.scala 193:17:@32229.4]
  assign x528_sub_1_io_flow = io_in_x267_TREADY; // @[Math.scala 194:20:@32230.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32253.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32254.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32256.4]
  assign RetimeWrapper_1_io_in = _T_330 ? 32'h0 : _T_332; // @[package.scala 94:16:@32255.4]
  assign x311_sum_1_clock = clock; // @[:@32262.4]
  assign x311_sum_1_reset = reset; // @[:@32263.4]
  assign x311_sum_1_io_a = x528_sub_1_io_result; // @[Math.scala 151:17:@32264.4]
  assign x311_sum_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 152:17:@32265.4]
  assign x311_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32266.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32272.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32273.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32275.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32274.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32281.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32282.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32284.4]
  assign RetimeWrapper_3_io_in = x311_sum_1_io_result; // @[package.scala 94:16:@32283.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32290.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32291.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32293.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@32292.4]
  assign RetimeWrapper_5_clock = clock; // @[:@32299.4]
  assign RetimeWrapper_5_reset = reset; // @[:@32300.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32302.4]
  assign RetimeWrapper_5_io_in = $unsigned(_T_272); // @[package.scala 94:16:@32301.4]
  assign RetimeWrapper_6_clock = clock; // @[:@32308.4]
  assign RetimeWrapper_6_reset = reset; // @[:@32309.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32311.4]
  assign RetimeWrapper_6_io_in = $unsigned(_T_260); // @[package.scala 94:16:@32310.4]
  assign RetimeWrapper_7_clock = clock; // @[:@32317.4]
  assign RetimeWrapper_7_reset = reset; // @[:@32318.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32320.4]
  assign RetimeWrapper_7_io_in = x547_x299_D1_0_number[31:0]; // @[package.scala 94:16:@32319.4]
  assign RetimeWrapper_8_clock = clock; // @[:@32328.4]
  assign RetimeWrapper_8_reset = reset; // @[:@32329.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32331.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32330.4]
  assign x313_rdcol_1_clock = clock; // @[:@32351.4]
  assign x313_rdcol_1_reset = reset; // @[:@32352.4]
  assign x313_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@32353.4]
  assign x313_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@32354.4]
  assign x313_rdcol_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32355.4]
  assign x317_sum_1_clock = clock; // @[:@32391.4]
  assign x317_sum_1_reset = reset; // @[:@32392.4]
  assign x317_sum_1_io_a = x528_sub_1_io_result; // @[Math.scala 151:17:@32393.4]
  assign x317_sum_1_io_b = _T_414 ? 32'h0 : _T_416; // @[Math.scala 152:17:@32394.4]
  assign x317_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32395.4]
  assign RetimeWrapper_9_clock = clock; // @[:@32401.4]
  assign RetimeWrapper_9_reset = reset; // @[:@32402.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32404.4]
  assign RetimeWrapper_9_io_in = $unsigned(_T_391); // @[package.scala 94:16:@32403.4]
  assign RetimeWrapper_10_clock = clock; // @[:@32410.4]
  assign RetimeWrapper_10_reset = reset; // @[:@32411.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32413.4]
  assign RetimeWrapper_10_io_in = x317_sum_1_io_result; // @[package.scala 94:16:@32412.4]
  assign RetimeWrapper_11_clock = clock; // @[:@32419.4]
  assign RetimeWrapper_11_reset = reset; // @[:@32420.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32422.4]
  assign RetimeWrapper_11_io_in = x547_x299_D1_0_number[63:32]; // @[package.scala 94:16:@32421.4]
  assign RetimeWrapper_12_clock = clock; // @[:@32430.4]
  assign RetimeWrapper_12_reset = reset; // @[:@32431.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32433.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32432.4]
  assign RetimeWrapper_13_clock = clock; // @[:@32451.4]
  assign RetimeWrapper_13_reset = reset; // @[:@32452.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32454.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@32453.4]
  assign RetimeWrapper_14_clock = clock; // @[:@32467.4]
  assign RetimeWrapper_14_reset = reset; // @[:@32468.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32470.4]
  assign RetimeWrapper_14_io_in = x313_rdcol_1_io_result; // @[package.scala 94:16:@32469.4]
  assign RetimeWrapper_15_clock = clock; // @[:@32483.4]
  assign RetimeWrapper_15_reset = reset; // @[:@32484.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32486.4]
  assign RetimeWrapper_15_io_in = $signed(_T_453) < $signed(32'sh0); // @[package.scala 94:16:@32485.4]
  assign RetimeWrapper_16_clock = clock; // @[:@32498.4]
  assign RetimeWrapper_16_reset = reset; // @[:@32499.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32501.4]
  assign RetimeWrapper_16_io_in = $unsigned(_T_391); // @[package.scala 94:16:@32500.4]
  assign RetimeWrapper_17_clock = clock; // @[:@32507.4]
  assign RetimeWrapper_17_reset = reset; // @[:@32508.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32510.4]
  assign RetimeWrapper_17_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32509.4]
  assign RetimeWrapper_18_clock = clock; // @[:@32516.4]
  assign RetimeWrapper_18_reset = reset; // @[:@32517.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32519.4]
  assign RetimeWrapper_18_io_in = x317_sum_1_io_result; // @[package.scala 94:16:@32518.4]
  assign RetimeWrapper_19_clock = clock; // @[:@32525.4]
  assign RetimeWrapper_19_reset = reset; // @[:@32526.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32528.4]
  assign RetimeWrapper_19_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@32527.4]
  assign RetimeWrapper_20_clock = clock; // @[:@32534.4]
  assign RetimeWrapper_20_reset = reset; // @[:@32535.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32537.4]
  assign RetimeWrapper_20_io_in = ~ x322; // @[package.scala 94:16:@32536.4]
  assign RetimeWrapper_21_clock = clock; // @[:@32543.4]
  assign RetimeWrapper_21_reset = reset; // @[:@32544.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32546.4]
  assign RetimeWrapper_21_io_in = $unsigned(_T_260); // @[package.scala 94:16:@32545.4]
  assign RetimeWrapper_22_clock = clock; // @[:@32555.4]
  assign RetimeWrapper_22_reset = reset; // @[:@32556.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32558.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32557.4]
  assign RetimeWrapper_23_clock = clock; // @[:@32576.4]
  assign RetimeWrapper_23_reset = reset; // @[:@32577.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32579.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@32578.4]
  assign RetimeWrapper_24_clock = clock; // @[:@32600.4]
  assign RetimeWrapper_24_reset = reset; // @[:@32601.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32603.4]
  assign RetimeWrapper_24_io_in = ~ x327; // @[package.scala 94:16:@32602.4]
  assign RetimeWrapper_25_clock = clock; // @[:@32609.4]
  assign RetimeWrapper_25_reset = reset; // @[:@32610.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32612.4]
  assign RetimeWrapper_25_io_in = x311_sum_1_io_result; // @[package.scala 94:16:@32611.4]
  assign RetimeWrapper_26_clock = clock; // @[:@32618.4]
  assign RetimeWrapper_26_reset = reset; // @[:@32619.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32621.4]
  assign RetimeWrapper_26_io_in = $unsigned(_T_272); // @[package.scala 94:16:@32620.4]
  assign RetimeWrapper_27_clock = clock; // @[:@32630.4]
  assign RetimeWrapper_27_reset = reset; // @[:@32631.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32633.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32632.4]
  assign x331_rdcol_1_clock = clock; // @[:@32653.4]
  assign x331_rdcol_1_reset = reset; // @[:@32654.4]
  assign x331_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@32655.4]
  assign x331_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@32656.4]
  assign x331_rdcol_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32657.4]
  assign RetimeWrapper_28_clock = clock; // @[:@32704.4]
  assign RetimeWrapper_28_reset = reset; // @[:@32705.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32707.4]
  assign RetimeWrapper_28_io_in = x528_sub_1_io_result; // @[package.scala 94:16:@32706.4]
  assign x337_sum_1_clock = clock; // @[:@32713.4]
  assign x337_sum_1_reset = reset; // @[:@32714.4]
  assign x337_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@32715.4]
  assign x337_sum_1_io_b = _T_608 ? 32'h0 : _T_610; // @[Math.scala 152:17:@32716.4]
  assign x337_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32717.4]
  assign RetimeWrapper_29_clock = clock; // @[:@32723.4]
  assign RetimeWrapper_29_reset = reset; // @[:@32724.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32726.4]
  assign RetimeWrapper_29_io_in = ~ x333; // @[package.scala 94:16:@32725.4]
  assign RetimeWrapper_30_clock = clock; // @[:@32732.4]
  assign RetimeWrapper_30_reset = reset; // @[:@32733.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32735.4]
  assign RetimeWrapper_30_io_in = $unsigned(_T_585); // @[package.scala 94:16:@32734.4]
  assign RetimeWrapper_31_clock = clock; // @[:@32741.4]
  assign RetimeWrapper_31_reset = reset; // @[:@32742.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32744.4]
  assign RetimeWrapper_31_io_in = x337_sum_1_io_result; // @[package.scala 94:16:@32743.4]
  assign RetimeWrapper_32_clock = clock; // @[:@32753.4]
  assign RetimeWrapper_32_reset = reset; // @[:@32754.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32756.4]
  assign RetimeWrapper_32_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32755.4]
  assign x340_rdcol_1_clock = clock; // @[:@32776.4]
  assign x340_rdcol_1_reset = reset; // @[:@32777.4]
  assign x340_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@32778.4]
  assign x340_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@32779.4]
  assign x340_rdcol_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32780.4]
  assign x346_sum_1_clock = clock; // @[:@32827.4]
  assign x346_sum_1_reset = reset; // @[:@32828.4]
  assign x346_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@32829.4]
  assign x346_sum_1_io_b = _T_699 ? 32'h0 : _T_701; // @[Math.scala 152:17:@32830.4]
  assign x346_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32831.4]
  assign RetimeWrapper_33_clock = clock; // @[:@32837.4]
  assign RetimeWrapper_33_reset = reset; // @[:@32838.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32840.4]
  assign RetimeWrapper_33_io_in = ~ x342; // @[package.scala 94:16:@32839.4]
  assign RetimeWrapper_34_clock = clock; // @[:@32846.4]
  assign RetimeWrapper_34_reset = reset; // @[:@32847.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32849.4]
  assign RetimeWrapper_34_io_in = $unsigned(_T_676); // @[package.scala 94:16:@32848.4]
  assign RetimeWrapper_35_clock = clock; // @[:@32855.4]
  assign RetimeWrapper_35_reset = reset; // @[:@32856.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32858.4]
  assign RetimeWrapper_35_io_in = x346_sum_1_io_result; // @[package.scala 94:16:@32857.4]
  assign RetimeWrapper_36_clock = clock; // @[:@32867.4]
  assign RetimeWrapper_36_reset = reset; // @[:@32868.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32870.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32869.4]
  assign x349_rdrow_1_clock = clock; // @[:@32890.4]
  assign x349_rdrow_1_reset = reset; // @[:@32891.4]
  assign x349_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@32892.4]
  assign x349_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@32893.4]
  assign x349_rdrow_1_io_flow = io_in_x267_TREADY; // @[Math.scala 194:20:@32894.4]
  assign x536_sub_1_clock = clock; // @[:@32962.4]
  assign x536_sub_1_reset = reset; // @[:@32963.4]
  assign x536_sub_1_io_a = _T_806[31:0]; // @[Math.scala 192:17:@32964.4]
  assign x536_sub_1_io_b = _T_809[31:0]; // @[Math.scala 193:17:@32965.4]
  assign x536_sub_1_io_flow = io_in_x267_TREADY; // @[Math.scala 194:20:@32966.4]
  assign RetimeWrapper_37_clock = clock; // @[:@32972.4]
  assign RetimeWrapper_37_reset = reset; // @[:@32973.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32975.4]
  assign RetimeWrapper_37_io_in = _T_414 ? 32'h0 : _T_416; // @[package.scala 94:16:@32974.4]
  assign x357_sum_1_clock = clock; // @[:@32981.4]
  assign x357_sum_1_reset = reset; // @[:@32982.4]
  assign x357_sum_1_io_a = x536_sub_1_io_result; // @[Math.scala 151:17:@32983.4]
  assign x357_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@32984.4]
  assign x357_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@32985.4]
  assign RetimeWrapper_38_clock = clock; // @[:@32991.4]
  assign RetimeWrapper_38_reset = reset; // @[:@32992.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32994.4]
  assign RetimeWrapper_38_io_in = $unsigned(_T_776); // @[package.scala 94:16:@32993.4]
  assign RetimeWrapper_39_clock = clock; // @[:@33000.4]
  assign RetimeWrapper_39_reset = reset; // @[:@33001.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33003.4]
  assign RetimeWrapper_39_io_in = ~ x352; // @[package.scala 94:16:@33002.4]
  assign RetimeWrapper_40_clock = clock; // @[:@33012.4]
  assign RetimeWrapper_40_reset = reset; // @[:@33013.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33015.4]
  assign RetimeWrapper_40_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33014.4]
  assign RetimeWrapper_41_clock = clock; // @[:@33033.4]
  assign RetimeWrapper_41_reset = reset; // @[:@33034.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33036.4]
  assign RetimeWrapper_41_io_in = $signed(_T_521) < $signed(32'sh0); // @[package.scala 94:16:@33035.4]
  assign RetimeWrapper_42_clock = clock; // @[:@33048.4]
  assign RetimeWrapper_42_reset = reset; // @[:@33049.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33051.4]
  assign RetimeWrapper_42_io_in = _T_330 ? 32'h0 : _T_332; // @[package.scala 94:16:@33050.4]
  assign x362_sum_1_clock = clock; // @[:@33059.4]
  assign x362_sum_1_reset = reset; // @[:@33060.4]
  assign x362_sum_1_io_a = x536_sub_1_io_result; // @[Math.scala 151:17:@33061.4]
  assign x362_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@33062.4]
  assign x362_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33063.4]
  assign RetimeWrapper_43_clock = clock; // @[:@33069.4]
  assign RetimeWrapper_43_reset = reset; // @[:@33070.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33072.4]
  assign RetimeWrapper_43_io_in = ~ x360; // @[package.scala 94:16:@33071.4]
  assign RetimeWrapper_44_clock = clock; // @[:@33081.4]
  assign RetimeWrapper_44_reset = reset; // @[:@33082.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33084.4]
  assign RetimeWrapper_44_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33083.4]
  assign RetimeWrapper_45_clock = clock; // @[:@33108.4]
  assign RetimeWrapper_45_reset = reset; // @[:@33109.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33111.4]
  assign RetimeWrapper_45_io_in = _T_608 ? 32'h0 : _T_610; // @[package.scala 94:16:@33110.4]
  assign x367_sum_1_clock = clock; // @[:@33117.4]
  assign x367_sum_1_reset = reset; // @[:@33118.4]
  assign x367_sum_1_io_a = x536_sub_1_io_result; // @[Math.scala 151:17:@33119.4]
  assign x367_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@33120.4]
  assign x367_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33121.4]
  assign RetimeWrapper_46_clock = clock; // @[:@33127.4]
  assign RetimeWrapper_46_reset = reset; // @[:@33128.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33130.4]
  assign RetimeWrapper_46_io_in = ~ x365; // @[package.scala 94:16:@33129.4]
  assign RetimeWrapper_47_clock = clock; // @[:@33139.4]
  assign RetimeWrapper_47_reset = reset; // @[:@33140.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33142.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33141.4]
  assign RetimeWrapper_48_clock = clock; // @[:@33166.4]
  assign RetimeWrapper_48_reset = reset; // @[:@33167.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33169.4]
  assign RetimeWrapper_48_io_in = _T_699 ? 32'h0 : _T_701; // @[package.scala 94:16:@33168.4]
  assign x372_sum_1_clock = clock; // @[:@33175.4]
  assign x372_sum_1_reset = reset; // @[:@33176.4]
  assign x372_sum_1_io_a = x536_sub_1_io_result; // @[Math.scala 151:17:@33177.4]
  assign x372_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@33178.4]
  assign x372_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33179.4]
  assign RetimeWrapper_49_clock = clock; // @[:@33185.4]
  assign RetimeWrapper_49_reset = reset; // @[:@33186.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33188.4]
  assign RetimeWrapper_49_io_in = ~ x370; // @[package.scala 94:16:@33187.4]
  assign RetimeWrapper_50_clock = clock; // @[:@33197.4]
  assign RetimeWrapper_50_reset = reset; // @[:@33198.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33200.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33199.4]
  assign x375_rdrow_1_clock = clock; // @[:@33220.4]
  assign x375_rdrow_1_reset = reset; // @[:@33221.4]
  assign x375_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@33222.4]
  assign x375_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@33223.4]
  assign x375_rdrow_1_io_flow = io_in_x267_TREADY; // @[Math.scala 194:20:@33224.4]
  assign x541_sub_1_clock = clock; // @[:@33292.4]
  assign x541_sub_1_reset = reset; // @[:@33293.4]
  assign x541_sub_1_io_a = _T_1016[31:0]; // @[Math.scala 192:17:@33294.4]
  assign x541_sub_1_io_b = _T_1019[31:0]; // @[Math.scala 193:17:@33295.4]
  assign x541_sub_1_io_flow = io_in_x267_TREADY; // @[Math.scala 194:20:@33296.4]
  assign x383_sum_1_clock = clock; // @[:@33302.4]
  assign x383_sum_1_reset = reset; // @[:@33303.4]
  assign x383_sum_1_io_a = x541_sub_1_io_result; // @[Math.scala 151:17:@33304.4]
  assign x383_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@33305.4]
  assign x383_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33306.4]
  assign RetimeWrapper_51_clock = clock; // @[:@33312.4]
  assign RetimeWrapper_51_reset = reset; // @[:@33313.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33315.4]
  assign RetimeWrapper_51_io_in = ~ x378; // @[package.scala 94:16:@33314.4]
  assign RetimeWrapper_52_clock = clock; // @[:@33321.4]
  assign RetimeWrapper_52_reset = reset; // @[:@33322.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33324.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_986); // @[package.scala 94:16:@33323.4]
  assign RetimeWrapper_53_clock = clock; // @[:@33333.4]
  assign RetimeWrapper_53_reset = reset; // @[:@33334.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33336.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33335.4]
  assign x388_sum_1_clock = clock; // @[:@33360.4]
  assign x388_sum_1_reset = reset; // @[:@33361.4]
  assign x388_sum_1_io_a = x541_sub_1_io_result; // @[Math.scala 151:17:@33362.4]
  assign x388_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@33363.4]
  assign x388_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33364.4]
  assign RetimeWrapper_54_clock = clock; // @[:@33370.4]
  assign RetimeWrapper_54_reset = reset; // @[:@33371.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33373.4]
  assign RetimeWrapper_54_io_in = ~ x386; // @[package.scala 94:16:@33372.4]
  assign RetimeWrapper_55_clock = clock; // @[:@33382.4]
  assign RetimeWrapper_55_reset = reset; // @[:@33383.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33385.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33384.4]
  assign x393_sum_1_clock = clock; // @[:@33409.4]
  assign x393_sum_1_reset = reset; // @[:@33410.4]
  assign x393_sum_1_io_a = x541_sub_1_io_result; // @[Math.scala 151:17:@33411.4]
  assign x393_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@33412.4]
  assign x393_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33413.4]
  assign RetimeWrapper_56_clock = clock; // @[:@33419.4]
  assign RetimeWrapper_56_reset = reset; // @[:@33420.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33422.4]
  assign RetimeWrapper_56_io_in = ~ x391; // @[package.scala 94:16:@33421.4]
  assign RetimeWrapper_57_clock = clock; // @[:@33431.4]
  assign RetimeWrapper_57_reset = reset; // @[:@33432.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33434.4]
  assign RetimeWrapper_57_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33433.4]
  assign x398_sum_1_clock = clock; // @[:@33460.4]
  assign x398_sum_1_reset = reset; // @[:@33461.4]
  assign x398_sum_1_io_a = x541_sub_1_io_result; // @[Math.scala 151:17:@33462.4]
  assign x398_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@33463.4]
  assign x398_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33464.4]
  assign RetimeWrapper_58_clock = clock; // @[:@33470.4]
  assign RetimeWrapper_58_reset = reset; // @[:@33471.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33473.4]
  assign RetimeWrapper_58_io_in = ~ x396; // @[package.scala 94:16:@33472.4]
  assign RetimeWrapper_59_clock = clock; // @[:@33482.4]
  assign RetimeWrapper_59_reset = reset; // @[:@33483.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33485.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33484.4]
  assign RetimeWrapper_60_clock = clock; // @[:@33505.4]
  assign RetimeWrapper_60_reset = reset; // @[:@33506.4]
  assign RetimeWrapper_60_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33508.4]
  assign RetimeWrapper_60_io_in = _GEN_6 << 1; // @[package.scala 94:16:@33507.4]
  assign RetimeWrapper_61_clock = clock; // @[:@33517.4]
  assign RetimeWrapper_61_reset = reset; // @[:@33518.4]
  assign RetimeWrapper_61_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33520.4]
  assign RetimeWrapper_61_io_in = _GEN_7 << 1; // @[package.scala 94:16:@33519.4]
  assign RetimeWrapper_62_clock = clock; // @[:@33529.4]
  assign RetimeWrapper_62_reset = reset; // @[:@33530.4]
  assign RetimeWrapper_62_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33532.4]
  assign RetimeWrapper_62_io_in = _GEN_8 << 2; // @[package.scala 94:16:@33531.4]
  assign RetimeWrapper_63_clock = clock; // @[:@33541.4]
  assign RetimeWrapper_63_reset = reset; // @[:@33542.4]
  assign RetimeWrapper_63_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33544.4]
  assign RetimeWrapper_63_io_in = _GEN_9 << 1; // @[package.scala 94:16:@33543.4]
  assign RetimeWrapper_64_clock = clock; // @[:@33553.4]
  assign RetimeWrapper_64_reset = reset; // @[:@33554.4]
  assign RetimeWrapper_64_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33556.4]
  assign RetimeWrapper_64_io_in = _GEN_10 << 1; // @[package.scala 94:16:@33555.4]
  assign RetimeWrapper_65_clock = clock; // @[:@33563.4]
  assign RetimeWrapper_65_reset = reset; // @[:@33564.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33566.4]
  assign RetimeWrapper_65_io_in = x301_lb_0_io_rPort_4_output_0; // @[package.scala 94:16:@33565.4]
  assign x406_x7_1_clock = clock; // @[:@33572.4]
  assign x406_x7_1_reset = reset; // @[:@33573.4]
  assign x406_x7_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@33574.4]
  assign x406_x7_1_io_b = _T_1144[31:0]; // @[Math.scala 152:17:@33575.4]
  assign x406_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33576.4]
  assign RetimeWrapper_66_clock = clock; // @[:@33582.4]
  assign RetimeWrapper_66_reset = reset; // @[:@33583.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33585.4]
  assign RetimeWrapper_66_io_in = x301_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@33584.4]
  assign x407_x8_1_clock = clock; // @[:@33591.4]
  assign x407_x8_1_reset = reset; // @[:@33592.4]
  assign x407_x8_1_io_a = RetimeWrapper_66_io_out; // @[Math.scala 151:17:@33593.4]
  assign x407_x8_1_io_b = _T_1149[31:0]; // @[Math.scala 152:17:@33594.4]
  assign x407_x8_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33595.4]
  assign x408_x7_1_clock = clock; // @[:@33601.4]
  assign x408_x7_1_reset = reset; // @[:@33602.4]
  assign x408_x7_1_io_a = _T_1154[31:0]; // @[Math.scala 151:17:@33603.4]
  assign x408_x7_1_io_b = _T_1159[31:0]; // @[Math.scala 152:17:@33604.4]
  assign x408_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33605.4]
  assign RetimeWrapper_67_clock = clock; // @[:@33611.4]
  assign RetimeWrapper_67_reset = reset; // @[:@33612.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33614.4]
  assign RetimeWrapper_67_io_in = x301_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@33613.4]
  assign x409_x8_1_clock = clock; // @[:@33620.4]
  assign x409_x8_1_reset = reset; // @[:@33621.4]
  assign x409_x8_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@33622.4]
  assign x409_x8_1_io_b = _T_1164[31:0]; // @[Math.scala 152:17:@33623.4]
  assign x409_x8_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33624.4]
  assign x410_x7_1_clock = clock; // @[:@33630.4]
  assign x410_x7_1_reset = reset; // @[:@33631.4]
  assign x410_x7_1_io_a = x406_x7_1_io_result; // @[Math.scala 151:17:@33632.4]
  assign x410_x7_1_io_b = x407_x8_1_io_result; // @[Math.scala 152:17:@33633.4]
  assign x410_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33634.4]
  assign x411_x8_1_clock = clock; // @[:@33640.4]
  assign x411_x8_1_reset = reset; // @[:@33641.4]
  assign x411_x8_1_io_a = x408_x7_1_io_result; // @[Math.scala 151:17:@33642.4]
  assign x411_x8_1_io_b = x409_x8_1_io_result; // @[Math.scala 152:17:@33643.4]
  assign x411_x8_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33644.4]
  assign x412_x7_1_clock = clock; // @[:@33650.4]
  assign x412_x7_1_reset = reset; // @[:@33651.4]
  assign x412_x7_1_io_a = x410_x7_1_io_result; // @[Math.scala 151:17:@33652.4]
  assign x412_x7_1_io_b = x411_x8_1_io_result; // @[Math.scala 152:17:@33653.4]
  assign x412_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33654.4]
  assign RetimeWrapper_68_clock = clock; // @[:@33660.4]
  assign RetimeWrapper_68_reset = reset; // @[:@33661.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33663.4]
  assign RetimeWrapper_68_io_in = x301_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@33662.4]
  assign x413_sum_1_clock = clock; // @[:@33669.4]
  assign x413_sum_1_reset = reset; // @[:@33670.4]
  assign x413_sum_1_io_a = x412_x7_1_io_result; // @[Math.scala 151:17:@33671.4]
  assign x413_sum_1_io_b = RetimeWrapper_68_io_out; // @[Math.scala 152:17:@33672.4]
  assign x413_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33673.4]
  assign x414_1_io_b = x413_sum_1_io_result; // @[Math.scala 721:17:@33681.4]
  assign x415_mul_1_clock = clock; // @[:@33690.4]
  assign x415_mul_1_io_a = x414_1_io_result; // @[Math.scala 263:17:@33692.4]
  assign x415_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@33693.4]
  assign x415_mul_1_io_flow = io_in_x267_TREADY; // @[Math.scala 265:20:@33694.4]
  assign x416_1_io_b = x415_mul_1_io_result; // @[Math.scala 721:17:@33702.4]
  assign RetimeWrapper_69_clock = clock; // @[:@33711.4]
  assign RetimeWrapper_69_reset = reset; // @[:@33712.4]
  assign RetimeWrapper_69_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33714.4]
  assign RetimeWrapper_69_io_in = _GEN_11 << 1; // @[package.scala 94:16:@33713.4]
  assign RetimeWrapper_70_clock = clock; // @[:@33723.4]
  assign RetimeWrapper_70_reset = reset; // @[:@33724.4]
  assign RetimeWrapper_70_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33726.4]
  assign RetimeWrapper_70_io_in = _GEN_12 << 1; // @[package.scala 94:16:@33725.4]
  assign RetimeWrapper_71_clock = clock; // @[:@33735.4]
  assign RetimeWrapper_71_reset = reset; // @[:@33736.4]
  assign RetimeWrapper_71_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33738.4]
  assign RetimeWrapper_71_io_in = _GEN_13 << 2; // @[package.scala 94:16:@33737.4]
  assign RetimeWrapper_72_clock = clock; // @[:@33747.4]
  assign RetimeWrapper_72_reset = reset; // @[:@33748.4]
  assign RetimeWrapper_72_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33750.4]
  assign RetimeWrapper_72_io_in = _GEN_14 << 1; // @[package.scala 94:16:@33749.4]
  assign RetimeWrapper_73_clock = clock; // @[:@33759.4]
  assign RetimeWrapper_73_reset = reset; // @[:@33760.4]
  assign RetimeWrapper_73_io_flow = io_in_x267_TREADY; // @[package.scala 95:18:@33762.4]
  assign RetimeWrapper_73_io_in = _GEN_15 << 1; // @[package.scala 94:16:@33761.4]
  assign RetimeWrapper_74_clock = clock; // @[:@33769.4]
  assign RetimeWrapper_74_reset = reset; // @[:@33770.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33772.4]
  assign RetimeWrapper_74_io_in = x301_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@33771.4]
  assign x422_x7_1_clock = clock; // @[:@33778.4]
  assign x422_x7_1_reset = reset; // @[:@33779.4]
  assign x422_x7_1_io_a = RetimeWrapper_74_io_out; // @[Math.scala 151:17:@33780.4]
  assign x422_x7_1_io_b = _T_1218[31:0]; // @[Math.scala 152:17:@33781.4]
  assign x422_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33782.4]
  assign RetimeWrapper_75_clock = clock; // @[:@33788.4]
  assign RetimeWrapper_75_reset = reset; // @[:@33789.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33791.4]
  assign RetimeWrapper_75_io_in = x301_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@33790.4]
  assign x423_x8_1_clock = clock; // @[:@33797.4]
  assign x423_x8_1_reset = reset; // @[:@33798.4]
  assign x423_x8_1_io_a = RetimeWrapper_75_io_out; // @[Math.scala 151:17:@33799.4]
  assign x423_x8_1_io_b = _T_1223[31:0]; // @[Math.scala 152:17:@33800.4]
  assign x423_x8_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33801.4]
  assign x424_x7_1_clock = clock; // @[:@33807.4]
  assign x424_x7_1_reset = reset; // @[:@33808.4]
  assign x424_x7_1_io_a = _T_1228[31:0]; // @[Math.scala 151:17:@33809.4]
  assign x424_x7_1_io_b = _T_1233[31:0]; // @[Math.scala 152:17:@33810.4]
  assign x424_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33811.4]
  assign RetimeWrapper_76_clock = clock; // @[:@33817.4]
  assign RetimeWrapper_76_reset = reset; // @[:@33818.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33820.4]
  assign RetimeWrapper_76_io_in = x301_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@33819.4]
  assign x425_x8_1_clock = clock; // @[:@33826.4]
  assign x425_x8_1_reset = reset; // @[:@33827.4]
  assign x425_x8_1_io_a = RetimeWrapper_76_io_out; // @[Math.scala 151:17:@33828.4]
  assign x425_x8_1_io_b = _T_1238[31:0]; // @[Math.scala 152:17:@33829.4]
  assign x425_x8_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33830.4]
  assign x426_x7_1_clock = clock; // @[:@33836.4]
  assign x426_x7_1_reset = reset; // @[:@33837.4]
  assign x426_x7_1_io_a = x422_x7_1_io_result; // @[Math.scala 151:17:@33838.4]
  assign x426_x7_1_io_b = x423_x8_1_io_result; // @[Math.scala 152:17:@33839.4]
  assign x426_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33840.4]
  assign x427_x8_1_clock = clock; // @[:@33846.4]
  assign x427_x8_1_reset = reset; // @[:@33847.4]
  assign x427_x8_1_io_a = x424_x7_1_io_result; // @[Math.scala 151:17:@33848.4]
  assign x427_x8_1_io_b = x425_x8_1_io_result; // @[Math.scala 152:17:@33849.4]
  assign x427_x8_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33850.4]
  assign x428_x7_1_clock = clock; // @[:@33856.4]
  assign x428_x7_1_reset = reset; // @[:@33857.4]
  assign x428_x7_1_io_a = x426_x7_1_io_result; // @[Math.scala 151:17:@33858.4]
  assign x428_x7_1_io_b = x427_x8_1_io_result; // @[Math.scala 152:17:@33859.4]
  assign x428_x7_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33860.4]
  assign RetimeWrapper_77_clock = clock; // @[:@33866.4]
  assign RetimeWrapper_77_reset = reset; // @[:@33867.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33869.4]
  assign RetimeWrapper_77_io_in = x301_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@33868.4]
  assign x429_sum_1_clock = clock; // @[:@33875.4]
  assign x429_sum_1_reset = reset; // @[:@33876.4]
  assign x429_sum_1_io_a = x428_x7_1_io_result; // @[Math.scala 151:17:@33877.4]
  assign x429_sum_1_io_b = RetimeWrapper_77_io_out; // @[Math.scala 152:17:@33878.4]
  assign x429_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@33879.4]
  assign x430_1_io_b = x429_sum_1_io_result; // @[Math.scala 721:17:@33887.4]
  assign x431_mul_1_clock = clock; // @[:@33896.4]
  assign x431_mul_1_io_a = x430_1_io_result; // @[Math.scala 263:17:@33898.4]
  assign x431_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@33899.4]
  assign x431_mul_1_io_flow = io_in_x267_TREADY; // @[Math.scala 265:20:@33900.4]
  assign x432_1_io_b = x431_mul_1_io_result; // @[Math.scala 721:17:@33908.4]
  assign RetimeWrapper_78_clock = clock; // @[:@33915.4]
  assign RetimeWrapper_78_reset = reset; // @[:@33916.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33918.4]
  assign RetimeWrapper_78_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33917.4]
  assign RetimeWrapper_79_clock = clock; // @[:@33924.4]
  assign RetimeWrapper_79_reset = reset; // @[:@33925.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33927.4]
  assign RetimeWrapper_79_io_in = x311_sum_1_io_result; // @[package.scala 94:16:@33926.4]
  assign RetimeWrapper_80_clock = clock; // @[:@33933.4]
  assign RetimeWrapper_80_reset = reset; // @[:@33934.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33936.4]
  assign RetimeWrapper_80_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33935.4]
  assign RetimeWrapper_81_clock = clock; // @[:@33942.4]
  assign RetimeWrapper_81_reset = reset; // @[:@33943.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33945.4]
  assign RetimeWrapper_81_io_in = $unsigned(_T_272); // @[package.scala 94:16:@33944.4]
  assign RetimeWrapper_82_clock = clock; // @[:@33951.4]
  assign RetimeWrapper_82_reset = reset; // @[:@33952.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33954.4]
  assign RetimeWrapper_82_io_in = $unsigned(_T_260); // @[package.scala 94:16:@33953.4]
  assign RetimeWrapper_83_clock = clock; // @[:@33960.4]
  assign RetimeWrapper_83_reset = reset; // @[:@33961.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33963.4]
  assign RetimeWrapper_83_io_in = x432_1_io_result; // @[package.scala 94:16:@33962.4]
  assign RetimeWrapper_84_clock = clock; // @[:@33971.4]
  assign RetimeWrapper_84_reset = reset; // @[:@33972.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33974.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33973.4]
  assign RetimeWrapper_85_clock = clock; // @[:@33992.4]
  assign RetimeWrapper_85_reset = reset; // @[:@33993.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33995.4]
  assign RetimeWrapper_85_io_in = x416_1_io_result; // @[package.scala 94:16:@33994.4]
  assign RetimeWrapper_86_clock = clock; // @[:@34001.4]
  assign RetimeWrapper_86_reset = reset; // @[:@34002.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34004.4]
  assign RetimeWrapper_86_io_in = $unsigned(_T_391); // @[package.scala 94:16:@34003.4]
  assign RetimeWrapper_87_clock = clock; // @[:@34010.4]
  assign RetimeWrapper_87_reset = reset; // @[:@34011.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34013.4]
  assign RetimeWrapper_87_io_in = x317_sum_1_io_result; // @[package.scala 94:16:@34012.4]
  assign RetimeWrapper_88_clock = clock; // @[:@34021.4]
  assign RetimeWrapper_88_reset = reset; // @[:@34022.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34024.4]
  assign RetimeWrapper_88_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34023.4]
  assign RetimeWrapper_89_clock = clock; // @[:@34042.4]
  assign RetimeWrapper_89_reset = reset; // @[:@34043.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34045.4]
  assign RetimeWrapper_89_io_in = $unsigned(_T_391); // @[package.scala 94:16:@34044.4]
  assign RetimeWrapper_90_clock = clock; // @[:@34051.4]
  assign RetimeWrapper_90_reset = reset; // @[:@34052.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34054.4]
  assign RetimeWrapper_90_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@34053.4]
  assign RetimeWrapper_91_clock = clock; // @[:@34060.4]
  assign RetimeWrapper_91_reset = reset; // @[:@34061.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34063.4]
  assign RetimeWrapper_91_io_in = x317_sum_1_io_result; // @[package.scala 94:16:@34062.4]
  assign RetimeWrapper_92_clock = clock; // @[:@34069.4]
  assign RetimeWrapper_92_reset = reset; // @[:@34070.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34072.4]
  assign RetimeWrapper_92_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@34071.4]
  assign RetimeWrapper_93_clock = clock; // @[:@34078.4]
  assign RetimeWrapper_93_reset = reset; // @[:@34079.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34081.4]
  assign RetimeWrapper_93_io_in = ~ x322; // @[package.scala 94:16:@34080.4]
  assign RetimeWrapper_94_clock = clock; // @[:@34087.4]
  assign RetimeWrapper_94_reset = reset; // @[:@34088.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34090.4]
  assign RetimeWrapper_94_io_in = $unsigned(_T_260); // @[package.scala 94:16:@34089.4]
  assign RetimeWrapper_95_clock = clock; // @[:@34099.4]
  assign RetimeWrapper_95_reset = reset; // @[:@34100.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34102.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34101.4]
  assign RetimeWrapper_96_clock = clock; // @[:@34120.4]
  assign RetimeWrapper_96_reset = reset; // @[:@34121.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34123.4]
  assign RetimeWrapper_96_io_in = ~ x327; // @[package.scala 94:16:@34122.4]
  assign RetimeWrapper_97_clock = clock; // @[:@34129.4]
  assign RetimeWrapper_97_reset = reset; // @[:@34130.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34132.4]
  assign RetimeWrapper_97_io_in = x311_sum_1_io_result; // @[package.scala 94:16:@34131.4]
  assign RetimeWrapper_98_clock = clock; // @[:@34138.4]
  assign RetimeWrapper_98_reset = reset; // @[:@34139.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34141.4]
  assign RetimeWrapper_98_io_in = $unsigned(_T_272); // @[package.scala 94:16:@34140.4]
  assign RetimeWrapper_99_clock = clock; // @[:@34150.4]
  assign RetimeWrapper_99_reset = reset; // @[:@34151.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34153.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34152.4]
  assign RetimeWrapper_100_clock = clock; // @[:@34171.4]
  assign RetimeWrapper_100_reset = reset; // @[:@34172.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34174.4]
  assign RetimeWrapper_100_io_in = ~ x333; // @[package.scala 94:16:@34173.4]
  assign RetimeWrapper_101_clock = clock; // @[:@34180.4]
  assign RetimeWrapper_101_reset = reset; // @[:@34181.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34183.4]
  assign RetimeWrapper_101_io_in = $unsigned(_T_585); // @[package.scala 94:16:@34182.4]
  assign RetimeWrapper_102_clock = clock; // @[:@34189.4]
  assign RetimeWrapper_102_reset = reset; // @[:@34190.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34192.4]
  assign RetimeWrapper_102_io_in = x337_sum_1_io_result; // @[package.scala 94:16:@34191.4]
  assign RetimeWrapper_103_clock = clock; // @[:@34201.4]
  assign RetimeWrapper_103_reset = reset; // @[:@34202.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34204.4]
  assign RetimeWrapper_103_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34203.4]
  assign RetimeWrapper_104_clock = clock; // @[:@34222.4]
  assign RetimeWrapper_104_reset = reset; // @[:@34223.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34225.4]
  assign RetimeWrapper_104_io_in = $unsigned(_T_776); // @[package.scala 94:16:@34224.4]
  assign RetimeWrapper_105_clock = clock; // @[:@34231.4]
  assign RetimeWrapper_105_reset = reset; // @[:@34232.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34234.4]
  assign RetimeWrapper_105_io_in = x357_sum_1_io_result; // @[package.scala 94:16:@34233.4]
  assign RetimeWrapper_106_clock = clock; // @[:@34240.4]
  assign RetimeWrapper_106_reset = reset; // @[:@34241.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34243.4]
  assign RetimeWrapper_106_io_in = ~ x352; // @[package.scala 94:16:@34242.4]
  assign RetimeWrapper_107_clock = clock; // @[:@34252.4]
  assign RetimeWrapper_107_reset = reset; // @[:@34253.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34255.4]
  assign RetimeWrapper_107_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34254.4]
  assign RetimeWrapper_108_clock = clock; // @[:@34273.4]
  assign RetimeWrapper_108_reset = reset; // @[:@34274.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34276.4]
  assign RetimeWrapper_108_io_in = ~ x360; // @[package.scala 94:16:@34275.4]
  assign RetimeWrapper_109_clock = clock; // @[:@34282.4]
  assign RetimeWrapper_109_reset = reset; // @[:@34283.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34285.4]
  assign RetimeWrapper_109_io_in = x362_sum_1_io_result; // @[package.scala 94:16:@34284.4]
  assign RetimeWrapper_110_clock = clock; // @[:@34294.4]
  assign RetimeWrapper_110_reset = reset; // @[:@34295.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34297.4]
  assign RetimeWrapper_110_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34296.4]
  assign RetimeWrapper_111_clock = clock; // @[:@34315.4]
  assign RetimeWrapper_111_reset = reset; // @[:@34316.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34318.4]
  assign RetimeWrapper_111_io_in = ~ x365; // @[package.scala 94:16:@34317.4]
  assign RetimeWrapper_112_clock = clock; // @[:@34324.4]
  assign RetimeWrapper_112_reset = reset; // @[:@34325.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34327.4]
  assign RetimeWrapper_112_io_in = x367_sum_1_io_result; // @[package.scala 94:16:@34326.4]
  assign RetimeWrapper_113_clock = clock; // @[:@34336.4]
  assign RetimeWrapper_113_reset = reset; // @[:@34337.4]
  assign RetimeWrapper_113_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34339.4]
  assign RetimeWrapper_113_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34338.4]
  assign x451_x9_1_clock = clock; // @[:@34369.4]
  assign x451_x9_1_reset = reset; // @[:@34370.4]
  assign x451_x9_1_io_a = x302_lb2_0_io_rPort_5_output_0; // @[Math.scala 151:17:@34371.4]
  assign x451_x9_1_io_b = _T_1518[31:0]; // @[Math.scala 152:17:@34372.4]
  assign x451_x9_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@34373.4]
  assign x452_x10_1_clock = clock; // @[:@34379.4]
  assign x452_x10_1_reset = reset; // @[:@34380.4]
  assign x452_x10_1_io_a = _T_1521[31:0]; // @[Math.scala 151:17:@34381.4]
  assign x452_x10_1_io_b = x302_lb2_0_io_rPort_2_output_0; // @[Math.scala 152:17:@34382.4]
  assign x452_x10_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@34383.4]
  assign x453_sum_1_clock = clock; // @[:@34389.4]
  assign x453_sum_1_reset = reset; // @[:@34390.4]
  assign x453_sum_1_io_a = x451_x9_1_io_result; // @[Math.scala 151:17:@34391.4]
  assign x453_sum_1_io_b = x452_x10_1_io_result; // @[Math.scala 152:17:@34392.4]
  assign x453_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@34393.4]
  assign x454_1_io_b = x453_sum_1_io_result; // @[Math.scala 721:17:@34401.4]
  assign x455_mul_1_clock = clock; // @[:@34410.4]
  assign x455_mul_1_io_a = x454_1_io_result; // @[Math.scala 263:17:@34412.4]
  assign x455_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@34413.4]
  assign x455_mul_1_io_flow = io_in_x267_TREADY; // @[Math.scala 265:20:@34414.4]
  assign x456_1_io_b = x455_mul_1_io_result; // @[Math.scala 721:17:@34424.4]
  assign x459_x9_1_clock = clock; // @[:@34441.4]
  assign x459_x9_1_reset = reset; // @[:@34442.4]
  assign x459_x9_1_io_a = x302_lb2_0_io_rPort_1_output_0; // @[Math.scala 151:17:@34443.4]
  assign x459_x9_1_io_b = _T_1548[31:0]; // @[Math.scala 152:17:@34444.4]
  assign x459_x9_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@34445.4]
  assign x460_x10_1_clock = clock; // @[:@34451.4]
  assign x460_x10_1_reset = reset; // @[:@34452.4]
  assign x460_x10_1_io_a = _T_1551[31:0]; // @[Math.scala 151:17:@34453.4]
  assign x460_x10_1_io_b = x302_lb2_0_io_rPort_4_output_0; // @[Math.scala 152:17:@34454.4]
  assign x460_x10_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@34455.4]
  assign x461_sum_1_clock = clock; // @[:@34461.4]
  assign x461_sum_1_reset = reset; // @[:@34462.4]
  assign x461_sum_1_io_a = x459_x9_1_io_result; // @[Math.scala 151:17:@34463.4]
  assign x461_sum_1_io_b = x460_x10_1_io_result; // @[Math.scala 152:17:@34464.4]
  assign x461_sum_1_io_flow = io_in_x267_TREADY; // @[Math.scala 153:20:@34465.4]
  assign x462_1_io_b = x461_sum_1_io_result; // @[Math.scala 721:17:@34473.4]
  assign x463_mul_1_clock = clock; // @[:@34482.4]
  assign x463_mul_1_io_a = x462_1_io_result; // @[Math.scala 263:17:@34484.4]
  assign x463_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@34485.4]
  assign x463_mul_1_io_flow = io_in_x267_TREADY; // @[Math.scala 265:20:@34486.4]
  assign x464_1_io_b = x463_mul_1_io_result; // @[Math.scala 721:17:@34494.4]
  assign RetimeWrapper_114_clock = clock; // @[:@34507.4]
  assign RetimeWrapper_114_reset = reset; // @[:@34508.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34510.4]
  assign RetimeWrapper_114_io_in = {x456_number,x464_number}; // @[package.scala 94:16:@34509.4]
  assign RetimeWrapper_115_clock = clock; // @[:@34516.4]
  assign RetimeWrapper_115_reset = reset; // @[:@34517.4]
  assign RetimeWrapper_115_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34519.4]
  assign RetimeWrapper_115_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@34518.4]
  assign RetimeWrapper_116_clock = clock; // @[:@34525.4]
  assign RetimeWrapper_116_reset = reset; // @[:@34526.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34528.4]
  assign RetimeWrapper_116_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@34527.4]
  assign RetimeWrapper_117_clock = clock; // @[:@34534.4]
  assign RetimeWrapper_117_reset = reset; // @[:@34535.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34537.4]
  assign RetimeWrapper_117_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34536.4]
endmodule
module x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1( // @[:@34555.2]
  input          clock, // @[:@34556.4]
  input          reset, // @[:@34557.4]
  input          io_in_x266_TVALID, // @[:@34558.4]
  output         io_in_x266_TREADY, // @[:@34558.4]
  input  [255:0] io_in_x266_TDATA, // @[:@34558.4]
  input  [7:0]   io_in_x266_TID, // @[:@34558.4]
  input  [7:0]   io_in_x266_TDEST, // @[:@34558.4]
  output         io_in_x267_TVALID, // @[:@34558.4]
  input          io_in_x267_TREADY, // @[:@34558.4]
  output [255:0] io_in_x267_TDATA, // @[:@34558.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@34558.4]
  input          io_sigsIn_smChildAcks_0, // @[:@34558.4]
  output         io_sigsOut_smDoneIn_0, // @[:@34558.4]
  input          io_rr // @[:@34558.4]
);
  wire  x294_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x294_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x294_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x294_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire [12:0] x294_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire [12:0] x294_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x294_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x294_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x294_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@34592.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34680.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34680.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34680.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34680.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34680.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34722.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34722.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34722.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34722.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34722.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@34730.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@34730.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@34730.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@34730.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@34730.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TREADY; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire [255:0] x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TDATA; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire [7:0] x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TID; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire [7:0] x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TDEST; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TVALID; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TREADY; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire [255:0] x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TDATA; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire [31:0] x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire [31:0] x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
  wire  _T_240; // @[package.scala 96:25:@34685.4 package.scala 96:25:@34686.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x470_outr_UnitPipe.scala 69:66:@34691.4]
  wire  _T_253; // @[package.scala 96:25:@34727.4 package.scala 96:25:@34728.4]
  wire  _T_259; // @[package.scala 96:25:@34735.4 package.scala 96:25:@34736.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@34738.4]
  wire  x469_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@34739.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@34747.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@34748.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@34760.4]
  x274_ctrchain x294_ctrchain ( // @[SpatialBlocks.scala 37:22:@34592.4]
    .clock(x294_ctrchain_clock),
    .reset(x294_ctrchain_reset),
    .io_input_reset(x294_ctrchain_io_input_reset),
    .io_input_enable(x294_ctrchain_io_input_enable),
    .io_output_counts_1(x294_ctrchain_io_output_counts_1),
    .io_output_counts_0(x294_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x294_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x294_ctrchain_io_output_oobs_1),
    .io_output_done(x294_ctrchain_io_output_done)
  );
  x469_inr_Foreach_SAMPLER_BOX_sm x469_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 32:18:@34652.4]
    .clock(x469_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x469_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x469_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x469_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x469_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x469_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x469_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x469_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x469_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34680.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34722.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@34730.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1 x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 701:24:@34764.4]
    .clock(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x266_TREADY(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TREADY),
    .io_in_x266_TDATA(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TDATA),
    .io_in_x266_TID(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TID),
    .io_in_x266_TDEST(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TDEST),
    .io_in_x267_TVALID(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TVALID),
    .io_in_x267_TREADY(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TREADY),
    .io_in_x267_TDATA(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TDATA),
    .io_sigsIn_backpressure(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@34685.4 package.scala 96:25:@34686.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x266_TVALID | x469_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x470_outr_UnitPipe.scala 69:66:@34691.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34727.4 package.scala 96:25:@34728.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@34735.4 package.scala 96:25:@34736.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@34738.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@34739.4]
  assign _T_264 = x469_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@34747.4]
  assign _T_265 = ~ x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@34748.4]
  assign _T_272 = x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@34760.4]
  assign io_in_x266_TREADY = x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TREADY; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 48:23:@34822.4]
  assign io_in_x267_TVALID = x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TVALID; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 49:23:@34832.4]
  assign io_in_x267_TDATA = x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TDATA; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 49:23:@34830.4]
  assign io_sigsOut_smDoneIn_0 = x469_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@34745.4]
  assign x294_ctrchain_clock = clock; // @[:@34593.4]
  assign x294_ctrchain_reset = reset; // @[:@34594.4]
  assign x294_ctrchain_io_input_reset = x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@34763.4]
  assign x294_ctrchain_io_input_enable = _T_272 & x469_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@34715.4 SpatialBlocks.scala 159:42:@34762.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@34653.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@34654.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_io_enable = x469_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x469_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@34742.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x470_outr_UnitPipe.scala 67:50:@34688.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@34744.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x267_TREADY | x469_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@34716.4]
  assign x469_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x470_outr_UnitPipe.scala 71:48:@34694.4]
  assign RetimeWrapper_clock = clock; // @[:@34681.4]
  assign RetimeWrapper_reset = reset; // @[:@34682.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34684.4]
  assign RetimeWrapper_io_in = x294_ctrchain_io_output_done; // @[package.scala 94:16:@34683.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34723.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34724.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34726.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@34725.4]
  assign RetimeWrapper_2_clock = clock; // @[:@34731.4]
  assign RetimeWrapper_2_reset = reset; // @[:@34732.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@34734.4]
  assign RetimeWrapper_2_io_in = x469_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@34733.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@34765.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@34766.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TDATA = io_in_x266_TDATA; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 48:23:@34821.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TID = io_in_x266_TID; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 48:23:@34817.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x266_TDEST = io_in_x266_TDEST; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 48:23:@34816.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x267_TREADY = io_in_x267_TREADY; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 49:23:@34831.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x267_TREADY | x469_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34849.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34847.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x469_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34845.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x294_ctrchain_io_output_counts_1[12]}},x294_ctrchain_io_output_counts_1}; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34840.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x294_ctrchain_io_output_counts_0[12]}},x294_ctrchain_io_output_counts_0}; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34839.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x294_ctrchain_io_output_oobs_0; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34837.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x294_ctrchain_io_output_oobs_1; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 706:22:@34838.4]
  assign x469_inr_Foreach_SAMPLER_BOX_kernelx469_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x469_inr_Foreach_SAMPLER_BOX.scala 705:18:@34833.4]
endmodule
module x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1( // @[:@34863.2]
  input          clock, // @[:@34864.4]
  input          reset, // @[:@34865.4]
  input          io_in_x266_TVALID, // @[:@34866.4]
  output         io_in_x266_TREADY, // @[:@34866.4]
  input  [255:0] io_in_x266_TDATA, // @[:@34866.4]
  input  [7:0]   io_in_x266_TID, // @[:@34866.4]
  input  [7:0]   io_in_x266_TDEST, // @[:@34866.4]
  output         io_in_x267_TVALID, // @[:@34866.4]
  input          io_in_x267_TREADY, // @[:@34866.4]
  output [255:0] io_in_x267_TDATA, // @[:@34866.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@34866.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@34866.4]
  input          io_sigsIn_smChildAcks_0, // @[:@34866.4]
  input          io_sigsIn_smChildAcks_1, // @[:@34866.4]
  output         io_sigsOut_smDoneIn_0, // @[:@34866.4]
  output         io_sigsOut_smDoneIn_1, // @[:@34866.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@34866.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@34866.4]
  input          io_rr // @[:@34866.4]
);
  wire  x269_fifoinraw_0_clock; // @[m_x269_fifoinraw_0.scala 27:17:@34880.4]
  wire  x269_fifoinraw_0_reset; // @[m_x269_fifoinraw_0.scala 27:17:@34880.4]
  wire  x270_fifoinpacked_0_clock; // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
  wire  x270_fifoinpacked_0_reset; // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
  wire  x270_fifoinpacked_0_io_wPort_0_en_0; // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
  wire  x270_fifoinpacked_0_io_full; // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
  wire  x270_fifoinpacked_0_io_active_0_in; // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
  wire  x270_fifoinpacked_0_io_active_0_out; // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
  wire  x271_fifooutraw_0_clock; // @[m_x271_fifooutraw_0.scala 27:17:@34928.4]
  wire  x271_fifooutraw_0_reset; // @[m_x271_fifooutraw_0.scala 27:17:@34928.4]
  wire  x274_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x274_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x274_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x274_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire [12:0] x274_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire [12:0] x274_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x274_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x274_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x274_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@34952.4]
  wire  x290_inr_Foreach_sm_clock; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_reset; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_enable; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_done; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_doneLatch; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_ctrDone; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_datapathEn; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_ctrInc; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_ctrRst; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_parentAck; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_backpressure; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  x290_inr_Foreach_sm_io_break; // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@35040.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@35086.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@35086.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@35086.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@35086.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@35086.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@35094.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@35094.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_clock; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_reset; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_wPort_0_en_0; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_full; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_active_0_in; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_active_0_out; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire [31:0] x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire [31:0] x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_rr; // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
  wire  x470_outr_UnitPipe_sm_clock; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_reset; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_enable; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_done; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_rst; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_ctrDone; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_ctrInc; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_parentAck; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  x470_outr_UnitPipe_sm_io_childAck_0; // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@35318.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@35318.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@35318.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@35318.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@35318.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@35326.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@35326.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@35326.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@35326.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@35326.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_clock; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_reset; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TVALID; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TREADY; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire [255:0] x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TDATA; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire [7:0] x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TID; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire [7:0] x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TDEST; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TVALID; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TREADY; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire [255:0] x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TDATA; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_rr; // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
  wire  _T_254; // @[package.scala 96:25:@35045.4 package.scala 96:25:@35046.4]
  wire  _T_260; // @[implicits.scala 47:10:@35049.4]
  wire  _T_261; // @[sm_x471_outr_UnitPipe.scala 70:41:@35050.4]
  wire  _T_262; // @[sm_x471_outr_UnitPipe.scala 70:78:@35051.4]
  wire  _T_263; // @[sm_x471_outr_UnitPipe.scala 70:76:@35052.4]
  wire  _T_275; // @[package.scala 96:25:@35091.4 package.scala 96:25:@35092.4]
  wire  _T_281; // @[package.scala 96:25:@35099.4 package.scala 96:25:@35100.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@35102.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@35111.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@35112.4]
  wire  _T_354; // @[package.scala 100:49:@35289.4]
  reg  _T_357; // @[package.scala 48:56:@35290.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@35323.4 package.scala 96:25:@35324.4]
  wire  _T_377; // @[package.scala 96:25:@35331.4 package.scala 96:25:@35332.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@35334.4]
  x269_fifoinraw_0 x269_fifoinraw_0 ( // @[m_x269_fifoinraw_0.scala 27:17:@34880.4]
    .clock(x269_fifoinraw_0_clock),
    .reset(x269_fifoinraw_0_reset)
  );
  x270_fifoinpacked_0 x270_fifoinpacked_0 ( // @[m_x270_fifoinpacked_0.scala 27:17:@34904.4]
    .clock(x270_fifoinpacked_0_clock),
    .reset(x270_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x270_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x270_fifoinpacked_0_io_full),
    .io_active_0_in(x270_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x270_fifoinpacked_0_io_active_0_out)
  );
  x269_fifoinraw_0 x271_fifooutraw_0 ( // @[m_x271_fifooutraw_0.scala 27:17:@34928.4]
    .clock(x271_fifooutraw_0_clock),
    .reset(x271_fifooutraw_0_reset)
  );
  x274_ctrchain x274_ctrchain ( // @[SpatialBlocks.scala 37:22:@34952.4]
    .clock(x274_ctrchain_clock),
    .reset(x274_ctrchain_reset),
    .io_input_reset(x274_ctrchain_io_input_reset),
    .io_input_enable(x274_ctrchain_io_input_enable),
    .io_output_counts_1(x274_ctrchain_io_output_counts_1),
    .io_output_counts_0(x274_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x274_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x274_ctrchain_io_output_oobs_1),
    .io_output_done(x274_ctrchain_io_output_done)
  );
  x290_inr_Foreach_sm x290_inr_Foreach_sm ( // @[sm_x290_inr_Foreach.scala 32:18:@35012.4]
    .clock(x290_inr_Foreach_sm_clock),
    .reset(x290_inr_Foreach_sm_reset),
    .io_enable(x290_inr_Foreach_sm_io_enable),
    .io_done(x290_inr_Foreach_sm_io_done),
    .io_doneLatch(x290_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x290_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x290_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x290_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x290_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x290_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x290_inr_Foreach_sm_io_backpressure),
    .io_break(x290_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@35040.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@35086.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@35094.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x290_inr_Foreach_kernelx290_inr_Foreach_concrete1 x290_inr_Foreach_kernelx290_inr_Foreach_concrete1 ( // @[sm_x290_inr_Foreach.scala 98:24:@35129.4]
    .clock(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_clock),
    .reset(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_reset),
    .io_in_x270_fifoinpacked_0_wPort_0_en_0(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_wPort_0_en_0),
    .io_in_x270_fifoinpacked_0_full(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_full),
    .io_in_x270_fifoinpacked_0_active_0_in(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_active_0_in),
    .io_in_x270_fifoinpacked_0_active_0_out(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x470_outr_UnitPipe_sm ( // @[sm_x470_outr_UnitPipe.scala 32:18:@35261.4]
    .clock(x470_outr_UnitPipe_sm_clock),
    .reset(x470_outr_UnitPipe_sm_reset),
    .io_enable(x470_outr_UnitPipe_sm_io_enable),
    .io_done(x470_outr_UnitPipe_sm_io_done),
    .io_rst(x470_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x470_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x470_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x470_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x470_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x470_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x470_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@35318.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@35326.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1 x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1 ( // @[sm_x470_outr_UnitPipe.scala 76:24:@35356.4]
    .clock(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_clock),
    .reset(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_reset),
    .io_in_x266_TVALID(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TVALID),
    .io_in_x266_TREADY(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TREADY),
    .io_in_x266_TDATA(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TDATA),
    .io_in_x266_TID(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TID),
    .io_in_x266_TDEST(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TDEST),
    .io_in_x267_TVALID(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TVALID),
    .io_in_x267_TREADY(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TREADY),
    .io_in_x267_TDATA(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TDATA),
    .io_sigsIn_smEnableOuts_0(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@35045.4 package.scala 96:25:@35046.4]
  assign _T_260 = x270_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@35049.4]
  assign _T_261 = ~ _T_260; // @[sm_x471_outr_UnitPipe.scala 70:41:@35050.4]
  assign _T_262 = ~ x270_fifoinpacked_0_io_active_0_out; // @[sm_x471_outr_UnitPipe.scala 70:78:@35051.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x471_outr_UnitPipe.scala 70:76:@35052.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@35091.4 package.scala 96:25:@35092.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@35099.4 package.scala 96:25:@35100.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@35102.4]
  assign _T_286 = x290_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@35111.4]
  assign _T_287 = ~ x290_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@35112.4]
  assign _T_354 = x470_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@35289.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@35323.4 package.scala 96:25:@35324.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@35331.4 package.scala 96:25:@35332.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@35334.4]
  assign io_in_x266_TREADY = x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TREADY; // @[sm_x470_outr_UnitPipe.scala 48:23:@35412.4]
  assign io_in_x267_TVALID = x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TVALID; // @[sm_x470_outr_UnitPipe.scala 49:23:@35422.4]
  assign io_in_x267_TDATA = x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TDATA; // @[sm_x470_outr_UnitPipe.scala 49:23:@35420.4]
  assign io_sigsOut_smDoneIn_0 = x290_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@35109.4]
  assign io_sigsOut_smDoneIn_1 = x470_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@35341.4]
  assign io_sigsOut_smCtrCopyDone_0 = x290_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@35128.4]
  assign io_sigsOut_smCtrCopyDone_1 = x470_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@35355.4]
  assign x269_fifoinraw_0_clock = clock; // @[:@34881.4]
  assign x269_fifoinraw_0_reset = reset; // @[:@34882.4]
  assign x270_fifoinpacked_0_clock = clock; // @[:@34905.4]
  assign x270_fifoinpacked_0_reset = reset; // @[:@34906.4]
  assign x270_fifoinpacked_0_io_wPort_0_en_0 = x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@35189.4]
  assign x270_fifoinpacked_0_io_active_0_in = x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@35188.4]
  assign x271_fifooutraw_0_clock = clock; // @[:@34929.4]
  assign x271_fifooutraw_0_reset = reset; // @[:@34930.4]
  assign x274_ctrchain_clock = clock; // @[:@34953.4]
  assign x274_ctrchain_reset = reset; // @[:@34954.4]
  assign x274_ctrchain_io_input_reset = x290_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@35127.4]
  assign x274_ctrchain_io_input_enable = x290_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@35079.4 SpatialBlocks.scala 159:42:@35126.4]
  assign x290_inr_Foreach_sm_clock = clock; // @[:@35013.4]
  assign x290_inr_Foreach_sm_reset = reset; // @[:@35014.4]
  assign x290_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@35106.4]
  assign x290_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x471_outr_UnitPipe.scala 69:38:@35048.4]
  assign x290_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@35108.4]
  assign x290_inr_Foreach_sm_io_backpressure = _T_263 | x290_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@35080.4]
  assign x290_inr_Foreach_sm_io_break = 1'h0; // @[sm_x471_outr_UnitPipe.scala 73:36:@35058.4]
  assign RetimeWrapper_clock = clock; // @[:@35041.4]
  assign RetimeWrapper_reset = reset; // @[:@35042.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@35044.4]
  assign RetimeWrapper_io_in = x274_ctrchain_io_output_done; // @[package.scala 94:16:@35043.4]
  assign RetimeWrapper_1_clock = clock; // @[:@35087.4]
  assign RetimeWrapper_1_reset = reset; // @[:@35088.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@35090.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@35089.4]
  assign RetimeWrapper_2_clock = clock; // @[:@35095.4]
  assign RetimeWrapper_2_reset = reset; // @[:@35096.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@35098.4]
  assign RetimeWrapper_2_io_in = x290_inr_Foreach_sm_io_done; // @[package.scala 94:16:@35097.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_clock = clock; // @[:@35130.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_reset = reset; // @[:@35131.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_full = x270_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@35183.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_in_x270_fifoinpacked_0_active_0_out = x270_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@35182.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x290_inr_Foreach_sm_io_doneLatch; // @[sm_x290_inr_Foreach.scala 103:22:@35212.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x290_inr_Foreach.scala 103:22:@35210.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_break = x290_inr_Foreach_sm_io_break; // @[sm_x290_inr_Foreach.scala 103:22:@35208.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x274_ctrchain_io_output_counts_1[12]}},x274_ctrchain_io_output_counts_1}; // @[sm_x290_inr_Foreach.scala 103:22:@35203.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x274_ctrchain_io_output_counts_0[12]}},x274_ctrchain_io_output_counts_0}; // @[sm_x290_inr_Foreach.scala 103:22:@35202.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x274_ctrchain_io_output_oobs_0; // @[sm_x290_inr_Foreach.scala 103:22:@35200.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x274_ctrchain_io_output_oobs_1; // @[sm_x290_inr_Foreach.scala 103:22:@35201.4]
  assign x290_inr_Foreach_kernelx290_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x290_inr_Foreach.scala 102:18:@35196.4]
  assign x470_outr_UnitPipe_sm_clock = clock; // @[:@35262.4]
  assign x470_outr_UnitPipe_sm_reset = reset; // @[:@35263.4]
  assign x470_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@35338.4]
  assign x470_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@35313.4]
  assign x470_outr_UnitPipe_sm_io_ctrDone = x470_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x471_outr_UnitPipe.scala 78:40:@35293.4]
  assign x470_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@35340.4]
  assign x470_outr_UnitPipe_sm_io_doneIn_0 = x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@35310.4]
  assign RetimeWrapper_3_clock = clock; // @[:@35319.4]
  assign RetimeWrapper_3_reset = reset; // @[:@35320.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@35322.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@35321.4]
  assign RetimeWrapper_4_clock = clock; // @[:@35327.4]
  assign RetimeWrapper_4_reset = reset; // @[:@35328.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@35330.4]
  assign RetimeWrapper_4_io_in = x470_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@35329.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_clock = clock; // @[:@35357.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_reset = reset; // @[:@35358.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TVALID = io_in_x266_TVALID; // @[sm_x470_outr_UnitPipe.scala 48:23:@35413.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TDATA = io_in_x266_TDATA; // @[sm_x470_outr_UnitPipe.scala 48:23:@35411.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TID = io_in_x266_TID; // @[sm_x470_outr_UnitPipe.scala 48:23:@35407.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x266_TDEST = io_in_x266_TDEST; // @[sm_x470_outr_UnitPipe.scala 48:23:@35406.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_in_x267_TREADY = io_in_x267_TREADY; // @[sm_x470_outr_UnitPipe.scala 49:23:@35421.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x470_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x470_outr_UnitPipe.scala 81:22:@35431.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x470_outr_UnitPipe_sm_io_childAck_0; // @[sm_x470_outr_UnitPipe.scala 81:22:@35429.4]
  assign x470_outr_UnitPipe_kernelx470_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x470_outr_UnitPipe.scala 80:18:@35423.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x493_outr_UnitPipe_sm( // @[:@35920.2]
  input   clock, // @[:@35921.4]
  input   reset, // @[:@35922.4]
  input   io_enable, // @[:@35923.4]
  output  io_done, // @[:@35923.4]
  input   io_parentAck, // @[:@35923.4]
  input   io_doneIn_0, // @[:@35923.4]
  input   io_doneIn_1, // @[:@35923.4]
  input   io_doneIn_2, // @[:@35923.4]
  output  io_enableOut_0, // @[:@35923.4]
  output  io_enableOut_1, // @[:@35923.4]
  output  io_enableOut_2, // @[:@35923.4]
  output  io_childAck_0, // @[:@35923.4]
  output  io_childAck_1, // @[:@35923.4]
  output  io_childAck_2, // @[:@35923.4]
  input   io_ctrCopyDone_0, // @[:@35923.4]
  input   io_ctrCopyDone_1, // @[:@35923.4]
  input   io_ctrCopyDone_2 // @[:@35923.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@35926.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@35926.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@35926.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@35926.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@35926.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@35926.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@35929.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@35929.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@35929.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@35929.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@35929.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@35929.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@35932.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@35932.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@35932.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@35932.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@35932.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@35932.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@35935.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@35935.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@35935.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@35935.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@35935.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@35935.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@35938.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@35938.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@35938.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@35938.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@35938.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@35938.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@35941.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@35941.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@35941.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@35941.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@35941.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@35941.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@35982.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@35982.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@35982.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@35982.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@35982.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@35982.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@35985.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@35985.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@35985.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@35985.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@35985.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@35985.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@35988.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@35988.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@35988.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@35988.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@35988.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@35988.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36039.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36039.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36039.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36039.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36039.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36053.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36053.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36053.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36053.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36053.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36071.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36071.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36071.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36071.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36071.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@36108.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@36108.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@36108.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@36108.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@36108.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@36140.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@36140.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@36140.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@36140.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@36140.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@36177.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@36177.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@36177.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@36177.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@36177.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@36191.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@36191.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@36191.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@36191.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@36191.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@36209.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@36209.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@36209.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@36209.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@36209.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@36266.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@36266.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@36266.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@36266.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@36266.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@36283.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@36283.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@36283.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@36283.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@36283.4]
  wire  _T_77; // @[Controllers.scala 80:47:@35944.4]
  wire  allDone; // @[Controllers.scala 80:47:@35945.4]
  wire  _T_151; // @[Controllers.scala 165:35:@36023.4]
  wire  _T_153; // @[Controllers.scala 165:60:@36024.4]
  wire  _T_154; // @[Controllers.scala 165:58:@36025.4]
  wire  _T_156; // @[Controllers.scala 165:76:@36026.4]
  wire  _T_157; // @[Controllers.scala 165:74:@36027.4]
  wire  _T_161; // @[Controllers.scala 165:109:@36030.4]
  wire  _T_164; // @[Controllers.scala 165:141:@36032.4]
  wire  _T_172; // @[package.scala 96:25:@36044.4 package.scala 96:25:@36045.4]
  wire  _T_176; // @[Controllers.scala 167:54:@36047.4]
  wire  _T_177; // @[Controllers.scala 167:52:@36048.4]
  wire  _T_184; // @[package.scala 96:25:@36058.4 package.scala 96:25:@36059.4]
  wire  _T_202; // @[package.scala 96:25:@36076.4 package.scala 96:25:@36077.4]
  wire  _T_206; // @[Controllers.scala 169:67:@36079.4]
  wire  _T_207; // @[Controllers.scala 169:86:@36080.4]
  wire  _T_219; // @[Controllers.scala 165:35:@36092.4]
  wire  _T_221; // @[Controllers.scala 165:60:@36093.4]
  wire  _T_222; // @[Controllers.scala 165:58:@36094.4]
  wire  _T_224; // @[Controllers.scala 165:76:@36095.4]
  wire  _T_225; // @[Controllers.scala 165:74:@36096.4]
  wire  _T_229; // @[Controllers.scala 165:109:@36099.4]
  wire  _T_232; // @[Controllers.scala 165:141:@36101.4]
  wire  _T_240; // @[package.scala 96:25:@36113.4 package.scala 96:25:@36114.4]
  wire  _T_244; // @[Controllers.scala 167:54:@36116.4]
  wire  _T_245; // @[Controllers.scala 167:52:@36117.4]
  wire  _T_252; // @[package.scala 96:25:@36127.4 package.scala 96:25:@36128.4]
  wire  _T_270; // @[package.scala 96:25:@36145.4 package.scala 96:25:@36146.4]
  wire  _T_274; // @[Controllers.scala 169:67:@36148.4]
  wire  _T_275; // @[Controllers.scala 169:86:@36149.4]
  wire  _T_287; // @[Controllers.scala 165:35:@36161.4]
  wire  _T_289; // @[Controllers.scala 165:60:@36162.4]
  wire  _T_290; // @[Controllers.scala 165:58:@36163.4]
  wire  _T_292; // @[Controllers.scala 165:76:@36164.4]
  wire  _T_293; // @[Controllers.scala 165:74:@36165.4]
  wire  _T_297; // @[Controllers.scala 165:109:@36168.4]
  wire  _T_300; // @[Controllers.scala 165:141:@36170.4]
  wire  _T_308; // @[package.scala 96:25:@36182.4 package.scala 96:25:@36183.4]
  wire  _T_312; // @[Controllers.scala 167:54:@36185.4]
  wire  _T_313; // @[Controllers.scala 167:52:@36186.4]
  wire  _T_320; // @[package.scala 96:25:@36196.4 package.scala 96:25:@36197.4]
  wire  _T_338; // @[package.scala 96:25:@36214.4 package.scala 96:25:@36215.4]
  wire  _T_342; // @[Controllers.scala 169:67:@36217.4]
  wire  _T_343; // @[Controllers.scala 169:86:@36218.4]
  wire  _T_358; // @[Controllers.scala 213:68:@36236.4]
  wire  _T_360; // @[Controllers.scala 213:90:@36238.4]
  wire  _T_362; // @[Controllers.scala 213:132:@36240.4]
  wire  _T_366; // @[Controllers.scala 213:68:@36245.4]
  wire  _T_368; // @[Controllers.scala 213:90:@36247.4]
  wire  _T_374; // @[Controllers.scala 213:68:@36253.4]
  wire  _T_376; // @[Controllers.scala 213:90:@36255.4]
  wire  _T_383; // @[package.scala 100:49:@36261.4]
  reg  _T_386; // @[package.scala 48:56:@36262.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@36264.4]
  reg  _T_400; // @[package.scala 48:56:@36280.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@35926.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@35929.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@35932.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@35935.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@35938.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@35941.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@35982.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@35985.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@35988.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36039.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36053.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36071.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@36108.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@36122.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@36140.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@36177.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@36191.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@36209.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@36266.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@36283.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@35944.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@35945.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@36023.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@36024.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@36025.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@36026.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@36027.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@36030.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@36032.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@36044.4 package.scala 96:25:@36045.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@36047.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@36048.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36058.4 package.scala 96:25:@36059.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36076.4 package.scala 96:25:@36077.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@36079.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@36080.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@36092.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@36093.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@36094.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@36095.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@36096.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@36099.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@36101.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@36113.4 package.scala 96:25:@36114.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@36116.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@36117.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@36127.4 package.scala 96:25:@36128.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@36145.4 package.scala 96:25:@36146.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@36148.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@36149.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@36161.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@36162.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@36163.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@36164.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@36165.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@36168.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@36170.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@36182.4 package.scala 96:25:@36183.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@36185.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@36186.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@36196.4 package.scala 96:25:@36197.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@36214.4 package.scala 96:25:@36215.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@36217.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@36218.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@36236.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@36238.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@36240.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@36245.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@36247.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@36253.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@36255.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@36261.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@36264.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@36290.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@36244.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@36252.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@36260.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@36231.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@36233.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@36235.4]
  assign active_0_clock = clock; // @[:@35927.4]
  assign active_0_reset = reset; // @[:@35928.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@36034.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@36038.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@35948.4]
  assign active_1_clock = clock; // @[:@35930.4]
  assign active_1_reset = reset; // @[:@35931.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@36103.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@36107.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@35949.4]
  assign active_2_clock = clock; // @[:@35933.4]
  assign active_2_reset = reset; // @[:@35934.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@36172.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@36176.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@35950.4]
  assign done_0_clock = clock; // @[:@35936.4]
  assign done_0_reset = reset; // @[:@35937.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@36084.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@35962.4 Controllers.scala 170:32:@36091.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@35951.4]
  assign done_1_clock = clock; // @[:@35939.4]
  assign done_1_reset = reset; // @[:@35940.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@36153.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@35971.4 Controllers.scala 170:32:@36160.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@35952.4]
  assign done_2_clock = clock; // @[:@35942.4]
  assign done_2_reset = reset; // @[:@35943.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@36222.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@35980.4 Controllers.scala 170:32:@36229.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@35953.4]
  assign iterDone_0_clock = clock; // @[:@35983.4]
  assign iterDone_0_reset = reset; // @[:@35984.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@36052.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@36002.4 Controllers.scala 168:36:@36068.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@35991.4]
  assign iterDone_1_clock = clock; // @[:@35986.4]
  assign iterDone_1_reset = reset; // @[:@35987.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@36121.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@36011.4 Controllers.scala 168:36:@36137.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@35992.4]
  assign iterDone_2_clock = clock; // @[:@35989.4]
  assign iterDone_2_reset = reset; // @[:@35990.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@36190.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@36020.4 Controllers.scala 168:36:@36206.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@35993.4]
  assign RetimeWrapper_clock = clock; // @[:@36040.4]
  assign RetimeWrapper_reset = reset; // @[:@36041.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36043.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@36042.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36054.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36055.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36057.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@36056.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36072.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36073.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36075.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@36074.4]
  assign RetimeWrapper_3_clock = clock; // @[:@36109.4]
  assign RetimeWrapper_3_reset = reset; // @[:@36110.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@36112.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@36111.4]
  assign RetimeWrapper_4_clock = clock; // @[:@36123.4]
  assign RetimeWrapper_4_reset = reset; // @[:@36124.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@36126.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@36125.4]
  assign RetimeWrapper_5_clock = clock; // @[:@36141.4]
  assign RetimeWrapper_5_reset = reset; // @[:@36142.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@36144.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@36143.4]
  assign RetimeWrapper_6_clock = clock; // @[:@36178.4]
  assign RetimeWrapper_6_reset = reset; // @[:@36179.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@36181.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@36180.4]
  assign RetimeWrapper_7_clock = clock; // @[:@36192.4]
  assign RetimeWrapper_7_reset = reset; // @[:@36193.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@36195.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@36194.4]
  assign RetimeWrapper_8_clock = clock; // @[:@36210.4]
  assign RetimeWrapper_8_reset = reset; // @[:@36211.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@36213.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@36212.4]
  assign RetimeWrapper_9_clock = clock; // @[:@36267.4]
  assign RetimeWrapper_9_reset = reset; // @[:@36268.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@36270.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@36269.4]
  assign RetimeWrapper_10_clock = clock; // @[:@36284.4]
  assign RetimeWrapper_10_reset = reset; // @[:@36285.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@36287.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@36286.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x479_inr_UnitPipe_sm( // @[:@36463.2]
  input   clock, // @[:@36464.4]
  input   reset, // @[:@36465.4]
  input   io_enable, // @[:@36466.4]
  output  io_done, // @[:@36466.4]
  output  io_doneLatch, // @[:@36466.4]
  input   io_ctrDone, // @[:@36466.4]
  output  io_datapathEn, // @[:@36466.4]
  output  io_ctrInc, // @[:@36466.4]
  input   io_parentAck, // @[:@36466.4]
  input   io_backpressure // @[:@36466.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@36468.4]
  wire  active_reset; // @[Controllers.scala 261:22:@36468.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@36468.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@36468.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@36468.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@36468.4]
  wire  done_clock; // @[Controllers.scala 262:20:@36471.4]
  wire  done_reset; // @[Controllers.scala 262:20:@36471.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@36471.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@36471.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@36471.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@36471.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36525.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36525.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36525.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36525.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36525.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36533.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36533.4]
  wire  _T_80; // @[Controllers.scala 264:48:@36476.4]
  wire  _T_81; // @[Controllers.scala 264:46:@36477.4]
  wire  _T_82; // @[Controllers.scala 264:62:@36478.4]
  wire  _T_83; // @[Controllers.scala 264:60:@36479.4]
  wire  _T_100; // @[package.scala 100:49:@36496.4]
  reg  _T_103; // @[package.scala 48:56:@36497.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@36505.4]
  wire  _T_116; // @[Controllers.scala 283:41:@36513.4]
  wire  _T_117; // @[Controllers.scala 283:59:@36514.4]
  wire  _T_119; // @[Controllers.scala 284:37:@36517.4]
  reg  _T_125; // @[package.scala 48:56:@36521.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@36543.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@36546.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@36548.4]
  wire  _T_152; // @[Controllers.scala 292:61:@36549.4]
  wire  _T_153; // @[Controllers.scala 292:24:@36550.4]
  SRFF active ( // @[Controllers.scala 261:22:@36468.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@36471.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36525.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36533.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@36476.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@36477.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@36478.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@36479.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@36496.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@36505.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@36513.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@36514.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@36517.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@36548.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@36549.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@36550.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@36524.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@36552.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@36516.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@36519.4]
  assign active_clock = clock; // @[:@36469.4]
  assign active_reset = reset; // @[:@36470.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@36481.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@36485.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@36486.4]
  assign done_clock = clock; // @[:@36472.4]
  assign done_reset = reset; // @[:@36473.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@36501.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@36494.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@36495.4]
  assign RetimeWrapper_clock = clock; // @[:@36526.4]
  assign RetimeWrapper_reset = reset; // @[:@36527.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36529.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@36528.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36534.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36535.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36537.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@36536.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1( // @[:@36627.2]
  output        io_in_x472_valid, // @[:@36630.4]
  output [63:0] io_in_x472_bits_addr, // @[:@36630.4]
  output [31:0] io_in_x472_bits_size, // @[:@36630.4]
  input  [63:0] io_in_x264_outdram_number, // @[:@36630.4]
  input         io_sigsIn_backpressure, // @[:@36630.4]
  input         io_sigsIn_datapathEn, // @[:@36630.4]
  input         io_rr // @[:@36630.4]
);
  wire [96:0] x476_tuple; // @[Cat.scala 30:58:@36644.4]
  wire  _T_135; // @[implicits.scala 55:10:@36647.4]
  assign x476_tuple = {33'h7e9000,io_in_x264_outdram_number}; // @[Cat.scala 30:58:@36644.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@36647.4]
  assign io_in_x472_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x479_inr_UnitPipe.scala 65:18:@36650.4]
  assign io_in_x472_bits_addr = x476_tuple[63:0]; // @[sm_x479_inr_UnitPipe.scala 66:22:@36652.4]
  assign io_in_x472_bits_size = x476_tuple[95:64]; // @[sm_x479_inr_UnitPipe.scala 67:22:@36654.4]
endmodule
module FF_13( // @[:@36656.2]
  input         clock, // @[:@36657.4]
  input         reset, // @[:@36658.4]
  output [22:0] io_rPort_0_output_0, // @[:@36659.4]
  input  [22:0] io_wPort_0_data_0, // @[:@36659.4]
  input         io_wPort_0_reset, // @[:@36659.4]
  input         io_wPort_0_en_0 // @[:@36659.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@36674.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@36676.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@36677.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@36676.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@36677.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@36679.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@36694.2]
  input         clock, // @[:@36695.4]
  input         reset, // @[:@36696.4]
  input         io_input_reset, // @[:@36697.4]
  input         io_input_enable, // @[:@36697.4]
  output [22:0] io_output_count_0, // @[:@36697.4]
  output        io_output_oobs_0, // @[:@36697.4]
  output        io_output_done // @[:@36697.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@36710.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@36710.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@36710.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@36710.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@36710.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@36710.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@36726.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@36726.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@36726.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@36726.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@36726.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@36726.4]
  wire  _T_36; // @[Counter.scala 264:45:@36729.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@36754.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@36755.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@36756.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@36757.4]
  wire  _T_57; // @[Counter.scala 293:18:@36759.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@36767.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@36770.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@36771.4]
  wire  _T_75; // @[Counter.scala 322:102:@36775.4]
  wire  _T_77; // @[Counter.scala 322:130:@36776.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@36710.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@36726.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@36729.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@36754.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@36755.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@36756.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@36757.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@36759.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@36767.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@36770.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@36771.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@36775.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@36776.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@36774.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@36778.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@36780.4]
  assign bases_0_clock = clock; // @[:@36711.4]
  assign bases_0_reset = reset; // @[:@36712.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@36773.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@36752.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@36753.4]
  assign SRFF_clock = clock; // @[:@36727.4]
  assign SRFF_reset = reset; // @[:@36728.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@36731.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@36733.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@36734.4]
endmodule
module x481_ctrchain( // @[:@36785.2]
  input         clock, // @[:@36786.4]
  input         reset, // @[:@36787.4]
  input         io_input_reset, // @[:@36788.4]
  input         io_input_enable, // @[:@36788.4]
  output [22:0] io_output_counts_0, // @[:@36788.4]
  output        io_output_oobs_0, // @[:@36788.4]
  output        io_output_done // @[:@36788.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@36790.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@36790.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@36790.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@36790.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@36790.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@36790.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@36790.4]
  reg  wasDone; // @[Counter.scala 542:24:@36799.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@36805.4]
  wire  _T_47; // @[Counter.scala 546:80:@36806.4]
  reg  doneLatch; // @[Counter.scala 550:26:@36811.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@36812.4]
  wire  _T_55; // @[Counter.scala 551:19:@36813.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@36790.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@36805.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@36806.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@36812.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@36813.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@36815.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@36817.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@36808.4]
  assign ctrs_0_clock = clock; // @[:@36791.4]
  assign ctrs_0_reset = reset; // @[:@36792.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@36796.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@36797.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x488_inr_Foreach_sm( // @[:@37005.2]
  input   clock, // @[:@37006.4]
  input   reset, // @[:@37007.4]
  input   io_enable, // @[:@37008.4]
  output  io_done, // @[:@37008.4]
  output  io_doneLatch, // @[:@37008.4]
  input   io_ctrDone, // @[:@37008.4]
  output  io_datapathEn, // @[:@37008.4]
  output  io_ctrInc, // @[:@37008.4]
  output  io_ctrRst, // @[:@37008.4]
  input   io_parentAck, // @[:@37008.4]
  input   io_backpressure, // @[:@37008.4]
  input   io_break // @[:@37008.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@37010.4]
  wire  active_reset; // @[Controllers.scala 261:22:@37010.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@37010.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@37010.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@37010.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@37010.4]
  wire  done_clock; // @[Controllers.scala 262:20:@37013.4]
  wire  done_reset; // @[Controllers.scala 262:20:@37013.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@37013.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@37013.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@37013.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@37013.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37047.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37047.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37047.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37047.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37047.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37069.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37069.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37069.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37069.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37069.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@37089.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@37089.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@37089.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@37089.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@37089.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@37105.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@37105.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@37105.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@37105.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@37105.4]
  wire  _T_80; // @[Controllers.scala 264:48:@37018.4]
  wire  _T_81; // @[Controllers.scala 264:46:@37019.4]
  wire  _T_82; // @[Controllers.scala 264:62:@37020.4]
  wire  _T_83; // @[Controllers.scala 264:60:@37021.4]
  wire  _T_100; // @[package.scala 100:49:@37038.4]
  reg  _T_103; // @[package.scala 48:56:@37039.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@37052.4 package.scala 96:25:@37053.4]
  wire  _T_110; // @[package.scala 100:49:@37054.4]
  reg  _T_113; // @[package.scala 48:56:@37055.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@37057.4]
  wire  _T_118; // @[Controllers.scala 283:41:@37062.4]
  wire  _T_119; // @[Controllers.scala 283:59:@37063.4]
  wire  _T_121; // @[Controllers.scala 284:37:@37066.4]
  wire  _T_124; // @[package.scala 96:25:@37074.4 package.scala 96:25:@37075.4]
  wire  _T_126; // @[package.scala 100:49:@37076.4]
  reg  _T_129; // @[package.scala 48:56:@37077.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@37099.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@37101.4]
  reg  _T_153; // @[package.scala 48:56:@37102.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@37110.4 package.scala 96:25:@37111.4]
  wire  _T_158; // @[Controllers.scala 292:61:@37112.4]
  wire  _T_159; // @[Controllers.scala 292:24:@37113.4]
  SRFF active ( // @[Controllers.scala 261:22:@37010.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@37013.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@37047.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@37069.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@37081.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@37089.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@37105.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@37018.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@37019.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@37020.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@37021.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@37038.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@37052.4 package.scala 96:25:@37053.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@37054.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@37057.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@37062.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@37063.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@37066.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37074.4 package.scala 96:25:@37075.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@37076.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@37101.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@37110.4 package.scala 96:25:@37111.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@37112.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@37113.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@37080.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@37115.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@37065.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@37068.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@37060.4]
  assign active_clock = clock; // @[:@37011.4]
  assign active_reset = reset; // @[:@37012.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@37023.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@37027.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@37028.4]
  assign done_clock = clock; // @[:@37014.4]
  assign done_reset = reset; // @[:@37015.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@37043.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@37036.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@37037.4]
  assign RetimeWrapper_clock = clock; // @[:@37048.4]
  assign RetimeWrapper_reset = reset; // @[:@37049.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@37051.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@37050.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37070.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37071.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@37073.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@37072.4]
  assign RetimeWrapper_2_clock = clock; // @[:@37082.4]
  assign RetimeWrapper_2_reset = reset; // @[:@37083.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@37085.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@37084.4]
  assign RetimeWrapper_3_clock = clock; // @[:@37090.4]
  assign RetimeWrapper_3_reset = reset; // @[:@37091.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@37093.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@37092.4]
  assign RetimeWrapper_4_clock = clock; // @[:@37106.4]
  assign RetimeWrapper_4_reset = reset; // @[:@37107.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@37109.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@37108.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x488_inr_Foreach_kernelx488_inr_Foreach_concrete1( // @[:@37322.2]
  input         clock, // @[:@37323.4]
  input         reset, // @[:@37324.4]
  output        io_in_x473_valid, // @[:@37325.4]
  output [31:0] io_in_x473_bits_wdata_0, // @[:@37325.4]
  output        io_in_x473_bits_wstrb, // @[:@37325.4]
  output [20:0] io_in_x268_outbuf_0_rPort_0_ofs_0, // @[:@37325.4]
  output        io_in_x268_outbuf_0_rPort_0_en_0, // @[:@37325.4]
  output        io_in_x268_outbuf_0_rPort_0_backpressure, // @[:@37325.4]
  input  [31:0] io_in_x268_outbuf_0_rPort_0_output_0, // @[:@37325.4]
  input         io_sigsIn_backpressure, // @[:@37325.4]
  input         io_sigsIn_datapathEn, // @[:@37325.4]
  input         io_sigsIn_break, // @[:@37325.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@37325.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@37325.4]
  input         io_rr // @[:@37325.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@37352.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@37352.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37381.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37381.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37381.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37381.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37381.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37390.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37390.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37390.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37390.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37390.4]
  wire  b483; // @[sm_x488_inr_Foreach.scala 62:18:@37360.4]
  wire  _T_274; // @[sm_x488_inr_Foreach.scala 67:129:@37364.4]
  wire  _T_278; // @[implicits.scala 55:10:@37367.4]
  wire  _T_279; // @[sm_x488_inr_Foreach.scala 67:146:@37368.4]
  wire [32:0] x486_tuple; // @[Cat.scala 30:58:@37378.4]
  wire  _T_290; // @[package.scala 96:25:@37395.4 package.scala 96:25:@37396.4]
  wire  _T_292; // @[implicits.scala 55:10:@37397.4]
  wire  x631_b483_D2; // @[package.scala 96:25:@37386.4 package.scala 96:25:@37387.4]
  wire  _T_293; // @[sm_x488_inr_Foreach.scala 74:112:@37398.4]
  wire [31:0] b482_number; // @[Math.scala 723:22:@37357.4 Math.scala 724:14:@37358.4]
  _ _ ( // @[Math.scala 720:24:@37352.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@37381.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@37390.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b483 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x488_inr_Foreach.scala 62:18:@37360.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x488_inr_Foreach.scala 67:129:@37364.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@37367.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x488_inr_Foreach.scala 67:146:@37368.4]
  assign x486_tuple = {1'h1,io_in_x268_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@37378.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37395.4 package.scala 96:25:@37396.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@37397.4]
  assign x631_b483_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@37386.4 package.scala 96:25:@37387.4]
  assign _T_293 = _T_292 & x631_b483_D2; // @[sm_x488_inr_Foreach.scala 74:112:@37398.4]
  assign b482_number = __io_result; // @[Math.scala 723:22:@37357.4 Math.scala 724:14:@37358.4]
  assign io_in_x473_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x488_inr_Foreach.scala 74:18:@37400.4]
  assign io_in_x473_bits_wdata_0 = x486_tuple[31:0]; // @[sm_x488_inr_Foreach.scala 75:26:@37402.4]
  assign io_in_x473_bits_wstrb = x486_tuple[32]; // @[sm_x488_inr_Foreach.scala 76:23:@37404.4]
  assign io_in_x268_outbuf_0_rPort_0_ofs_0 = b482_number[20:0]; // @[MemInterfaceType.scala 107:54:@37371.4]
  assign io_in_x268_outbuf_0_rPort_0_en_0 = _T_279 & b483; // @[MemInterfaceType.scala 110:79:@37373.4]
  assign io_in_x268_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@37372.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@37355.4]
  assign RetimeWrapper_clock = clock; // @[:@37382.4]
  assign RetimeWrapper_reset = reset; // @[:@37383.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37385.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@37384.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37391.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37392.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37394.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37393.4]
endmodule
module x492_inr_UnitPipe_sm( // @[:@37560.2]
  input   clock, // @[:@37561.4]
  input   reset, // @[:@37562.4]
  input   io_enable, // @[:@37563.4]
  output  io_done, // @[:@37563.4]
  output  io_doneLatch, // @[:@37563.4]
  input   io_ctrDone, // @[:@37563.4]
  output  io_datapathEn, // @[:@37563.4]
  output  io_ctrInc, // @[:@37563.4]
  input   io_parentAck // @[:@37563.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@37565.4]
  wire  active_reset; // @[Controllers.scala 261:22:@37565.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@37565.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@37565.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@37565.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@37565.4]
  wire  done_clock; // @[Controllers.scala 262:20:@37568.4]
  wire  done_reset; // @[Controllers.scala 262:20:@37568.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@37568.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@37568.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@37568.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@37568.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37602.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37602.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37602.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37602.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37602.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37624.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37624.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37624.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37624.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37624.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@37636.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@37636.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@37636.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@37636.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@37636.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@37644.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@37644.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@37644.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@37644.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@37644.4]
  wire  _T_80; // @[Controllers.scala 264:48:@37573.4]
  wire  _T_81; // @[Controllers.scala 264:46:@37574.4]
  wire  _T_82; // @[Controllers.scala 264:62:@37575.4]
  wire  _T_100; // @[package.scala 100:49:@37593.4]
  reg  _T_103; // @[package.scala 48:56:@37594.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@37617.4]
  wire  _T_124; // @[package.scala 96:25:@37629.4 package.scala 96:25:@37630.4]
  wire  _T_126; // @[package.scala 100:49:@37631.4]
  reg  _T_129; // @[package.scala 48:56:@37632.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@37654.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@37656.4]
  reg  _T_153; // @[package.scala 48:56:@37657.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@37659.4]
  wire  _T_156; // @[Controllers.scala 292:61:@37660.4]
  wire  _T_157; // @[Controllers.scala 292:24:@37661.4]
  SRFF active ( // @[Controllers.scala 261:22:@37565.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@37568.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@37602.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@37624.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@37636.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@37644.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@37573.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@37574.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@37575.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@37593.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@37617.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37629.4 package.scala 96:25:@37630.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@37631.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@37656.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@37659.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@37660.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@37661.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@37635.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@37663.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@37620.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@37623.4]
  assign active_clock = clock; // @[:@37566.4]
  assign active_reset = reset; // @[:@37567.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@37578.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@37582.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@37583.4]
  assign done_clock = clock; // @[:@37569.4]
  assign done_reset = reset; // @[:@37570.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@37598.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@37591.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@37592.4]
  assign RetimeWrapper_clock = clock; // @[:@37603.4]
  assign RetimeWrapper_reset = reset; // @[:@37604.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@37606.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@37605.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37625.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37626.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@37628.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@37627.4]
  assign RetimeWrapper_2_clock = clock; // @[:@37637.4]
  assign RetimeWrapper_2_reset = reset; // @[:@37638.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@37640.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@37639.4]
  assign RetimeWrapper_3_clock = clock; // @[:@37645.4]
  assign RetimeWrapper_3_reset = reset; // @[:@37646.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@37648.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@37647.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1( // @[:@37738.2]
  output  io_in_x474_ready, // @[:@37741.4]
  input   io_sigsIn_datapathEn // @[:@37741.4]
);
  assign io_in_x474_ready = io_sigsIn_datapathEn; // @[sm_x492_inr_UnitPipe.scala 57:18:@37753.4]
endmodule
module x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1( // @[:@37756.2]
  input         clock, // @[:@37757.4]
  input         reset, // @[:@37758.4]
  input         io_in_x472_ready, // @[:@37759.4]
  output        io_in_x472_valid, // @[:@37759.4]
  output [63:0] io_in_x472_bits_addr, // @[:@37759.4]
  output [31:0] io_in_x472_bits_size, // @[:@37759.4]
  input  [63:0] io_in_x264_outdram_number, // @[:@37759.4]
  input         io_in_x473_ready, // @[:@37759.4]
  output        io_in_x473_valid, // @[:@37759.4]
  output [31:0] io_in_x473_bits_wdata_0, // @[:@37759.4]
  output        io_in_x473_bits_wstrb, // @[:@37759.4]
  output [20:0] io_in_x268_outbuf_0_rPort_0_ofs_0, // @[:@37759.4]
  output        io_in_x268_outbuf_0_rPort_0_en_0, // @[:@37759.4]
  output        io_in_x268_outbuf_0_rPort_0_backpressure, // @[:@37759.4]
  input  [31:0] io_in_x268_outbuf_0_rPort_0_output_0, // @[:@37759.4]
  output        io_in_x474_ready, // @[:@37759.4]
  input         io_in_x474_valid, // @[:@37759.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@37759.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@37759.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@37759.4]
  input         io_sigsIn_smChildAcks_0, // @[:@37759.4]
  input         io_sigsIn_smChildAcks_1, // @[:@37759.4]
  input         io_sigsIn_smChildAcks_2, // @[:@37759.4]
  output        io_sigsOut_smDoneIn_0, // @[:@37759.4]
  output        io_sigsOut_smDoneIn_1, // @[:@37759.4]
  output        io_sigsOut_smDoneIn_2, // @[:@37759.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@37759.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@37759.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@37759.4]
  input         io_rr // @[:@37759.4]
);
  wire  x479_inr_UnitPipe_sm_clock; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_reset; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_enable; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_done; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_doneLatch; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_ctrDone; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_datapathEn; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_ctrInc; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_parentAck; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  x479_inr_UnitPipe_sm_io_backpressure; // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37883.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37883.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37883.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37883.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37883.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37891.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37891.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37891.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37891.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37891.4]
  wire  x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_valid; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire [63:0] x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_bits_addr; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire [31:0] x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_bits_size; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire [63:0] x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x264_outdram_number; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire  x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire  x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire  x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_rr; // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
  wire  x481_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire  x481_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire  x481_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire  x481_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire [22:0] x481_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire  x481_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire  x481_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@37989.4]
  wire  x488_inr_Foreach_sm_clock; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_reset; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_enable; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_done; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_doneLatch; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_ctrDone; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_datapathEn; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_ctrInc; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_ctrRst; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_parentAck; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_backpressure; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  x488_inr_Foreach_sm_io_break; // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38070.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38070.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38070.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38070.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38070.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38110.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38110.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38110.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38110.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38110.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@38118.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@38118.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@38118.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@38118.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@38118.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_clock; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_reset; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_valid; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire [31:0] x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_bits_wdata_0; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_bits_wstrb; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire [20:0] x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_en_0; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire [31:0] x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_output_0; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire [31:0] x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_rr; // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
  wire  x492_inr_UnitPipe_sm_clock; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_reset; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_enable; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_done; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_doneLatch; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_ctrDone; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_datapathEn; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_ctrInc; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  x492_inr_UnitPipe_sm_io_parentAck; // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@38330.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@38330.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@38330.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@38330.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@38330.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@38338.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@38338.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@38338.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@38338.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@38338.4]
  wire  x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1_io_in_x474_ready; // @[sm_x492_inr_UnitPipe.scala 60:24:@38368.4]
  wire  x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x492_inr_UnitPipe.scala 60:24:@38368.4]
  wire  _T_359; // @[package.scala 100:49:@37854.4]
  reg  _T_362; // @[package.scala 48:56:@37855.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@37888.4 package.scala 96:25:@37889.4]
  wire  _T_381; // @[package.scala 96:25:@37896.4 package.scala 96:25:@37897.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@37899.4]
  wire  _T_454; // @[package.scala 96:25:@38075.4 package.scala 96:25:@38076.4]
  wire  _T_468; // @[package.scala 96:25:@38115.4 package.scala 96:25:@38116.4]
  wire  _T_474; // @[package.scala 96:25:@38123.4 package.scala 96:25:@38124.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@38126.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@38135.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@38136.4]
  wire  _T_547; // @[package.scala 100:49:@38301.4]
  reg  _T_550; // @[package.scala 48:56:@38302.4]
  reg [31:0] _RAND_1;
  wire  x492_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x493_outr_UnitPipe.scala 101:55:@38308.4]
  wire  _T_563; // @[package.scala 96:25:@38335.4 package.scala 96:25:@38336.4]
  wire  _T_569; // @[package.scala 96:25:@38343.4 package.scala 96:25:@38344.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@38346.4]
  wire  x492_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@38347.4]
  x479_inr_UnitPipe_sm x479_inr_UnitPipe_sm ( // @[sm_x479_inr_UnitPipe.scala 33:18:@37826.4]
    .clock(x479_inr_UnitPipe_sm_clock),
    .reset(x479_inr_UnitPipe_sm_reset),
    .io_enable(x479_inr_UnitPipe_sm_io_enable),
    .io_done(x479_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x479_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x479_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x479_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x479_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x479_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x479_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@37883.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@37891.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1 x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1 ( // @[sm_x479_inr_UnitPipe.scala 69:24:@37921.4]
    .io_in_x472_valid(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_valid),
    .io_in_x472_bits_addr(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_bits_addr),
    .io_in_x472_bits_size(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_bits_size),
    .io_in_x264_outdram_number(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x264_outdram_number),
    .io_sigsIn_backpressure(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_rr)
  );
  x481_ctrchain x481_ctrchain ( // @[SpatialBlocks.scala 37:22:@37989.4]
    .clock(x481_ctrchain_clock),
    .reset(x481_ctrchain_reset),
    .io_input_reset(x481_ctrchain_io_input_reset),
    .io_input_enable(x481_ctrchain_io_input_enable),
    .io_output_counts_0(x481_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x481_ctrchain_io_output_oobs_0),
    .io_output_done(x481_ctrchain_io_output_done)
  );
  x488_inr_Foreach_sm x488_inr_Foreach_sm ( // @[sm_x488_inr_Foreach.scala 33:18:@38042.4]
    .clock(x488_inr_Foreach_sm_clock),
    .reset(x488_inr_Foreach_sm_reset),
    .io_enable(x488_inr_Foreach_sm_io_enable),
    .io_done(x488_inr_Foreach_sm_io_done),
    .io_doneLatch(x488_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x488_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x488_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x488_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x488_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x488_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x488_inr_Foreach_sm_io_backpressure),
    .io_break(x488_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38070.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38110.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@38118.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x488_inr_Foreach_kernelx488_inr_Foreach_concrete1 x488_inr_Foreach_kernelx488_inr_Foreach_concrete1 ( // @[sm_x488_inr_Foreach.scala 78:24:@38153.4]
    .clock(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_clock),
    .reset(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_reset),
    .io_in_x473_valid(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_valid),
    .io_in_x473_bits_wdata_0(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_bits_wdata_0),
    .io_in_x473_bits_wstrb(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_bits_wstrb),
    .io_in_x268_outbuf_0_rPort_0_ofs_0(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0),
    .io_in_x268_outbuf_0_rPort_0_en_0(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_en_0),
    .io_in_x268_outbuf_0_rPort_0_backpressure(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure),
    .io_in_x268_outbuf_0_rPort_0_output_0(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_output_0),
    .io_sigsIn_backpressure(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_rr)
  );
  x492_inr_UnitPipe_sm x492_inr_UnitPipe_sm ( // @[sm_x492_inr_UnitPipe.scala 32:18:@38273.4]
    .clock(x492_inr_UnitPipe_sm_clock),
    .reset(x492_inr_UnitPipe_sm_reset),
    .io_enable(x492_inr_UnitPipe_sm_io_enable),
    .io_done(x492_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x492_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x492_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x492_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x492_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x492_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@38330.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@38338.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1 x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1 ( // @[sm_x492_inr_UnitPipe.scala 60:24:@38368.4]
    .io_in_x474_ready(x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1_io_in_x474_ready),
    .io_sigsIn_datapathEn(x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x479_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@37854.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@37888.4 package.scala 96:25:@37889.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37896.4 package.scala 96:25:@37897.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@37899.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@38075.4 package.scala 96:25:@38076.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@38115.4 package.scala 96:25:@38116.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@38123.4 package.scala 96:25:@38124.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@38126.4]
  assign _T_479 = x488_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@38135.4]
  assign _T_480 = ~ x488_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@38136.4]
  assign _T_547 = x492_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@38301.4]
  assign x492_inr_UnitPipe_sigsIn_forwardpressure = io_in_x474_valid | x492_inr_UnitPipe_sm_io_doneLatch; // @[sm_x493_outr_UnitPipe.scala 101:55:@38308.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@38335.4 package.scala 96:25:@38336.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@38343.4 package.scala 96:25:@38344.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@38346.4]
  assign x492_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@38347.4]
  assign io_in_x472_valid = x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_valid; // @[sm_x479_inr_UnitPipe.scala 49:23:@37959.4]
  assign io_in_x472_bits_addr = x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_bits_addr; // @[sm_x479_inr_UnitPipe.scala 49:23:@37958.4]
  assign io_in_x472_bits_size = x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x472_bits_size; // @[sm_x479_inr_UnitPipe.scala 49:23:@37957.4]
  assign io_in_x473_valid = x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_valid; // @[sm_x488_inr_Foreach.scala 49:23:@38203.4]
  assign io_in_x473_bits_wdata_0 = x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_bits_wdata_0; // @[sm_x488_inr_Foreach.scala 49:23:@38202.4]
  assign io_in_x473_bits_wstrb = x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x473_bits_wstrb; // @[sm_x488_inr_Foreach.scala 49:23:@38201.4]
  assign io_in_x268_outbuf_0_rPort_0_ofs_0 = x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@38208.4]
  assign io_in_x268_outbuf_0_rPort_0_en_0 = x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@38207.4]
  assign io_in_x268_outbuf_0_rPort_0_backpressure = x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@38206.4]
  assign io_in_x474_ready = x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1_io_in_x474_ready; // @[sm_x492_inr_UnitPipe.scala 46:23:@38404.4]
  assign io_sigsOut_smDoneIn_0 = x479_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@37906.4]
  assign io_sigsOut_smDoneIn_1 = x488_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@38133.4]
  assign io_sigsOut_smDoneIn_2 = x492_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@38353.4]
  assign io_sigsOut_smCtrCopyDone_0 = x479_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@37920.4]
  assign io_sigsOut_smCtrCopyDone_1 = x488_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@38152.4]
  assign io_sigsOut_smCtrCopyDone_2 = x492_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@38367.4]
  assign x479_inr_UnitPipe_sm_clock = clock; // @[:@37827.4]
  assign x479_inr_UnitPipe_sm_reset = reset; // @[:@37828.4]
  assign x479_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@37903.4]
  assign x479_inr_UnitPipe_sm_io_ctrDone = x479_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x493_outr_UnitPipe.scala 77:39:@37858.4]
  assign x479_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@37905.4]
  assign x479_inr_UnitPipe_sm_io_backpressure = io_in_x472_ready | x479_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@37877.4]
  assign RetimeWrapper_clock = clock; // @[:@37884.4]
  assign RetimeWrapper_reset = reset; // @[:@37885.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@37887.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@37886.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37892.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37893.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@37895.4]
  assign RetimeWrapper_1_io_in = x479_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@37894.4]
  assign x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_in_x264_outdram_number = io_in_x264_outdram_number; // @[sm_x479_inr_UnitPipe.scala 50:31:@37961.4]
  assign x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x472_ready | x479_inr_UnitPipe_sm_io_doneLatch; // @[sm_x479_inr_UnitPipe.scala 74:22:@37976.4]
  assign x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x479_inr_UnitPipe_sm_io_datapathEn; // @[sm_x479_inr_UnitPipe.scala 74:22:@37974.4]
  assign x479_inr_UnitPipe_kernelx479_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x479_inr_UnitPipe.scala 73:18:@37962.4]
  assign x481_ctrchain_clock = clock; // @[:@37990.4]
  assign x481_ctrchain_reset = reset; // @[:@37991.4]
  assign x481_ctrchain_io_input_reset = x488_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@38151.4]
  assign x481_ctrchain_io_input_enable = x488_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@38103.4 SpatialBlocks.scala 159:42:@38150.4]
  assign x488_inr_Foreach_sm_clock = clock; // @[:@38043.4]
  assign x488_inr_Foreach_sm_reset = reset; // @[:@38044.4]
  assign x488_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@38130.4]
  assign x488_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x493_outr_UnitPipe.scala 90:38:@38078.4]
  assign x488_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@38132.4]
  assign x488_inr_Foreach_sm_io_backpressure = io_in_x473_ready | x488_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@38104.4]
  assign x488_inr_Foreach_sm_io_break = 1'h0; // @[sm_x493_outr_UnitPipe.scala 94:36:@38084.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38071.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38072.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38074.4]
  assign RetimeWrapper_2_io_in = x481_ctrchain_io_output_done; // @[package.scala 94:16:@38073.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38111.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38112.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38114.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@38113.4]
  assign RetimeWrapper_4_clock = clock; // @[:@38119.4]
  assign RetimeWrapper_4_reset = reset; // @[:@38120.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@38122.4]
  assign RetimeWrapper_4_io_in = x488_inr_Foreach_sm_io_done; // @[package.scala 94:16:@38121.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_clock = clock; // @[:@38154.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_reset = reset; // @[:@38155.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_in_x268_outbuf_0_rPort_0_output_0 = io_in_x268_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@38205.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x473_ready | x488_inr_Foreach_sm_io_doneLatch; // @[sm_x488_inr_Foreach.scala 83:22:@38224.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x488_inr_Foreach.scala 83:22:@38222.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_break = x488_inr_Foreach_sm_io_break; // @[sm_x488_inr_Foreach.scala 83:22:@38220.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x481_ctrchain_io_output_counts_0[22]}},x481_ctrchain_io_output_counts_0}; // @[sm_x488_inr_Foreach.scala 83:22:@38215.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x481_ctrchain_io_output_oobs_0; // @[sm_x488_inr_Foreach.scala 83:22:@38214.4]
  assign x488_inr_Foreach_kernelx488_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x488_inr_Foreach.scala 82:18:@38210.4]
  assign x492_inr_UnitPipe_sm_clock = clock; // @[:@38274.4]
  assign x492_inr_UnitPipe_sm_reset = reset; // @[:@38275.4]
  assign x492_inr_UnitPipe_sm_io_enable = x492_inr_UnitPipe_sigsIn_baseEn & x492_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@38350.4]
  assign x492_inr_UnitPipe_sm_io_ctrDone = x492_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x493_outr_UnitPipe.scala 99:39:@38305.4]
  assign x492_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@38352.4]
  assign RetimeWrapper_5_clock = clock; // @[:@38331.4]
  assign RetimeWrapper_5_reset = reset; // @[:@38332.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@38334.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@38333.4]
  assign RetimeWrapper_6_clock = clock; // @[:@38339.4]
  assign RetimeWrapper_6_reset = reset; // @[:@38340.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@38342.4]
  assign RetimeWrapper_6_io_in = x492_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@38341.4]
  assign x492_inr_UnitPipe_kernelx492_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x492_inr_UnitPipe_sm_io_datapathEn; // @[sm_x492_inr_UnitPipe.scala 65:22:@38417.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x542_kernelx542_concrete1( // @[:@38433.2]
  input          clock, // @[:@38434.4]
  input          reset, // @[:@38435.4]
  input          io_in_x472_ready, // @[:@38436.4]
  output         io_in_x472_valid, // @[:@38436.4]
  output [63:0]  io_in_x472_bits_addr, // @[:@38436.4]
  output [31:0]  io_in_x472_bits_size, // @[:@38436.4]
  input          io_in_x266_TVALID, // @[:@38436.4]
  output         io_in_x266_TREADY, // @[:@38436.4]
  input  [255:0] io_in_x266_TDATA, // @[:@38436.4]
  input  [7:0]   io_in_x266_TID, // @[:@38436.4]
  input  [7:0]   io_in_x266_TDEST, // @[:@38436.4]
  input  [63:0]  io_in_x264_outdram_number, // @[:@38436.4]
  output         io_in_x267_TVALID, // @[:@38436.4]
  input          io_in_x267_TREADY, // @[:@38436.4]
  output [255:0] io_in_x267_TDATA, // @[:@38436.4]
  input          io_in_x473_ready, // @[:@38436.4]
  output         io_in_x473_valid, // @[:@38436.4]
  output [31:0]  io_in_x473_bits_wdata_0, // @[:@38436.4]
  output         io_in_x473_bits_wstrb, // @[:@38436.4]
  output [20:0]  io_in_x268_outbuf_0_rPort_0_ofs_0, // @[:@38436.4]
  output         io_in_x268_outbuf_0_rPort_0_en_0, // @[:@38436.4]
  output         io_in_x268_outbuf_0_rPort_0_backpressure, // @[:@38436.4]
  input  [31:0]  io_in_x268_outbuf_0_rPort_0_output_0, // @[:@38436.4]
  output         io_in_x474_ready, // @[:@38436.4]
  input          io_in_x474_valid, // @[:@38436.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@38436.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@38436.4]
  input          io_sigsIn_smChildAcks_0, // @[:@38436.4]
  input          io_sigsIn_smChildAcks_1, // @[:@38436.4]
  output         io_sigsOut_smDoneIn_0, // @[:@38436.4]
  output         io_sigsOut_smDoneIn_1, // @[:@38436.4]
  input          io_rr // @[:@38436.4]
);
  wire  x471_outr_UnitPipe_sm_clock; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_reset; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_enable; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_done; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_parentAck; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_childAck_0; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_childAck_1; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  x471_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38571.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38571.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38571.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38571.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38571.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38579.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38579.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38579.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38579.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38579.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_clock; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_reset; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TVALID; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TREADY; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire [255:0] x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TDATA; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire [7:0] x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TID; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire [7:0] x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TDEST; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TVALID; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TREADY; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire [255:0] x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TDATA; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_rr; // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
  wire  x493_outr_UnitPipe_sm_clock; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_reset; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_enable; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_done; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_parentAck; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_childAck_0; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_childAck_1; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_childAck_2; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  x493_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38860.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38868.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38868.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38868.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38868.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38868.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_clock; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_reset; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_ready; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_valid; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire [63:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_bits_addr; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire [31:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_bits_size; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire [63:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x264_outdram_number; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_ready; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_valid; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire [31:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_bits_wdata_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_bits_wstrb; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire [20:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_en_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire [31:0] x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_output_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x474_ready; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x474_valid; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_rr; // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
  wire  _T_408; // @[package.scala 96:25:@38576.4 package.scala 96:25:@38577.4]
  wire  _T_414; // @[package.scala 96:25:@38584.4 package.scala 96:25:@38585.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@38587.4]
  wire  _T_508; // @[package.scala 96:25:@38865.4 package.scala 96:25:@38866.4]
  wire  _T_514; // @[package.scala 96:25:@38873.4 package.scala 96:25:@38874.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@38876.4]
  x471_outr_UnitPipe_sm x471_outr_UnitPipe_sm ( // @[sm_x471_outr_UnitPipe.scala 32:18:@38509.4]
    .clock(x471_outr_UnitPipe_sm_clock),
    .reset(x471_outr_UnitPipe_sm_reset),
    .io_enable(x471_outr_UnitPipe_sm_io_enable),
    .io_done(x471_outr_UnitPipe_sm_io_done),
    .io_parentAck(x471_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x471_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x471_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x471_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x471_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x471_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x471_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x471_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x471_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@38571.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@38579.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1 x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1 ( // @[sm_x471_outr_UnitPipe.scala 87:24:@38610.4]
    .clock(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_clock),
    .reset(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_reset),
    .io_in_x266_TVALID(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TVALID),
    .io_in_x266_TREADY(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TREADY),
    .io_in_x266_TDATA(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TDATA),
    .io_in_x266_TID(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TID),
    .io_in_x266_TDEST(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TDEST),
    .io_in_x267_TVALID(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TVALID),
    .io_in_x267_TREADY(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TREADY),
    .io_in_x267_TDATA(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TDATA),
    .io_sigsIn_smEnableOuts_0(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_rr)
  );
  x493_outr_UnitPipe_sm x493_outr_UnitPipe_sm ( // @[sm_x493_outr_UnitPipe.scala 36:18:@38788.4]
    .clock(x493_outr_UnitPipe_sm_clock),
    .reset(x493_outr_UnitPipe_sm_reset),
    .io_enable(x493_outr_UnitPipe_sm_io_enable),
    .io_done(x493_outr_UnitPipe_sm_io_done),
    .io_parentAck(x493_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x493_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x493_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x493_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x493_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x493_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x493_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x493_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x493_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x493_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x493_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x493_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x493_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38860.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38868.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1 x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1 ( // @[sm_x493_outr_UnitPipe.scala 108:24:@38900.4]
    .clock(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_clock),
    .reset(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_reset),
    .io_in_x472_ready(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_ready),
    .io_in_x472_valid(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_valid),
    .io_in_x472_bits_addr(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_bits_addr),
    .io_in_x472_bits_size(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_bits_size),
    .io_in_x264_outdram_number(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x264_outdram_number),
    .io_in_x473_ready(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_ready),
    .io_in_x473_valid(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_valid),
    .io_in_x473_bits_wdata_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_bits_wdata_0),
    .io_in_x473_bits_wstrb(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_bits_wstrb),
    .io_in_x268_outbuf_0_rPort_0_ofs_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0),
    .io_in_x268_outbuf_0_rPort_0_en_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_en_0),
    .io_in_x268_outbuf_0_rPort_0_backpressure(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure),
    .io_in_x268_outbuf_0_rPort_0_output_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_output_0),
    .io_in_x474_ready(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x474_ready),
    .io_in_x474_valid(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x474_valid),
    .io_sigsIn_smEnableOuts_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@38576.4 package.scala 96:25:@38577.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38584.4 package.scala 96:25:@38585.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@38587.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@38865.4 package.scala 96:25:@38866.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@38873.4 package.scala 96:25:@38874.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@38876.4]
  assign io_in_x472_valid = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_valid; // @[sm_x493_outr_UnitPipe.scala 58:23:@38982.4]
  assign io_in_x472_bits_addr = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_bits_addr; // @[sm_x493_outr_UnitPipe.scala 58:23:@38981.4]
  assign io_in_x472_bits_size = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_bits_size; // @[sm_x493_outr_UnitPipe.scala 58:23:@38980.4]
  assign io_in_x266_TREADY = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TREADY; // @[sm_x471_outr_UnitPipe.scala 48:23:@38678.4]
  assign io_in_x267_TVALID = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TVALID; // @[sm_x471_outr_UnitPipe.scala 49:23:@38688.4]
  assign io_in_x267_TDATA = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TDATA; // @[sm_x471_outr_UnitPipe.scala 49:23:@38686.4]
  assign io_in_x473_valid = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_valid; // @[sm_x493_outr_UnitPipe.scala 60:23:@38987.4]
  assign io_in_x473_bits_wdata_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_bits_wdata_0; // @[sm_x493_outr_UnitPipe.scala 60:23:@38986.4]
  assign io_in_x473_bits_wstrb = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_bits_wstrb; // @[sm_x493_outr_UnitPipe.scala 60:23:@38985.4]
  assign io_in_x268_outbuf_0_rPort_0_ofs_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@38992.4]
  assign io_in_x268_outbuf_0_rPort_0_en_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@38991.4]
  assign io_in_x268_outbuf_0_rPort_0_backpressure = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@38990.4]
  assign io_in_x474_ready = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x474_ready; // @[sm_x493_outr_UnitPipe.scala 62:23:@38996.4]
  assign io_sigsOut_smDoneIn_0 = x471_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@38594.4]
  assign io_sigsOut_smDoneIn_1 = x493_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@38883.4]
  assign x471_outr_UnitPipe_sm_clock = clock; // @[:@38510.4]
  assign x471_outr_UnitPipe_sm_reset = reset; // @[:@38511.4]
  assign x471_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@38591.4]
  assign x471_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@38593.4]
  assign x471_outr_UnitPipe_sm_io_doneIn_0 = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@38561.4]
  assign x471_outr_UnitPipe_sm_io_doneIn_1 = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@38562.4]
  assign x471_outr_UnitPipe_sm_io_ctrCopyDone_0 = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@38608.4]
  assign x471_outr_UnitPipe_sm_io_ctrCopyDone_1 = x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@38609.4]
  assign RetimeWrapper_clock = clock; // @[:@38572.4]
  assign RetimeWrapper_reset = reset; // @[:@38573.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@38575.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@38574.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38580.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38581.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@38583.4]
  assign RetimeWrapper_1_io_in = x471_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@38582.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_clock = clock; // @[:@38611.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_reset = reset; // @[:@38612.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TVALID = io_in_x266_TVALID; // @[sm_x471_outr_UnitPipe.scala 48:23:@38679.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TDATA = io_in_x266_TDATA; // @[sm_x471_outr_UnitPipe.scala 48:23:@38677.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TID = io_in_x266_TID; // @[sm_x471_outr_UnitPipe.scala 48:23:@38673.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x266_TDEST = io_in_x266_TDEST; // @[sm_x471_outr_UnitPipe.scala 48:23:@38672.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_in_x267_TREADY = io_in_x267_TREADY; // @[sm_x471_outr_UnitPipe.scala 49:23:@38687.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x471_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x471_outr_UnitPipe.scala 92:22:@38704.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x471_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x471_outr_UnitPipe.scala 92:22:@38705.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x471_outr_UnitPipe_sm_io_childAck_0; // @[sm_x471_outr_UnitPipe.scala 92:22:@38700.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x471_outr_UnitPipe_sm_io_childAck_1; // @[sm_x471_outr_UnitPipe.scala 92:22:@38701.4]
  assign x471_outr_UnitPipe_kernelx471_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x471_outr_UnitPipe.scala 91:18:@38689.4]
  assign x493_outr_UnitPipe_sm_clock = clock; // @[:@38789.4]
  assign x493_outr_UnitPipe_sm_reset = reset; // @[:@38790.4]
  assign x493_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@38880.4]
  assign x493_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@38882.4]
  assign x493_outr_UnitPipe_sm_io_doneIn_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@38848.4]
  assign x493_outr_UnitPipe_sm_io_doneIn_1 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@38849.4]
  assign x493_outr_UnitPipe_sm_io_doneIn_2 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@38850.4]
  assign x493_outr_UnitPipe_sm_io_ctrCopyDone_0 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@38897.4]
  assign x493_outr_UnitPipe_sm_io_ctrCopyDone_1 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@38898.4]
  assign x493_outr_UnitPipe_sm_io_ctrCopyDone_2 = x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@38899.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38861.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38862.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38864.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@38863.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38869.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38870.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38872.4]
  assign RetimeWrapper_3_io_in = x493_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@38871.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_clock = clock; // @[:@38901.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_reset = reset; // @[:@38902.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x472_ready = io_in_x472_ready; // @[sm_x493_outr_UnitPipe.scala 58:23:@38983.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x264_outdram_number = io_in_x264_outdram_number; // @[sm_x493_outr_UnitPipe.scala 59:31:@38984.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x473_ready = io_in_x473_ready; // @[sm_x493_outr_UnitPipe.scala 60:23:@38988.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x268_outbuf_0_rPort_0_output_0 = io_in_x268_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@38989.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_in_x474_valid = io_in_x474_valid; // @[sm_x493_outr_UnitPipe.scala 62:23:@38995.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x493_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x493_outr_UnitPipe.scala 113:22:@39019.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x493_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x493_outr_UnitPipe.scala 113:22:@39020.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x493_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x493_outr_UnitPipe.scala 113:22:@39021.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x493_outr_UnitPipe_sm_io_childAck_0; // @[sm_x493_outr_UnitPipe.scala 113:22:@39013.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x493_outr_UnitPipe_sm_io_childAck_1; // @[sm_x493_outr_UnitPipe.scala 113:22:@39014.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x493_outr_UnitPipe_sm_io_childAck_2; // @[sm_x493_outr_UnitPipe.scala 113:22:@39015.4]
  assign x493_outr_UnitPipe_kernelx493_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x493_outr_UnitPipe.scala 112:18:@38997.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@39049.2]
  input          clock, // @[:@39050.4]
  input          reset, // @[:@39051.4]
  input          io_in_x472_ready, // @[:@39052.4]
  output         io_in_x472_valid, // @[:@39052.4]
  output [63:0]  io_in_x472_bits_addr, // @[:@39052.4]
  output [31:0]  io_in_x472_bits_size, // @[:@39052.4]
  input          io_in_x266_TVALID, // @[:@39052.4]
  output         io_in_x266_TREADY, // @[:@39052.4]
  input  [255:0] io_in_x266_TDATA, // @[:@39052.4]
  input  [7:0]   io_in_x266_TID, // @[:@39052.4]
  input  [7:0]   io_in_x266_TDEST, // @[:@39052.4]
  input  [63:0]  io_in_x264_outdram_number, // @[:@39052.4]
  output         io_in_x267_TVALID, // @[:@39052.4]
  input          io_in_x267_TREADY, // @[:@39052.4]
  output [255:0] io_in_x267_TDATA, // @[:@39052.4]
  input          io_in_x473_ready, // @[:@39052.4]
  output         io_in_x473_valid, // @[:@39052.4]
  output [31:0]  io_in_x473_bits_wdata_0, // @[:@39052.4]
  output         io_in_x473_bits_wstrb, // @[:@39052.4]
  output         io_in_x474_ready, // @[:@39052.4]
  input          io_in_x474_valid, // @[:@39052.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@39052.4]
  input          io_sigsIn_smChildAcks_0, // @[:@39052.4]
  output         io_sigsOut_smDoneIn_0, // @[:@39052.4]
  input          io_rr // @[:@39052.4]
);
  wire  x268_outbuf_0_clock; // @[m_x268_outbuf_0.scala 27:17:@39062.4]
  wire  x268_outbuf_0_reset; // @[m_x268_outbuf_0.scala 27:17:@39062.4]
  wire [20:0] x268_outbuf_0_io_rPort_0_ofs_0; // @[m_x268_outbuf_0.scala 27:17:@39062.4]
  wire  x268_outbuf_0_io_rPort_0_en_0; // @[m_x268_outbuf_0.scala 27:17:@39062.4]
  wire  x268_outbuf_0_io_rPort_0_backpressure; // @[m_x268_outbuf_0.scala 27:17:@39062.4]
  wire [31:0] x268_outbuf_0_io_rPort_0_output_0; // @[m_x268_outbuf_0.scala 27:17:@39062.4]
  wire  x542_sm_clock; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_reset; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_enable; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_done; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_ctrDone; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_ctrInc; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_parentAck; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_doneIn_0; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_doneIn_1; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_enableOut_0; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_enableOut_1; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_childAck_0; // @[sm_x542.scala 37:18:@39120.4]
  wire  x542_sm_io_childAck_1; // @[sm_x542.scala 37:18:@39120.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39195.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39195.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39195.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39195.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39195.4]
  wire  x542_kernelx542_concrete1_clock; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_reset; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x472_ready; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x472_valid; // @[sm_x542.scala 102:24:@39224.4]
  wire [63:0] x542_kernelx542_concrete1_io_in_x472_bits_addr; // @[sm_x542.scala 102:24:@39224.4]
  wire [31:0] x542_kernelx542_concrete1_io_in_x472_bits_size; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x266_TVALID; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x266_TREADY; // @[sm_x542.scala 102:24:@39224.4]
  wire [255:0] x542_kernelx542_concrete1_io_in_x266_TDATA; // @[sm_x542.scala 102:24:@39224.4]
  wire [7:0] x542_kernelx542_concrete1_io_in_x266_TID; // @[sm_x542.scala 102:24:@39224.4]
  wire [7:0] x542_kernelx542_concrete1_io_in_x266_TDEST; // @[sm_x542.scala 102:24:@39224.4]
  wire [63:0] x542_kernelx542_concrete1_io_in_x264_outdram_number; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x267_TVALID; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x267_TREADY; // @[sm_x542.scala 102:24:@39224.4]
  wire [255:0] x542_kernelx542_concrete1_io_in_x267_TDATA; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x473_ready; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x473_valid; // @[sm_x542.scala 102:24:@39224.4]
  wire [31:0] x542_kernelx542_concrete1_io_in_x473_bits_wdata_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x473_bits_wstrb; // @[sm_x542.scala 102:24:@39224.4]
  wire [20:0] x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_en_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure; // @[sm_x542.scala 102:24:@39224.4]
  wire [31:0] x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_output_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x474_ready; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_in_x474_valid; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x542.scala 102:24:@39224.4]
  wire  x542_kernelx542_concrete1_io_rr; // @[sm_x542.scala 102:24:@39224.4]
  wire  _T_266; // @[package.scala 100:49:@39153.4]
  reg  _T_269; // @[package.scala 48:56:@39154.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@39192.4 package.scala 96:25:@39193.4]
  wire  _T_289; // @[package.scala 96:25:@39200.4 package.scala 96:25:@39201.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@39203.4]
  x268_outbuf_0 x268_outbuf_0 ( // @[m_x268_outbuf_0.scala 27:17:@39062.4]
    .clock(x268_outbuf_0_clock),
    .reset(x268_outbuf_0_reset),
    .io_rPort_0_ofs_0(x268_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x268_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x268_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x268_outbuf_0_io_rPort_0_output_0)
  );
  x542_sm x542_sm ( // @[sm_x542.scala 37:18:@39120.4]
    .clock(x542_sm_clock),
    .reset(x542_sm_reset),
    .io_enable(x542_sm_io_enable),
    .io_done(x542_sm_io_done),
    .io_ctrDone(x542_sm_io_ctrDone),
    .io_ctrInc(x542_sm_io_ctrInc),
    .io_parentAck(x542_sm_io_parentAck),
    .io_doneIn_0(x542_sm_io_doneIn_0),
    .io_doneIn_1(x542_sm_io_doneIn_1),
    .io_enableOut_0(x542_sm_io_enableOut_0),
    .io_enableOut_1(x542_sm_io_enableOut_1),
    .io_childAck_0(x542_sm_io_childAck_0),
    .io_childAck_1(x542_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39187.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39195.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x542_kernelx542_concrete1 x542_kernelx542_concrete1 ( // @[sm_x542.scala 102:24:@39224.4]
    .clock(x542_kernelx542_concrete1_clock),
    .reset(x542_kernelx542_concrete1_reset),
    .io_in_x472_ready(x542_kernelx542_concrete1_io_in_x472_ready),
    .io_in_x472_valid(x542_kernelx542_concrete1_io_in_x472_valid),
    .io_in_x472_bits_addr(x542_kernelx542_concrete1_io_in_x472_bits_addr),
    .io_in_x472_bits_size(x542_kernelx542_concrete1_io_in_x472_bits_size),
    .io_in_x266_TVALID(x542_kernelx542_concrete1_io_in_x266_TVALID),
    .io_in_x266_TREADY(x542_kernelx542_concrete1_io_in_x266_TREADY),
    .io_in_x266_TDATA(x542_kernelx542_concrete1_io_in_x266_TDATA),
    .io_in_x266_TID(x542_kernelx542_concrete1_io_in_x266_TID),
    .io_in_x266_TDEST(x542_kernelx542_concrete1_io_in_x266_TDEST),
    .io_in_x264_outdram_number(x542_kernelx542_concrete1_io_in_x264_outdram_number),
    .io_in_x267_TVALID(x542_kernelx542_concrete1_io_in_x267_TVALID),
    .io_in_x267_TREADY(x542_kernelx542_concrete1_io_in_x267_TREADY),
    .io_in_x267_TDATA(x542_kernelx542_concrete1_io_in_x267_TDATA),
    .io_in_x473_ready(x542_kernelx542_concrete1_io_in_x473_ready),
    .io_in_x473_valid(x542_kernelx542_concrete1_io_in_x473_valid),
    .io_in_x473_bits_wdata_0(x542_kernelx542_concrete1_io_in_x473_bits_wdata_0),
    .io_in_x473_bits_wstrb(x542_kernelx542_concrete1_io_in_x473_bits_wstrb),
    .io_in_x268_outbuf_0_rPort_0_ofs_0(x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0),
    .io_in_x268_outbuf_0_rPort_0_en_0(x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_en_0),
    .io_in_x268_outbuf_0_rPort_0_backpressure(x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure),
    .io_in_x268_outbuf_0_rPort_0_output_0(x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_output_0),
    .io_in_x474_ready(x542_kernelx542_concrete1_io_in_x474_ready),
    .io_in_x474_valid(x542_kernelx542_concrete1_io_in_x474_valid),
    .io_sigsIn_smEnableOuts_0(x542_kernelx542_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x542_kernelx542_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x542_kernelx542_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x542_kernelx542_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x542_kernelx542_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x542_kernelx542_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x542_kernelx542_concrete1_io_rr)
  );
  assign _T_266 = x542_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39153.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@39192.4 package.scala 96:25:@39193.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39200.4 package.scala 96:25:@39201.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@39203.4]
  assign io_in_x472_valid = x542_kernelx542_concrete1_io_in_x472_valid; // @[sm_x542.scala 63:23:@39305.4]
  assign io_in_x472_bits_addr = x542_kernelx542_concrete1_io_in_x472_bits_addr; // @[sm_x542.scala 63:23:@39304.4]
  assign io_in_x472_bits_size = x542_kernelx542_concrete1_io_in_x472_bits_size; // @[sm_x542.scala 63:23:@39303.4]
  assign io_in_x266_TREADY = x542_kernelx542_concrete1_io_in_x266_TREADY; // @[sm_x542.scala 64:23:@39314.4]
  assign io_in_x267_TVALID = x542_kernelx542_concrete1_io_in_x267_TVALID; // @[sm_x542.scala 66:23:@39325.4]
  assign io_in_x267_TDATA = x542_kernelx542_concrete1_io_in_x267_TDATA; // @[sm_x542.scala 66:23:@39323.4]
  assign io_in_x473_valid = x542_kernelx542_concrete1_io_in_x473_valid; // @[sm_x542.scala 67:23:@39328.4]
  assign io_in_x473_bits_wdata_0 = x542_kernelx542_concrete1_io_in_x473_bits_wdata_0; // @[sm_x542.scala 67:23:@39327.4]
  assign io_in_x473_bits_wstrb = x542_kernelx542_concrete1_io_in_x473_bits_wstrb; // @[sm_x542.scala 67:23:@39326.4]
  assign io_in_x474_ready = x542_kernelx542_concrete1_io_in_x474_ready; // @[sm_x542.scala 69:23:@39337.4]
  assign io_sigsOut_smDoneIn_0 = x542_sm_io_done; // @[SpatialBlocks.scala 156:53:@39210.4]
  assign x268_outbuf_0_clock = clock; // @[:@39063.4]
  assign x268_outbuf_0_reset = reset; // @[:@39064.4]
  assign x268_outbuf_0_io_rPort_0_ofs_0 = x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@39333.4]
  assign x268_outbuf_0_io_rPort_0_en_0 = x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@39332.4]
  assign x268_outbuf_0_io_rPort_0_backpressure = x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@39331.4]
  assign x542_sm_clock = clock; // @[:@39121.4]
  assign x542_sm_reset = reset; // @[:@39122.4]
  assign x542_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@39207.4]
  assign x542_sm_io_ctrDone = x542_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@39157.4]
  assign x542_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@39209.4]
  assign x542_sm_io_doneIn_0 = x542_kernelx542_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@39177.4]
  assign x542_sm_io_doneIn_1 = x542_kernelx542_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@39178.4]
  assign RetimeWrapper_clock = clock; // @[:@39188.4]
  assign RetimeWrapper_reset = reset; // @[:@39189.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39191.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@39190.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39196.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39197.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39199.4]
  assign RetimeWrapper_1_io_in = x542_sm_io_done; // @[package.scala 94:16:@39198.4]
  assign x542_kernelx542_concrete1_clock = clock; // @[:@39225.4]
  assign x542_kernelx542_concrete1_reset = reset; // @[:@39226.4]
  assign x542_kernelx542_concrete1_io_in_x472_ready = io_in_x472_ready; // @[sm_x542.scala 63:23:@39306.4]
  assign x542_kernelx542_concrete1_io_in_x266_TVALID = io_in_x266_TVALID; // @[sm_x542.scala 64:23:@39315.4]
  assign x542_kernelx542_concrete1_io_in_x266_TDATA = io_in_x266_TDATA; // @[sm_x542.scala 64:23:@39313.4]
  assign x542_kernelx542_concrete1_io_in_x266_TID = io_in_x266_TID; // @[sm_x542.scala 64:23:@39309.4]
  assign x542_kernelx542_concrete1_io_in_x266_TDEST = io_in_x266_TDEST; // @[sm_x542.scala 64:23:@39308.4]
  assign x542_kernelx542_concrete1_io_in_x264_outdram_number = io_in_x264_outdram_number; // @[sm_x542.scala 65:31:@39316.4]
  assign x542_kernelx542_concrete1_io_in_x267_TREADY = io_in_x267_TREADY; // @[sm_x542.scala 66:23:@39324.4]
  assign x542_kernelx542_concrete1_io_in_x473_ready = io_in_x473_ready; // @[sm_x542.scala 67:23:@39329.4]
  assign x542_kernelx542_concrete1_io_in_x268_outbuf_0_rPort_0_output_0 = x268_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@39330.4]
  assign x542_kernelx542_concrete1_io_in_x474_valid = io_in_x474_valid; // @[sm_x542.scala 69:23:@39336.4]
  assign x542_kernelx542_concrete1_io_sigsIn_smEnableOuts_0 = x542_sm_io_enableOut_0; // @[sm_x542.scala 107:22:@39348.4]
  assign x542_kernelx542_concrete1_io_sigsIn_smEnableOuts_1 = x542_sm_io_enableOut_1; // @[sm_x542.scala 107:22:@39349.4]
  assign x542_kernelx542_concrete1_io_sigsIn_smChildAcks_0 = x542_sm_io_childAck_0; // @[sm_x542.scala 107:22:@39344.4]
  assign x542_kernelx542_concrete1_io_sigsIn_smChildAcks_1 = x542_sm_io_childAck_1; // @[sm_x542.scala 107:22:@39345.4]
  assign x542_kernelx542_concrete1_io_rr = io_rr; // @[sm_x542.scala 106:18:@39338.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@39371.2]
  input          clock, // @[:@39372.4]
  input          reset, // @[:@39373.4]
  input          io_enable, // @[:@39374.4]
  output         io_done, // @[:@39374.4]
  input          io_reset, // @[:@39374.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@39374.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@39374.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@39374.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@39374.4]
  output         io_memStreams_loads_0_data_ready, // @[:@39374.4]
  input          io_memStreams_loads_0_data_valid, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@39374.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@39374.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@39374.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@39374.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@39374.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@39374.4]
  input          io_memStreams_stores_0_data_ready, // @[:@39374.4]
  output         io_memStreams_stores_0_data_valid, // @[:@39374.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@39374.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@39374.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@39374.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@39374.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@39374.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@39374.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@39374.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@39374.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@39374.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@39374.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@39374.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@39374.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@39374.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@39374.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@39374.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@39374.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@39374.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@39374.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@39374.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@39374.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@39374.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@39374.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@39374.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@39374.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@39374.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@39374.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@39374.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@39374.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@39374.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@39374.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@39374.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@39374.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@39374.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@39374.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@39374.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@39374.4]
  output         io_heap_0_req_valid, // @[:@39374.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@39374.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@39374.4]
  input          io_heap_0_resp_valid, // @[:@39374.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@39374.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@39374.4]
  input  [63:0]  io_argIns_0, // @[:@39374.4]
  input  [63:0]  io_argIns_1, // @[:@39374.4]
  input          io_argOuts_0_port_ready, // @[:@39374.4]
  output         io_argOuts_0_port_valid, // @[:@39374.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@39374.4]
  input  [63:0]  io_argOuts_0_echo // @[:@39374.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@39522.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@39522.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@39522.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@39522.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39540.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39540.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@39549.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@39549.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@39549.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@39549.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@39549.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@39549.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@39588.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39620.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39620.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39620.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39620.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39620.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x472_ready; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x472_valid; // @[sm_RootController.scala 91:24:@39682.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x472_bits_addr; // @[sm_RootController.scala 91:24:@39682.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x472_bits_size; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x266_TVALID; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x266_TREADY; // @[sm_RootController.scala 91:24:@39682.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x266_TDATA; // @[sm_RootController.scala 91:24:@39682.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x266_TID; // @[sm_RootController.scala 91:24:@39682.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x266_TDEST; // @[sm_RootController.scala 91:24:@39682.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x264_outdram_number; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x267_TVALID; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x267_TREADY; // @[sm_RootController.scala 91:24:@39682.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x267_TDATA; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x473_ready; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x473_valid; // @[sm_RootController.scala 91:24:@39682.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x473_bits_wdata_0; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x473_bits_wstrb; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x474_ready; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_in_x474_valid; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@39682.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@39682.4]
  wire  _T_599; // @[package.scala 96:25:@39545.4 package.scala 96:25:@39546.4]
  wire  _T_664; // @[Main.scala 46:50:@39616.4]
  wire  _T_665; // @[Main.scala 46:59:@39617.4]
  wire  _T_677; // @[package.scala 100:49:@39637.4]
  reg  _T_680; // @[package.scala 48:56:@39638.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@39522.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39540.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@39549.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@39588.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39620.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@39682.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x472_ready(RootController_kernelRootController_concrete1_io_in_x472_ready),
    .io_in_x472_valid(RootController_kernelRootController_concrete1_io_in_x472_valid),
    .io_in_x472_bits_addr(RootController_kernelRootController_concrete1_io_in_x472_bits_addr),
    .io_in_x472_bits_size(RootController_kernelRootController_concrete1_io_in_x472_bits_size),
    .io_in_x266_TVALID(RootController_kernelRootController_concrete1_io_in_x266_TVALID),
    .io_in_x266_TREADY(RootController_kernelRootController_concrete1_io_in_x266_TREADY),
    .io_in_x266_TDATA(RootController_kernelRootController_concrete1_io_in_x266_TDATA),
    .io_in_x266_TID(RootController_kernelRootController_concrete1_io_in_x266_TID),
    .io_in_x266_TDEST(RootController_kernelRootController_concrete1_io_in_x266_TDEST),
    .io_in_x264_outdram_number(RootController_kernelRootController_concrete1_io_in_x264_outdram_number),
    .io_in_x267_TVALID(RootController_kernelRootController_concrete1_io_in_x267_TVALID),
    .io_in_x267_TREADY(RootController_kernelRootController_concrete1_io_in_x267_TREADY),
    .io_in_x267_TDATA(RootController_kernelRootController_concrete1_io_in_x267_TDATA),
    .io_in_x473_ready(RootController_kernelRootController_concrete1_io_in_x473_ready),
    .io_in_x473_valid(RootController_kernelRootController_concrete1_io_in_x473_valid),
    .io_in_x473_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x473_bits_wdata_0),
    .io_in_x473_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x473_bits_wstrb),
    .io_in_x474_ready(RootController_kernelRootController_concrete1_io_in_x474_ready),
    .io_in_x474_valid(RootController_kernelRootController_concrete1_io_in_x474_valid),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@39545.4 package.scala 96:25:@39546.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@39616.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@39617.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39637.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@39636.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x472_valid; // @[sm_RootController.scala 60:23:@39745.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x472_bits_addr; // @[sm_RootController.scala 60:23:@39744.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x472_bits_size; // @[sm_RootController.scala 60:23:@39743.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x473_valid; // @[sm_RootController.scala 64:23:@39768.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x473_bits_wdata_0; // @[sm_RootController.scala 64:23:@39767.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x473_bits_wstrb; // @[sm_RootController.scala 64:23:@39766.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x474_ready; // @[sm_RootController.scala 65:23:@39772.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x266_TREADY; // @[sm_RootController.scala 61:23:@39754.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x267_TVALID; // @[sm_RootController.scala 63:23:@39765.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x267_TDATA; // @[sm_RootController.scala 63:23:@39763.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 63:23:@39762.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 63:23:@39761.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 63:23:@39760.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 63:23:@39759.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 63:23:@39758.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 63:23:@39757.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@39523.4]
  assign SingleCounter_reset = reset; // @[:@39524.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@39538.4]
  assign RetimeWrapper_clock = clock; // @[:@39541.4]
  assign RetimeWrapper_reset = reset; // @[:@39542.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39544.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@39543.4]
  assign SRFF_clock = clock; // @[:@39550.4]
  assign SRFF_reset = reset; // @[:@39551.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@39800.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@39634.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@39635.4]
  assign RootController_sm_clock = clock; // @[:@39589.4]
  assign RootController_sm_reset = reset; // @[:@39590.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@39633.4 SpatialBlocks.scala 140:18:@39667.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@39661.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@39641.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@39629.4 SpatialBlocks.scala 142:21:@39669.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@39658.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39621.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39622.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39624.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@39623.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@39683.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@39684.4]
  assign RootController_kernelRootController_concrete1_io_in_x472_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 60:23:@39746.4]
  assign RootController_kernelRootController_concrete1_io_in_x266_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 61:23:@39755.4]
  assign RootController_kernelRootController_concrete1_io_in_x266_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 61:23:@39753.4]
  assign RootController_kernelRootController_concrete1_io_in_x266_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 61:23:@39749.4]
  assign RootController_kernelRootController_concrete1_io_in_x266_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 61:23:@39748.4]
  assign RootController_kernelRootController_concrete1_io_in_x264_outdram_number = io_argIns_1; // @[sm_RootController.scala 62:31:@39756.4]
  assign RootController_kernelRootController_concrete1_io_in_x267_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 63:23:@39764.4]
  assign RootController_kernelRootController_concrete1_io_in_x473_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 64:23:@39769.4]
  assign RootController_kernelRootController_concrete1_io_in_x474_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 65:23:@39771.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@39781.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@39779.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@39773.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@39802.2]
  input        clock, // @[:@39803.4]
  input        reset, // @[:@39804.4]
  input        io_enable, // @[:@39805.4]
  output [5:0] io_out, // @[:@39805.4]
  output [5:0] io_next // @[:@39805.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@39807.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@39808.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@39809.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@39814.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@39808.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@39809.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@39814.6]
  assign io_out = count; // @[Counter.scala 25:10:@39817.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@39818.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_33( // @[:@39854.2]
  input         clock, // @[:@39855.4]
  input         reset, // @[:@39856.4]
  input  [5:0]  io_raddr, // @[:@39857.4]
  input         io_wen, // @[:@39857.4]
  input  [5:0]  io_waddr, // @[:@39857.4]
  input  [63:0] io_wdata_addr, // @[:@39857.4]
  input  [31:0] io_wdata_size, // @[:@39857.4]
  output [63:0] io_rdata_addr, // @[:@39857.4]
  output [31:0] io_rdata_size // @[:@39857.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@39859.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@39859.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@39859.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@39859.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@39859.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@39859.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@39859.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@39859.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@39859.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@39873.4]
  wire  _T_20; // @[SRAM.scala 182:49:@39878.4]
  wire  _T_21; // @[SRAM.scala 182:37:@39879.4]
  reg  _T_24; // @[SRAM.scala 182:29:@39880.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@39883.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@39885.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@39859.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@39873.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@39878.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@39879.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@39885.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@39894.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@39893.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@39874.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@39875.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@39871.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@39877.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@39876.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@39872.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@39870.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@39869.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@39896.2]
  input         clock, // @[:@39897.4]
  input         reset, // @[:@39898.4]
  output        io_in_ready, // @[:@39899.4]
  input         io_in_valid, // @[:@39899.4]
  input  [63:0] io_in_bits_addr, // @[:@39899.4]
  input  [31:0] io_in_bits_size, // @[:@39899.4]
  input         io_out_ready, // @[:@39899.4]
  output        io_out_valid, // @[:@39899.4]
  output [63:0] io_out_bits_addr, // @[:@39899.4]
  output [31:0] io_out_bits_size // @[:@39899.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@40295.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@40295.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@40295.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@40295.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@40295.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@40305.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@40305.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@40305.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@40305.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@40305.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@40320.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@40320.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@40320.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@40320.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@40320.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@40320.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@40320.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@40320.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@40320.4]
  wire  writeEn; // @[FIFO.scala 30:29:@40293.4]
  wire  readEn; // @[FIFO.scala 31:29:@40294.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@40315.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@40316.4]
  wire  _T_824; // @[FIFO.scala 45:27:@40317.4]
  wire  empty; // @[FIFO.scala 45:24:@40318.4]
  wire  full; // @[FIFO.scala 46:23:@40319.4]
  wire  _T_827; // @[FIFO.scala 83:17:@40332.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@40333.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@40295.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@40305.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_33 SRAM ( // @[FIFO.scala 73:19:@40320.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@40293.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@40294.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@40316.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@40317.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@40318.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@40319.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@40332.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@40333.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@40339.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@40337.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@40330.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@40329.4]
  assign enqCounter_clock = clock; // @[:@40296.4]
  assign enqCounter_reset = reset; // @[:@40297.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@40303.4]
  assign deqCounter_clock = clock; // @[:@40306.4]
  assign deqCounter_reset = reset; // @[:@40307.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@40313.4]
  assign SRAM_clock = clock; // @[:@40321.4]
  assign SRAM_reset = reset; // @[:@40322.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@40324.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@40325.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@40326.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@40328.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@40327.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@40341.2]
  input        clock, // @[:@40342.4]
  input        reset, // @[:@40343.4]
  input        io_enable, // @[:@40344.4]
  output [3:0] io_out // @[:@40344.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@40346.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@40347.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@40348.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@40353.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@40347.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@40348.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@40353.6]
  assign io_out = count; // @[Counter.scala 25:10:@40356.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@40377.2]
  input        clock, // @[:@40378.4]
  input        reset, // @[:@40379.4]
  input        io_reset, // @[:@40380.4]
  input        io_enable, // @[:@40380.4]
  input  [1:0] io_stride, // @[:@40380.4]
  output [1:0] io_out, // @[:@40380.4]
  output [1:0] io_next // @[:@40380.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@40382.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@40383.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@40384.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@40389.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@40385.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@40383.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@40384.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@40389.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@40385.4]
  assign io_out = count; // @[Counter.scala 25:10:@40392.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@40393.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_34( // @[:@40429.2]
  input         clock, // @[:@40430.4]
  input         reset, // @[:@40431.4]
  input  [1:0]  io_raddr, // @[:@40432.4]
  input         io_wen, // @[:@40432.4]
  input  [1:0]  io_waddr, // @[:@40432.4]
  input  [31:0] io_wdata, // @[:@40432.4]
  output [31:0] io_rdata, // @[:@40432.4]
  input         io_backpressure // @[:@40432.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@40434.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@40434.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@40434.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@40434.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@40434.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@40434.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@40434.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@40434.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@40434.4]
  wire  _T_19; // @[SRAM.scala 182:49:@40452.4]
  wire  _T_20; // @[SRAM.scala 182:37:@40453.4]
  reg  _T_23; // @[SRAM.scala 182:29:@40454.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@40456.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@40434.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@40452.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@40453.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@40461.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@40448.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@40449.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@40446.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@40451.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@40450.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@40447.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@40445.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@40444.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@40463.2]
  input         clock, // @[:@40464.4]
  input         reset, // @[:@40465.4]
  output        io_in_ready, // @[:@40466.4]
  input         io_in_valid, // @[:@40466.4]
  input  [31:0] io_in_bits, // @[:@40466.4]
  input         io_out_ready, // @[:@40466.4]
  output        io_out_valid, // @[:@40466.4]
  output [31:0] io_out_bits // @[:@40466.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@40492.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@40492.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@40492.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@40492.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@40492.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@40492.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@40492.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@40502.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@40502.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@40502.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@40502.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@40502.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@40502.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@40502.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@40517.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@40517.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@40517.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@40517.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@40517.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@40517.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@40517.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@40517.4]
  wire  writeEn; // @[FIFO.scala 30:29:@40490.4]
  wire  readEn; // @[FIFO.scala 31:29:@40491.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@40512.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@40513.4]
  wire  _T_104; // @[FIFO.scala 45:27:@40514.4]
  wire  empty; // @[FIFO.scala 45:24:@40515.4]
  wire  full; // @[FIFO.scala 46:23:@40516.4]
  wire  _T_107; // @[FIFO.scala 83:17:@40527.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@40528.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@40492.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@40502.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_34 SRAM ( // @[FIFO.scala 73:19:@40517.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@40490.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@40491.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@40513.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@40514.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@40515.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@40516.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@40527.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@40528.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@40534.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@40532.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@40525.4]
  assign enqCounter_clock = clock; // @[:@40493.4]
  assign enqCounter_reset = reset; // @[:@40494.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@40500.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@40501.4]
  assign deqCounter_clock = clock; // @[:@40503.4]
  assign deqCounter_reset = reset; // @[:@40504.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@40510.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@40511.4]
  assign SRAM_clock = clock; // @[:@40518.4]
  assign SRAM_reset = reset; // @[:@40519.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@40521.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@40522.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@40523.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@40524.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@40526.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@42921.2]
  input         clock, // @[:@42922.4]
  input         reset, // @[:@42923.4]
  output        io_in_ready, // @[:@42924.4]
  input         io_in_valid, // @[:@42924.4]
  input  [31:0] io_in_bits_0, // @[:@42924.4]
  input         io_out_ready, // @[:@42924.4]
  output        io_out_valid, // @[:@42924.4]
  output [31:0] io_out_bits_0, // @[:@42924.4]
  output [31:0] io_out_bits_1, // @[:@42924.4]
  output [31:0] io_out_bits_2, // @[:@42924.4]
  output [31:0] io_out_bits_3, // @[:@42924.4]
  output [31:0] io_out_bits_4, // @[:@42924.4]
  output [31:0] io_out_bits_5, // @[:@42924.4]
  output [31:0] io_out_bits_6, // @[:@42924.4]
  output [31:0] io_out_bits_7, // @[:@42924.4]
  output [31:0] io_out_bits_8, // @[:@42924.4]
  output [31:0] io_out_bits_9, // @[:@42924.4]
  output [31:0] io_out_bits_10, // @[:@42924.4]
  output [31:0] io_out_bits_11, // @[:@42924.4]
  output [31:0] io_out_bits_12, // @[:@42924.4]
  output [31:0] io_out_bits_13, // @[:@42924.4]
  output [31:0] io_out_bits_14, // @[:@42924.4]
  output [31:0] io_out_bits_15 // @[:@42924.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@42928.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@42928.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@42928.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@42928.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@42939.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@42939.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@42939.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@42939.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@42952.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@42952.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@42987.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@42987.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@43022.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@43022.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@43057.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@43057.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@43092.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@43092.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@43127.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@43127.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@43162.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@43162.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@43162.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@43162.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@43162.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@43162.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@43162.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@43162.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@43197.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@43197.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@43197.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@43197.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@43197.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@43197.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@43197.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@43197.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@43232.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@43232.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@43232.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@43232.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@43232.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@43232.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@43232.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@43232.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@43267.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@43267.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@43267.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@43267.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@43267.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@43267.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@43267.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@43267.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@43302.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@43302.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@43302.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@43302.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@43302.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@43302.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@43302.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@43302.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@43337.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@43337.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@43337.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@43337.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@43337.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@43337.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@43337.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@43337.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@43372.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@43372.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@43372.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@43372.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@43372.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@43372.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@43372.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@43372.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@43407.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@43407.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@43407.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@43407.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@43407.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@43407.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@43407.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@43407.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@43442.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@43442.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@43442.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@43442.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@43442.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@43442.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@43442.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@43442.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@43477.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@43477.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@43477.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@43477.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@43477.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@43477.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@43477.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@43477.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@42927.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@42950.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@42977.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@43012.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@43047.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@43082.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@43117.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@43152.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@43187.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@43222.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@43257.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@43292.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@43327.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@43362.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@43397.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@43432.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@43467.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@43502.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43513.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43514.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43515.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43516.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43517.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43518.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43519.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43520.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43521.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43522.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43523.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43524.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43525.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43526.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43527.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@43544.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43528.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@43563.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@43564.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@43565.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@43566.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@43567.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@43568.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@43569.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@43570.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@43571.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@43572.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@43573.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@43574.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@43575.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@43576.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@42928.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@42939.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@42952.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@42987.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@43022.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@43057.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@43092.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@43127.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@43162.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@43197.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@43232.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@43267.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@43302.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@43337.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@43372.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@43407.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@43442.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@43477.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@42927.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@42950.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@42977.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@43012.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@43047.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@43082.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@43117.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@43152.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@43187.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@43222.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@43257.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@43292.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@43327.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@43362.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@43397.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@43432.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@43467.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@43502.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43513.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43514.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43515.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43516.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43517.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43518.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43519.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43520.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43521.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43522.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43523.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43524.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43525.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43526.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43527.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@43544.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@43512.4 FIFOVec.scala 49:42:@43528.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@43563.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@43564.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@43565.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@43566.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@43567.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@43568.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@43569.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@43570.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@43571.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@43572.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@43573.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@43574.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@43575.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@43576.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@43545.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@43579.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@43887.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@43888.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@43889.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@43890.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@43891.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@43892.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@43893.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@43894.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@43895.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@43896.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@43897.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@43898.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@43899.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@43900.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@43901.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@43902.4]
  assign enqCounter_clock = clock; // @[:@42929.4]
  assign enqCounter_reset = reset; // @[:@42930.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@42937.4]
  assign deqCounter_clock = clock; // @[:@42940.4]
  assign deqCounter_reset = reset; // @[:@42941.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@42948.4]
  assign fifos_0_clock = clock; // @[:@42953.4]
  assign fifos_0_reset = reset; // @[:@42954.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@42980.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42982.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42986.4]
  assign fifos_1_clock = clock; // @[:@42988.4]
  assign fifos_1_reset = reset; // @[:@42989.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@43015.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43017.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43021.4]
  assign fifos_2_clock = clock; // @[:@43023.4]
  assign fifos_2_reset = reset; // @[:@43024.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@43050.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43052.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43056.4]
  assign fifos_3_clock = clock; // @[:@43058.4]
  assign fifos_3_reset = reset; // @[:@43059.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@43085.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43087.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43091.4]
  assign fifos_4_clock = clock; // @[:@43093.4]
  assign fifos_4_reset = reset; // @[:@43094.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@43120.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43122.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43126.4]
  assign fifos_5_clock = clock; // @[:@43128.4]
  assign fifos_5_reset = reset; // @[:@43129.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@43155.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43157.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43161.4]
  assign fifos_6_clock = clock; // @[:@43163.4]
  assign fifos_6_reset = reset; // @[:@43164.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@43190.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43192.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43196.4]
  assign fifos_7_clock = clock; // @[:@43198.4]
  assign fifos_7_reset = reset; // @[:@43199.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@43225.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43227.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43231.4]
  assign fifos_8_clock = clock; // @[:@43233.4]
  assign fifos_8_reset = reset; // @[:@43234.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@43260.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43262.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43266.4]
  assign fifos_9_clock = clock; // @[:@43268.4]
  assign fifos_9_reset = reset; // @[:@43269.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@43295.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43297.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43301.4]
  assign fifos_10_clock = clock; // @[:@43303.4]
  assign fifos_10_reset = reset; // @[:@43304.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@43330.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43332.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43336.4]
  assign fifos_11_clock = clock; // @[:@43338.4]
  assign fifos_11_reset = reset; // @[:@43339.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@43365.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43367.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43371.4]
  assign fifos_12_clock = clock; // @[:@43373.4]
  assign fifos_12_reset = reset; // @[:@43374.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@43400.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43402.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43406.4]
  assign fifos_13_clock = clock; // @[:@43408.4]
  assign fifos_13_reset = reset; // @[:@43409.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@43435.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43437.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43441.4]
  assign fifos_14_clock = clock; // @[:@43443.4]
  assign fifos_14_reset = reset; // @[:@43444.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@43470.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43472.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43476.4]
  assign fifos_15_clock = clock; // @[:@43478.4]
  assign fifos_15_reset = reset; // @[:@43479.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@43505.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43507.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43511.4]
endmodule
module FFRAM( // @[:@43976.2]
  input        clock, // @[:@43977.4]
  input        reset, // @[:@43978.4]
  input  [1:0] io_raddr, // @[:@43979.4]
  input        io_wen, // @[:@43979.4]
  input  [1:0] io_waddr, // @[:@43979.4]
  input        io_wdata, // @[:@43979.4]
  output       io_rdata, // @[:@43979.4]
  input        io_banks_0_wdata_valid, // @[:@43979.4]
  input        io_banks_0_wdata_bits, // @[:@43979.4]
  input        io_banks_1_wdata_valid, // @[:@43979.4]
  input        io_banks_1_wdata_bits, // @[:@43979.4]
  input        io_banks_2_wdata_valid, // @[:@43979.4]
  input        io_banks_2_wdata_bits, // @[:@43979.4]
  input        io_banks_3_wdata_valid, // @[:@43979.4]
  input        io_banks_3_wdata_bits // @[:@43979.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@43983.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@43984.4]
  wire  _T_89; // @[SRAM.scala 148:25:@43985.4]
  wire  _T_90; // @[SRAM.scala 148:15:@43986.4]
  wire  _T_91; // @[SRAM.scala 149:15:@43988.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@43987.4]
  reg  regs_1; // @[SRAM.scala 145:20:@43994.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@43995.4]
  wire  _T_98; // @[SRAM.scala 148:25:@43996.4]
  wire  _T_99; // @[SRAM.scala 148:15:@43997.4]
  wire  _T_100; // @[SRAM.scala 149:15:@43999.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@43998.4]
  reg  regs_2; // @[SRAM.scala 145:20:@44005.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@44006.4]
  wire  _T_107; // @[SRAM.scala 148:25:@44007.4]
  wire  _T_108; // @[SRAM.scala 148:15:@44008.4]
  wire  _T_109; // @[SRAM.scala 149:15:@44010.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@44009.4]
  reg  regs_3; // @[SRAM.scala 145:20:@44016.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@44017.4]
  wire  _T_116; // @[SRAM.scala 148:25:@44018.4]
  wire  _T_117; // @[SRAM.scala 148:15:@44019.4]
  wire  _T_118; // @[SRAM.scala 149:15:@44021.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@44020.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@44030.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@44030.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@43984.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@43985.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@43986.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43988.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@43987.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@43995.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@43996.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@43997.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43999.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@43998.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@44006.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@44007.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@44008.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44010.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@44009.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@44017.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@44018.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@44019.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44021.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@44020.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@44030.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@44030.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@44030.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@44032.2]
  input   clock, // @[:@44033.4]
  input   reset, // @[:@44034.4]
  output  io_in_ready, // @[:@44035.4]
  input   io_in_valid, // @[:@44035.4]
  input   io_in_bits, // @[:@44035.4]
  input   io_out_ready, // @[:@44035.4]
  output  io_out_valid, // @[:@44035.4]
  output  io_out_bits // @[:@44035.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@44061.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@44061.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@44061.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@44061.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@44061.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@44061.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@44061.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@44071.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@44071.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@44071.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@44071.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@44071.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@44071.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@44071.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@44086.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@44086.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@44086.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@44086.4]
  wire  writeEn; // @[FIFO.scala 30:29:@44059.4]
  wire  readEn; // @[FIFO.scala 31:29:@44060.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@44081.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@44082.4]
  wire  _T_104; // @[FIFO.scala 45:27:@44083.4]
  wire  empty; // @[FIFO.scala 45:24:@44084.4]
  wire  full; // @[FIFO.scala 46:23:@44085.4]
  wire  _T_157; // @[FIFO.scala 83:17:@44172.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@44173.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@44061.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@44071.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@44086.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@44059.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@44060.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@44082.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@44083.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@44084.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@44085.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@44172.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@44173.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@44179.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@44177.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@44111.4]
  assign enqCounter_clock = clock; // @[:@44062.4]
  assign enqCounter_reset = reset; // @[:@44063.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@44069.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@44070.4]
  assign deqCounter_clock = clock; // @[:@44072.4]
  assign deqCounter_reset = reset; // @[:@44073.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@44079.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@44080.4]
  assign FFRAM_clock = clock; // @[:@44087.4]
  assign FFRAM_reset = reset; // @[:@44088.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@44107.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@44108.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@44109.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@44110.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44113.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44112.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44116.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44115.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44119.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44118.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@44122.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@44121.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@47796.2]
  input   clock, // @[:@47797.4]
  input   reset, // @[:@47798.4]
  output  io_in_ready, // @[:@47799.4]
  input   io_in_valid, // @[:@47799.4]
  input   io_in_bits_0, // @[:@47799.4]
  input   io_out_ready, // @[:@47799.4]
  output  io_out_valid, // @[:@47799.4]
  output  io_out_bits_0, // @[:@47799.4]
  output  io_out_bits_1, // @[:@47799.4]
  output  io_out_bits_2, // @[:@47799.4]
  output  io_out_bits_3, // @[:@47799.4]
  output  io_out_bits_4, // @[:@47799.4]
  output  io_out_bits_5, // @[:@47799.4]
  output  io_out_bits_6, // @[:@47799.4]
  output  io_out_bits_7, // @[:@47799.4]
  output  io_out_bits_8, // @[:@47799.4]
  output  io_out_bits_9, // @[:@47799.4]
  output  io_out_bits_10, // @[:@47799.4]
  output  io_out_bits_11, // @[:@47799.4]
  output  io_out_bits_12, // @[:@47799.4]
  output  io_out_bits_13, // @[:@47799.4]
  output  io_out_bits_14, // @[:@47799.4]
  output  io_out_bits_15 // @[:@47799.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@47803.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@47803.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@47803.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@47803.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@47814.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@47814.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@47814.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@47814.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@47827.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@47862.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@47897.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@47932.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@47967.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@48002.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@48037.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@48072.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@48107.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@48142.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@48177.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@48212.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@48247.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@48282.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@48317.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@48352.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@48352.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@47802.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@47825.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@47852.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@47887.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@47922.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@47957.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@47992.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@48027.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@48062.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@48097.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@48132.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@48167.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@48202.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@48237.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@48272.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@48307.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@48342.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@48377.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48388.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48389.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48390.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48391.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48392.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48393.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48394.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48395.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48396.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48397.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48398.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48399.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48400.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48401.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48402.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@48419.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48403.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@48438.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@48439.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@48440.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@48441.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@48442.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@48443.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@48444.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@48445.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@48446.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@48447.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@48448.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@48449.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@48450.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@48451.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@47803.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@47814.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@47827.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@47862.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@47897.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@47932.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@47967.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@48002.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@48037.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@48072.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@48107.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@48142.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@48177.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@48212.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@48247.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@48282.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@48317.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@48352.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@47802.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@47825.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@47852.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@47887.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@47922.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@47957.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@47992.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@48027.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@48062.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@48097.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@48132.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@48167.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@48202.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@48237.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@48272.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@48307.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@48342.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@48377.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48388.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48389.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48390.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48391.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48392.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48393.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48394.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48395.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48396.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48397.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48398.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48399.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48400.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48401.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48402.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@48419.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@48387.4 FIFOVec.scala 49:42:@48403.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@48438.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@48439.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@48440.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@48441.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@48442.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@48443.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@48444.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@48445.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@48446.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@48447.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@48448.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@48449.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@48450.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@48451.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@48420.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@48454.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@48762.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@48763.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@48764.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@48765.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@48766.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@48767.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@48768.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@48769.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@48770.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@48771.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@48772.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@48773.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@48774.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@48775.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@48776.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@48777.4]
  assign enqCounter_clock = clock; // @[:@47804.4]
  assign enqCounter_reset = reset; // @[:@47805.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@47812.4]
  assign deqCounter_clock = clock; // @[:@47815.4]
  assign deqCounter_reset = reset; // @[:@47816.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@47823.4]
  assign fifos_0_clock = clock; // @[:@47828.4]
  assign fifos_0_reset = reset; // @[:@47829.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@47855.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@47857.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@47861.4]
  assign fifos_1_clock = clock; // @[:@47863.4]
  assign fifos_1_reset = reset; // @[:@47864.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@47890.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@47892.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@47896.4]
  assign fifos_2_clock = clock; // @[:@47898.4]
  assign fifos_2_reset = reset; // @[:@47899.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@47925.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@47927.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@47931.4]
  assign fifos_3_clock = clock; // @[:@47933.4]
  assign fifos_3_reset = reset; // @[:@47934.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@47960.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@47962.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@47966.4]
  assign fifos_4_clock = clock; // @[:@47968.4]
  assign fifos_4_reset = reset; // @[:@47969.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@47995.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@47997.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48001.4]
  assign fifos_5_clock = clock; // @[:@48003.4]
  assign fifos_5_reset = reset; // @[:@48004.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@48030.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48032.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48036.4]
  assign fifos_6_clock = clock; // @[:@48038.4]
  assign fifos_6_reset = reset; // @[:@48039.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@48065.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48067.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48071.4]
  assign fifos_7_clock = clock; // @[:@48073.4]
  assign fifos_7_reset = reset; // @[:@48074.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@48100.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48102.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48106.4]
  assign fifos_8_clock = clock; // @[:@48108.4]
  assign fifos_8_reset = reset; // @[:@48109.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@48135.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48137.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48141.4]
  assign fifos_9_clock = clock; // @[:@48143.4]
  assign fifos_9_reset = reset; // @[:@48144.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@48170.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48172.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48176.4]
  assign fifos_10_clock = clock; // @[:@48178.4]
  assign fifos_10_reset = reset; // @[:@48179.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@48205.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48207.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48211.4]
  assign fifos_11_clock = clock; // @[:@48213.4]
  assign fifos_11_reset = reset; // @[:@48214.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@48240.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48242.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48246.4]
  assign fifos_12_clock = clock; // @[:@48248.4]
  assign fifos_12_reset = reset; // @[:@48249.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@48275.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48277.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48281.4]
  assign fifos_13_clock = clock; // @[:@48283.4]
  assign fifos_13_reset = reset; // @[:@48284.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@48310.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48312.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48316.4]
  assign fifos_14_clock = clock; // @[:@48318.4]
  assign fifos_14_reset = reset; // @[:@48319.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@48345.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48347.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48351.4]
  assign fifos_15_clock = clock; // @[:@48353.4]
  assign fifos_15_reset = reset; // @[:@48354.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@48380.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@48382.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@48386.4]
endmodule
module FIFOWidthConvert( // @[:@48779.2]
  input         clock, // @[:@48780.4]
  input         reset, // @[:@48781.4]
  output        io_in_ready, // @[:@48782.4]
  input         io_in_valid, // @[:@48782.4]
  input  [31:0] io_in_bits_data_0, // @[:@48782.4]
  input         io_in_bits_strobe, // @[:@48782.4]
  input         io_out_ready, // @[:@48782.4]
  output        io_out_valid, // @[:@48782.4]
  output [31:0] io_out_bits_data_0, // @[:@48782.4]
  output [31:0] io_out_bits_data_1, // @[:@48782.4]
  output [31:0] io_out_bits_data_2, // @[:@48782.4]
  output [31:0] io_out_bits_data_3, // @[:@48782.4]
  output [31:0] io_out_bits_data_4, // @[:@48782.4]
  output [31:0] io_out_bits_data_5, // @[:@48782.4]
  output [31:0] io_out_bits_data_6, // @[:@48782.4]
  output [31:0] io_out_bits_data_7, // @[:@48782.4]
  output [31:0] io_out_bits_data_8, // @[:@48782.4]
  output [31:0] io_out_bits_data_9, // @[:@48782.4]
  output [31:0] io_out_bits_data_10, // @[:@48782.4]
  output [31:0] io_out_bits_data_11, // @[:@48782.4]
  output [31:0] io_out_bits_data_12, // @[:@48782.4]
  output [31:0] io_out_bits_data_13, // @[:@48782.4]
  output [31:0] io_out_bits_data_14, // @[:@48782.4]
  output [31:0] io_out_bits_data_15, // @[:@48782.4]
  output [63:0] io_out_bits_strobe // @[:@48782.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@48784.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@48825.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@48884.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@48890.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@48948.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@48954.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@48955.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@48959.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@48963.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@48967.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@48971.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@48975.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@48979.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@48983.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@48987.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@48991.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@48995.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@48999.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@49003.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@49007.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@49011.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@49015.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@49092.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@49101.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@49110.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@49119.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@49128.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@49137.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@49145.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@48784.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@48825.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@48884.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@48890.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@48948.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@48954.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@48955.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@48959.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@48963.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@48967.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@48971.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@48975.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@48979.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@48983.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@48987.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@48991.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@48995.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@48999.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@49003.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@49007.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@49011.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@49015.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@49092.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@49101.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@49110.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@49119.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@49128.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@49137.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@49145.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@48874.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@48875.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@48924.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@48925.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@48926.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@48927.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@48928.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@48929.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@48930.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@48931.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@48932.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@48933.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@48934.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@48935.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@48936.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@48937.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@48938.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@48939.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@49147.4]
  assign FIFOVec_clock = clock; // @[:@48785.4]
  assign FIFOVec_reset = reset; // @[:@48786.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@48871.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@48870.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@49148.4]
  assign FIFOVec_1_clock = clock; // @[:@48826.4]
  assign FIFOVec_1_reset = reset; // @[:@48827.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@48873.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@48872.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@49149.4]
endmodule
module FFRAM_16( // @[:@49187.2]
  input        clock, // @[:@49188.4]
  input        reset, // @[:@49189.4]
  input  [5:0] io_raddr, // @[:@49190.4]
  input        io_wen, // @[:@49190.4]
  input  [5:0] io_waddr, // @[:@49190.4]
  input        io_wdata, // @[:@49190.4]
  output       io_rdata, // @[:@49190.4]
  input        io_banks_0_wdata_valid, // @[:@49190.4]
  input        io_banks_0_wdata_bits, // @[:@49190.4]
  input        io_banks_1_wdata_valid, // @[:@49190.4]
  input        io_banks_1_wdata_bits, // @[:@49190.4]
  input        io_banks_2_wdata_valid, // @[:@49190.4]
  input        io_banks_2_wdata_bits, // @[:@49190.4]
  input        io_banks_3_wdata_valid, // @[:@49190.4]
  input        io_banks_3_wdata_bits, // @[:@49190.4]
  input        io_banks_4_wdata_valid, // @[:@49190.4]
  input        io_banks_4_wdata_bits, // @[:@49190.4]
  input        io_banks_5_wdata_valid, // @[:@49190.4]
  input        io_banks_5_wdata_bits, // @[:@49190.4]
  input        io_banks_6_wdata_valid, // @[:@49190.4]
  input        io_banks_6_wdata_bits, // @[:@49190.4]
  input        io_banks_7_wdata_valid, // @[:@49190.4]
  input        io_banks_7_wdata_bits, // @[:@49190.4]
  input        io_banks_8_wdata_valid, // @[:@49190.4]
  input        io_banks_8_wdata_bits, // @[:@49190.4]
  input        io_banks_9_wdata_valid, // @[:@49190.4]
  input        io_banks_9_wdata_bits, // @[:@49190.4]
  input        io_banks_10_wdata_valid, // @[:@49190.4]
  input        io_banks_10_wdata_bits, // @[:@49190.4]
  input        io_banks_11_wdata_valid, // @[:@49190.4]
  input        io_banks_11_wdata_bits, // @[:@49190.4]
  input        io_banks_12_wdata_valid, // @[:@49190.4]
  input        io_banks_12_wdata_bits, // @[:@49190.4]
  input        io_banks_13_wdata_valid, // @[:@49190.4]
  input        io_banks_13_wdata_bits, // @[:@49190.4]
  input        io_banks_14_wdata_valid, // @[:@49190.4]
  input        io_banks_14_wdata_bits, // @[:@49190.4]
  input        io_banks_15_wdata_valid, // @[:@49190.4]
  input        io_banks_15_wdata_bits, // @[:@49190.4]
  input        io_banks_16_wdata_valid, // @[:@49190.4]
  input        io_banks_16_wdata_bits, // @[:@49190.4]
  input        io_banks_17_wdata_valid, // @[:@49190.4]
  input        io_banks_17_wdata_bits, // @[:@49190.4]
  input        io_banks_18_wdata_valid, // @[:@49190.4]
  input        io_banks_18_wdata_bits, // @[:@49190.4]
  input        io_banks_19_wdata_valid, // @[:@49190.4]
  input        io_banks_19_wdata_bits, // @[:@49190.4]
  input        io_banks_20_wdata_valid, // @[:@49190.4]
  input        io_banks_20_wdata_bits, // @[:@49190.4]
  input        io_banks_21_wdata_valid, // @[:@49190.4]
  input        io_banks_21_wdata_bits, // @[:@49190.4]
  input        io_banks_22_wdata_valid, // @[:@49190.4]
  input        io_banks_22_wdata_bits, // @[:@49190.4]
  input        io_banks_23_wdata_valid, // @[:@49190.4]
  input        io_banks_23_wdata_bits, // @[:@49190.4]
  input        io_banks_24_wdata_valid, // @[:@49190.4]
  input        io_banks_24_wdata_bits, // @[:@49190.4]
  input        io_banks_25_wdata_valid, // @[:@49190.4]
  input        io_banks_25_wdata_bits, // @[:@49190.4]
  input        io_banks_26_wdata_valid, // @[:@49190.4]
  input        io_banks_26_wdata_bits, // @[:@49190.4]
  input        io_banks_27_wdata_valid, // @[:@49190.4]
  input        io_banks_27_wdata_bits, // @[:@49190.4]
  input        io_banks_28_wdata_valid, // @[:@49190.4]
  input        io_banks_28_wdata_bits, // @[:@49190.4]
  input        io_banks_29_wdata_valid, // @[:@49190.4]
  input        io_banks_29_wdata_bits, // @[:@49190.4]
  input        io_banks_30_wdata_valid, // @[:@49190.4]
  input        io_banks_30_wdata_bits, // @[:@49190.4]
  input        io_banks_31_wdata_valid, // @[:@49190.4]
  input        io_banks_31_wdata_bits, // @[:@49190.4]
  input        io_banks_32_wdata_valid, // @[:@49190.4]
  input        io_banks_32_wdata_bits, // @[:@49190.4]
  input        io_banks_33_wdata_valid, // @[:@49190.4]
  input        io_banks_33_wdata_bits, // @[:@49190.4]
  input        io_banks_34_wdata_valid, // @[:@49190.4]
  input        io_banks_34_wdata_bits, // @[:@49190.4]
  input        io_banks_35_wdata_valid, // @[:@49190.4]
  input        io_banks_35_wdata_bits, // @[:@49190.4]
  input        io_banks_36_wdata_valid, // @[:@49190.4]
  input        io_banks_36_wdata_bits, // @[:@49190.4]
  input        io_banks_37_wdata_valid, // @[:@49190.4]
  input        io_banks_37_wdata_bits, // @[:@49190.4]
  input        io_banks_38_wdata_valid, // @[:@49190.4]
  input        io_banks_38_wdata_bits, // @[:@49190.4]
  input        io_banks_39_wdata_valid, // @[:@49190.4]
  input        io_banks_39_wdata_bits, // @[:@49190.4]
  input        io_banks_40_wdata_valid, // @[:@49190.4]
  input        io_banks_40_wdata_bits, // @[:@49190.4]
  input        io_banks_41_wdata_valid, // @[:@49190.4]
  input        io_banks_41_wdata_bits, // @[:@49190.4]
  input        io_banks_42_wdata_valid, // @[:@49190.4]
  input        io_banks_42_wdata_bits, // @[:@49190.4]
  input        io_banks_43_wdata_valid, // @[:@49190.4]
  input        io_banks_43_wdata_bits, // @[:@49190.4]
  input        io_banks_44_wdata_valid, // @[:@49190.4]
  input        io_banks_44_wdata_bits, // @[:@49190.4]
  input        io_banks_45_wdata_valid, // @[:@49190.4]
  input        io_banks_45_wdata_bits, // @[:@49190.4]
  input        io_banks_46_wdata_valid, // @[:@49190.4]
  input        io_banks_46_wdata_bits, // @[:@49190.4]
  input        io_banks_47_wdata_valid, // @[:@49190.4]
  input        io_banks_47_wdata_bits, // @[:@49190.4]
  input        io_banks_48_wdata_valid, // @[:@49190.4]
  input        io_banks_48_wdata_bits, // @[:@49190.4]
  input        io_banks_49_wdata_valid, // @[:@49190.4]
  input        io_banks_49_wdata_bits, // @[:@49190.4]
  input        io_banks_50_wdata_valid, // @[:@49190.4]
  input        io_banks_50_wdata_bits, // @[:@49190.4]
  input        io_banks_51_wdata_valid, // @[:@49190.4]
  input        io_banks_51_wdata_bits, // @[:@49190.4]
  input        io_banks_52_wdata_valid, // @[:@49190.4]
  input        io_banks_52_wdata_bits, // @[:@49190.4]
  input        io_banks_53_wdata_valid, // @[:@49190.4]
  input        io_banks_53_wdata_bits, // @[:@49190.4]
  input        io_banks_54_wdata_valid, // @[:@49190.4]
  input        io_banks_54_wdata_bits, // @[:@49190.4]
  input        io_banks_55_wdata_valid, // @[:@49190.4]
  input        io_banks_55_wdata_bits, // @[:@49190.4]
  input        io_banks_56_wdata_valid, // @[:@49190.4]
  input        io_banks_56_wdata_bits, // @[:@49190.4]
  input        io_banks_57_wdata_valid, // @[:@49190.4]
  input        io_banks_57_wdata_bits, // @[:@49190.4]
  input        io_banks_58_wdata_valid, // @[:@49190.4]
  input        io_banks_58_wdata_bits, // @[:@49190.4]
  input        io_banks_59_wdata_valid, // @[:@49190.4]
  input        io_banks_59_wdata_bits, // @[:@49190.4]
  input        io_banks_60_wdata_valid, // @[:@49190.4]
  input        io_banks_60_wdata_bits, // @[:@49190.4]
  input        io_banks_61_wdata_valid, // @[:@49190.4]
  input        io_banks_61_wdata_bits, // @[:@49190.4]
  input        io_banks_62_wdata_valid, // @[:@49190.4]
  input        io_banks_62_wdata_bits, // @[:@49190.4]
  input        io_banks_63_wdata_valid, // @[:@49190.4]
  input        io_banks_63_wdata_bits // @[:@49190.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@49194.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@49195.4]
  wire  _T_689; // @[SRAM.scala 148:25:@49196.4]
  wire  _T_690; // @[SRAM.scala 148:15:@49197.4]
  wire  _T_691; // @[SRAM.scala 149:15:@49199.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@49198.4]
  reg  regs_1; // @[SRAM.scala 145:20:@49205.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@49206.4]
  wire  _T_698; // @[SRAM.scala 148:25:@49207.4]
  wire  _T_699; // @[SRAM.scala 148:15:@49208.4]
  wire  _T_700; // @[SRAM.scala 149:15:@49210.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@49209.4]
  reg  regs_2; // @[SRAM.scala 145:20:@49216.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@49217.4]
  wire  _T_707; // @[SRAM.scala 148:25:@49218.4]
  wire  _T_708; // @[SRAM.scala 148:15:@49219.4]
  wire  _T_709; // @[SRAM.scala 149:15:@49221.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@49220.4]
  reg  regs_3; // @[SRAM.scala 145:20:@49227.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@49228.4]
  wire  _T_716; // @[SRAM.scala 148:25:@49229.4]
  wire  _T_717; // @[SRAM.scala 148:15:@49230.4]
  wire  _T_718; // @[SRAM.scala 149:15:@49232.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@49231.4]
  reg  regs_4; // @[SRAM.scala 145:20:@49238.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@49239.4]
  wire  _T_725; // @[SRAM.scala 148:25:@49240.4]
  wire  _T_726; // @[SRAM.scala 148:15:@49241.4]
  wire  _T_727; // @[SRAM.scala 149:15:@49243.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@49242.4]
  reg  regs_5; // @[SRAM.scala 145:20:@49249.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@49250.4]
  wire  _T_734; // @[SRAM.scala 148:25:@49251.4]
  wire  _T_735; // @[SRAM.scala 148:15:@49252.4]
  wire  _T_736; // @[SRAM.scala 149:15:@49254.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@49253.4]
  reg  regs_6; // @[SRAM.scala 145:20:@49260.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@49261.4]
  wire  _T_743; // @[SRAM.scala 148:25:@49262.4]
  wire  _T_744; // @[SRAM.scala 148:15:@49263.4]
  wire  _T_745; // @[SRAM.scala 149:15:@49265.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@49264.4]
  reg  regs_7; // @[SRAM.scala 145:20:@49271.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@49272.4]
  wire  _T_752; // @[SRAM.scala 148:25:@49273.4]
  wire  _T_753; // @[SRAM.scala 148:15:@49274.4]
  wire  _T_754; // @[SRAM.scala 149:15:@49276.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@49275.4]
  reg  regs_8; // @[SRAM.scala 145:20:@49282.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@49283.4]
  wire  _T_761; // @[SRAM.scala 148:25:@49284.4]
  wire  _T_762; // @[SRAM.scala 148:15:@49285.4]
  wire  _T_763; // @[SRAM.scala 149:15:@49287.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@49286.4]
  reg  regs_9; // @[SRAM.scala 145:20:@49293.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@49294.4]
  wire  _T_770; // @[SRAM.scala 148:25:@49295.4]
  wire  _T_771; // @[SRAM.scala 148:15:@49296.4]
  wire  _T_772; // @[SRAM.scala 149:15:@49298.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@49297.4]
  reg  regs_10; // @[SRAM.scala 145:20:@49304.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@49305.4]
  wire  _T_779; // @[SRAM.scala 148:25:@49306.4]
  wire  _T_780; // @[SRAM.scala 148:15:@49307.4]
  wire  _T_781; // @[SRAM.scala 149:15:@49309.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@49308.4]
  reg  regs_11; // @[SRAM.scala 145:20:@49315.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@49316.4]
  wire  _T_788; // @[SRAM.scala 148:25:@49317.4]
  wire  _T_789; // @[SRAM.scala 148:15:@49318.4]
  wire  _T_790; // @[SRAM.scala 149:15:@49320.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@49319.4]
  reg  regs_12; // @[SRAM.scala 145:20:@49326.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@49327.4]
  wire  _T_797; // @[SRAM.scala 148:25:@49328.4]
  wire  _T_798; // @[SRAM.scala 148:15:@49329.4]
  wire  _T_799; // @[SRAM.scala 149:15:@49331.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@49330.4]
  reg  regs_13; // @[SRAM.scala 145:20:@49337.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@49338.4]
  wire  _T_806; // @[SRAM.scala 148:25:@49339.4]
  wire  _T_807; // @[SRAM.scala 148:15:@49340.4]
  wire  _T_808; // @[SRAM.scala 149:15:@49342.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@49341.4]
  reg  regs_14; // @[SRAM.scala 145:20:@49348.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@49349.4]
  wire  _T_815; // @[SRAM.scala 148:25:@49350.4]
  wire  _T_816; // @[SRAM.scala 148:15:@49351.4]
  wire  _T_817; // @[SRAM.scala 149:15:@49353.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@49352.4]
  reg  regs_15; // @[SRAM.scala 145:20:@49359.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@49360.4]
  wire  _T_824; // @[SRAM.scala 148:25:@49361.4]
  wire  _T_825; // @[SRAM.scala 148:15:@49362.4]
  wire  _T_826; // @[SRAM.scala 149:15:@49364.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@49363.4]
  reg  regs_16; // @[SRAM.scala 145:20:@49370.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@49371.4]
  wire  _T_833; // @[SRAM.scala 148:25:@49372.4]
  wire  _T_834; // @[SRAM.scala 148:15:@49373.4]
  wire  _T_835; // @[SRAM.scala 149:15:@49375.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@49374.4]
  reg  regs_17; // @[SRAM.scala 145:20:@49381.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@49382.4]
  wire  _T_842; // @[SRAM.scala 148:25:@49383.4]
  wire  _T_843; // @[SRAM.scala 148:15:@49384.4]
  wire  _T_844; // @[SRAM.scala 149:15:@49386.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@49385.4]
  reg  regs_18; // @[SRAM.scala 145:20:@49392.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@49393.4]
  wire  _T_851; // @[SRAM.scala 148:25:@49394.4]
  wire  _T_852; // @[SRAM.scala 148:15:@49395.4]
  wire  _T_853; // @[SRAM.scala 149:15:@49397.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@49396.4]
  reg  regs_19; // @[SRAM.scala 145:20:@49403.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@49404.4]
  wire  _T_860; // @[SRAM.scala 148:25:@49405.4]
  wire  _T_861; // @[SRAM.scala 148:15:@49406.4]
  wire  _T_862; // @[SRAM.scala 149:15:@49408.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@49407.4]
  reg  regs_20; // @[SRAM.scala 145:20:@49414.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@49415.4]
  wire  _T_869; // @[SRAM.scala 148:25:@49416.4]
  wire  _T_870; // @[SRAM.scala 148:15:@49417.4]
  wire  _T_871; // @[SRAM.scala 149:15:@49419.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@49418.4]
  reg  regs_21; // @[SRAM.scala 145:20:@49425.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@49426.4]
  wire  _T_878; // @[SRAM.scala 148:25:@49427.4]
  wire  _T_879; // @[SRAM.scala 148:15:@49428.4]
  wire  _T_880; // @[SRAM.scala 149:15:@49430.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@49429.4]
  reg  regs_22; // @[SRAM.scala 145:20:@49436.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@49437.4]
  wire  _T_887; // @[SRAM.scala 148:25:@49438.4]
  wire  _T_888; // @[SRAM.scala 148:15:@49439.4]
  wire  _T_889; // @[SRAM.scala 149:15:@49441.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@49440.4]
  reg  regs_23; // @[SRAM.scala 145:20:@49447.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@49448.4]
  wire  _T_896; // @[SRAM.scala 148:25:@49449.4]
  wire  _T_897; // @[SRAM.scala 148:15:@49450.4]
  wire  _T_898; // @[SRAM.scala 149:15:@49452.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@49451.4]
  reg  regs_24; // @[SRAM.scala 145:20:@49458.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@49459.4]
  wire  _T_905; // @[SRAM.scala 148:25:@49460.4]
  wire  _T_906; // @[SRAM.scala 148:15:@49461.4]
  wire  _T_907; // @[SRAM.scala 149:15:@49463.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@49462.4]
  reg  regs_25; // @[SRAM.scala 145:20:@49469.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@49470.4]
  wire  _T_914; // @[SRAM.scala 148:25:@49471.4]
  wire  _T_915; // @[SRAM.scala 148:15:@49472.4]
  wire  _T_916; // @[SRAM.scala 149:15:@49474.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@49473.4]
  reg  regs_26; // @[SRAM.scala 145:20:@49480.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@49481.4]
  wire  _T_923; // @[SRAM.scala 148:25:@49482.4]
  wire  _T_924; // @[SRAM.scala 148:15:@49483.4]
  wire  _T_925; // @[SRAM.scala 149:15:@49485.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@49484.4]
  reg  regs_27; // @[SRAM.scala 145:20:@49491.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@49492.4]
  wire  _T_932; // @[SRAM.scala 148:25:@49493.4]
  wire  _T_933; // @[SRAM.scala 148:15:@49494.4]
  wire  _T_934; // @[SRAM.scala 149:15:@49496.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@49495.4]
  reg  regs_28; // @[SRAM.scala 145:20:@49502.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@49503.4]
  wire  _T_941; // @[SRAM.scala 148:25:@49504.4]
  wire  _T_942; // @[SRAM.scala 148:15:@49505.4]
  wire  _T_943; // @[SRAM.scala 149:15:@49507.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@49506.4]
  reg  regs_29; // @[SRAM.scala 145:20:@49513.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@49514.4]
  wire  _T_950; // @[SRAM.scala 148:25:@49515.4]
  wire  _T_951; // @[SRAM.scala 148:15:@49516.4]
  wire  _T_952; // @[SRAM.scala 149:15:@49518.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@49517.4]
  reg  regs_30; // @[SRAM.scala 145:20:@49524.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@49525.4]
  wire  _T_959; // @[SRAM.scala 148:25:@49526.4]
  wire  _T_960; // @[SRAM.scala 148:15:@49527.4]
  wire  _T_961; // @[SRAM.scala 149:15:@49529.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@49528.4]
  reg  regs_31; // @[SRAM.scala 145:20:@49535.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@49536.4]
  wire  _T_968; // @[SRAM.scala 148:25:@49537.4]
  wire  _T_969; // @[SRAM.scala 148:15:@49538.4]
  wire  _T_970; // @[SRAM.scala 149:15:@49540.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@49539.4]
  reg  regs_32; // @[SRAM.scala 145:20:@49546.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@49547.4]
  wire  _T_977; // @[SRAM.scala 148:25:@49548.4]
  wire  _T_978; // @[SRAM.scala 148:15:@49549.4]
  wire  _T_979; // @[SRAM.scala 149:15:@49551.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@49550.4]
  reg  regs_33; // @[SRAM.scala 145:20:@49557.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@49558.4]
  wire  _T_986; // @[SRAM.scala 148:25:@49559.4]
  wire  _T_987; // @[SRAM.scala 148:15:@49560.4]
  wire  _T_988; // @[SRAM.scala 149:15:@49562.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@49561.4]
  reg  regs_34; // @[SRAM.scala 145:20:@49568.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@49569.4]
  wire  _T_995; // @[SRAM.scala 148:25:@49570.4]
  wire  _T_996; // @[SRAM.scala 148:15:@49571.4]
  wire  _T_997; // @[SRAM.scala 149:15:@49573.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@49572.4]
  reg  regs_35; // @[SRAM.scala 145:20:@49579.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@49580.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@49581.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@49582.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@49584.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@49583.4]
  reg  regs_36; // @[SRAM.scala 145:20:@49590.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@49591.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@49592.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@49593.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@49595.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@49594.4]
  reg  regs_37; // @[SRAM.scala 145:20:@49601.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@49602.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@49603.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@49604.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@49606.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@49605.4]
  reg  regs_38; // @[SRAM.scala 145:20:@49612.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@49613.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@49614.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@49615.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@49617.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@49616.4]
  reg  regs_39; // @[SRAM.scala 145:20:@49623.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@49624.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@49625.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@49626.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@49628.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@49627.4]
  reg  regs_40; // @[SRAM.scala 145:20:@49634.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@49635.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@49636.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@49637.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@49639.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@49638.4]
  reg  regs_41; // @[SRAM.scala 145:20:@49645.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@49646.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@49647.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@49648.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@49650.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@49649.4]
  reg  regs_42; // @[SRAM.scala 145:20:@49656.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@49657.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@49658.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@49659.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@49661.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@49660.4]
  reg  regs_43; // @[SRAM.scala 145:20:@49667.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@49668.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@49669.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@49670.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@49672.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@49671.4]
  reg  regs_44; // @[SRAM.scala 145:20:@49678.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@49679.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@49680.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@49681.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@49683.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@49682.4]
  reg  regs_45; // @[SRAM.scala 145:20:@49689.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@49690.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@49691.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@49692.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@49694.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@49693.4]
  reg  regs_46; // @[SRAM.scala 145:20:@49700.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@49701.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@49702.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@49703.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@49705.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@49704.4]
  reg  regs_47; // @[SRAM.scala 145:20:@49711.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@49712.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@49713.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@49714.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@49716.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@49715.4]
  reg  regs_48; // @[SRAM.scala 145:20:@49722.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@49723.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@49724.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@49725.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@49727.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@49726.4]
  reg  regs_49; // @[SRAM.scala 145:20:@49733.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@49734.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@49735.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@49736.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@49738.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@49737.4]
  reg  regs_50; // @[SRAM.scala 145:20:@49744.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@49745.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@49746.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@49747.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@49749.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@49748.4]
  reg  regs_51; // @[SRAM.scala 145:20:@49755.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@49756.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@49757.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@49758.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@49760.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@49759.4]
  reg  regs_52; // @[SRAM.scala 145:20:@49766.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@49767.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@49768.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@49769.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@49771.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@49770.4]
  reg  regs_53; // @[SRAM.scala 145:20:@49777.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@49778.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@49779.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@49780.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@49782.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@49781.4]
  reg  regs_54; // @[SRAM.scala 145:20:@49788.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@49789.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@49790.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@49791.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@49793.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@49792.4]
  reg  regs_55; // @[SRAM.scala 145:20:@49799.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@49800.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@49801.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@49802.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@49804.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@49803.4]
  reg  regs_56; // @[SRAM.scala 145:20:@49810.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@49811.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@49812.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@49813.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@49815.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@49814.4]
  reg  regs_57; // @[SRAM.scala 145:20:@49821.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@49822.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@49823.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@49824.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@49826.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@49825.4]
  reg  regs_58; // @[SRAM.scala 145:20:@49832.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@49833.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@49834.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@49835.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@49837.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@49836.4]
  reg  regs_59; // @[SRAM.scala 145:20:@49843.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@49844.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@49845.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@49846.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@49848.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@49847.4]
  reg  regs_60; // @[SRAM.scala 145:20:@49854.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@49855.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@49856.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@49857.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@49859.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@49858.4]
  reg  regs_61; // @[SRAM.scala 145:20:@49865.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@49866.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@49867.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@49868.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@49870.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@49869.4]
  reg  regs_62; // @[SRAM.scala 145:20:@49876.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@49877.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@49878.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@49879.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@49881.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@49880.4]
  reg  regs_63; // @[SRAM.scala 145:20:@49887.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@49888.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@49889.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@49890.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@49892.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@49891.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@49961.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@49961.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@49195.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@49196.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@49197.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49199.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@49198.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@49206.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@49207.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@49208.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49210.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@49209.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@49217.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@49218.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@49219.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49221.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@49220.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@49228.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@49229.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@49230.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49232.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@49231.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@49239.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@49240.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@49241.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49243.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@49242.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@49250.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@49251.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@49252.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49254.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@49253.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@49261.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@49262.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@49263.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49265.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@49264.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@49272.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@49273.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@49274.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49276.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@49275.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@49283.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@49284.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@49285.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49287.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@49286.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@49294.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@49295.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@49296.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49298.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@49297.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@49305.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@49306.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@49307.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49309.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@49308.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@49316.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@49317.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@49318.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49320.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@49319.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@49327.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@49328.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@49329.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49331.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@49330.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@49338.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@49339.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@49340.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49342.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@49341.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@49349.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@49350.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@49351.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49353.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@49352.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@49360.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@49361.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@49362.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49364.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@49363.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@49371.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@49372.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@49373.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49375.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@49374.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@49382.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@49383.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@49384.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49386.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@49385.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@49393.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@49394.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@49395.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49397.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@49396.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@49404.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@49405.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@49406.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49408.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@49407.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@49415.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@49416.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@49417.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49419.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@49418.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@49426.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@49427.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@49428.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49430.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@49429.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@49437.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@49438.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@49439.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49441.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@49440.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@49448.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@49449.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@49450.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49452.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@49451.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@49459.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@49460.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@49461.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49463.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@49462.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@49470.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@49471.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@49472.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49474.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@49473.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@49481.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@49482.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@49483.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49485.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@49484.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@49492.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@49493.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@49494.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49496.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@49495.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@49503.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@49504.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@49505.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49507.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@49506.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@49514.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@49515.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@49516.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49518.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@49517.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@49525.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@49526.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@49527.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49529.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@49528.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@49536.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@49537.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@49538.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49540.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@49539.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@49547.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@49548.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@49549.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49551.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@49550.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@49558.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@49559.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@49560.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49562.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@49561.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@49569.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@49570.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@49571.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49573.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@49572.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@49580.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@49581.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@49582.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49584.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@49583.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@49591.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@49592.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@49593.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49595.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@49594.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@49602.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@49603.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@49604.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49606.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@49605.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@49613.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@49614.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@49615.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49617.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@49616.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@49624.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@49625.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@49626.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49628.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@49627.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@49635.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@49636.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@49637.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49639.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@49638.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@49646.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@49647.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@49648.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49650.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@49649.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@49657.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@49658.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@49659.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49661.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@49660.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@49668.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@49669.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@49670.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49672.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@49671.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@49679.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@49680.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@49681.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49683.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@49682.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@49690.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@49691.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@49692.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49694.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@49693.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@49701.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@49702.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@49703.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49705.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@49704.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@49712.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@49713.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@49714.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49716.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@49715.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@49723.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@49724.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@49725.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49727.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@49726.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@49734.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@49735.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@49736.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49738.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@49737.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@49745.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@49746.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@49747.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49749.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@49748.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@49756.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@49757.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@49758.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49760.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@49759.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@49767.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@49768.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@49769.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49771.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@49770.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@49778.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@49779.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@49780.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49782.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@49781.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@49789.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@49790.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@49791.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49793.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@49792.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@49800.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@49801.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@49802.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49804.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@49803.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@49811.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@49812.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@49813.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49815.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@49814.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@49822.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@49823.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@49824.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49826.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@49825.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@49833.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@49834.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@49835.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49837.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@49836.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@49844.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@49845.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@49846.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49848.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@49847.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@49855.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@49856.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@49857.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49859.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@49858.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@49866.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@49867.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@49868.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49870.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@49869.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@49877.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@49878.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@49879.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49881.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@49880.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@49888.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@49889.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@49890.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@49892.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@49891.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@49961.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@49961.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@49961.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@49963.2]
  input   clock, // @[:@49964.4]
  input   reset, // @[:@49965.4]
  output  io_in_ready, // @[:@49966.4]
  input   io_in_valid, // @[:@49966.4]
  input   io_in_bits, // @[:@49966.4]
  input   io_out_ready, // @[:@49966.4]
  output  io_out_valid, // @[:@49966.4]
  output  io_out_bits, // @[:@49966.4]
  input   io_banks_0_wdata_valid, // @[:@49966.4]
  input   io_banks_0_wdata_bits, // @[:@49966.4]
  input   io_banks_1_wdata_valid, // @[:@49966.4]
  input   io_banks_1_wdata_bits, // @[:@49966.4]
  input   io_banks_2_wdata_valid, // @[:@49966.4]
  input   io_banks_2_wdata_bits, // @[:@49966.4]
  input   io_banks_3_wdata_valid, // @[:@49966.4]
  input   io_banks_3_wdata_bits, // @[:@49966.4]
  input   io_banks_4_wdata_valid, // @[:@49966.4]
  input   io_banks_4_wdata_bits, // @[:@49966.4]
  input   io_banks_5_wdata_valid, // @[:@49966.4]
  input   io_banks_5_wdata_bits, // @[:@49966.4]
  input   io_banks_6_wdata_valid, // @[:@49966.4]
  input   io_banks_6_wdata_bits, // @[:@49966.4]
  input   io_banks_7_wdata_valid, // @[:@49966.4]
  input   io_banks_7_wdata_bits, // @[:@49966.4]
  input   io_banks_8_wdata_valid, // @[:@49966.4]
  input   io_banks_8_wdata_bits, // @[:@49966.4]
  input   io_banks_9_wdata_valid, // @[:@49966.4]
  input   io_banks_9_wdata_bits, // @[:@49966.4]
  input   io_banks_10_wdata_valid, // @[:@49966.4]
  input   io_banks_10_wdata_bits, // @[:@49966.4]
  input   io_banks_11_wdata_valid, // @[:@49966.4]
  input   io_banks_11_wdata_bits, // @[:@49966.4]
  input   io_banks_12_wdata_valid, // @[:@49966.4]
  input   io_banks_12_wdata_bits, // @[:@49966.4]
  input   io_banks_13_wdata_valid, // @[:@49966.4]
  input   io_banks_13_wdata_bits, // @[:@49966.4]
  input   io_banks_14_wdata_valid, // @[:@49966.4]
  input   io_banks_14_wdata_bits, // @[:@49966.4]
  input   io_banks_15_wdata_valid, // @[:@49966.4]
  input   io_banks_15_wdata_bits, // @[:@49966.4]
  input   io_banks_16_wdata_valid, // @[:@49966.4]
  input   io_banks_16_wdata_bits, // @[:@49966.4]
  input   io_banks_17_wdata_valid, // @[:@49966.4]
  input   io_banks_17_wdata_bits, // @[:@49966.4]
  input   io_banks_18_wdata_valid, // @[:@49966.4]
  input   io_banks_18_wdata_bits, // @[:@49966.4]
  input   io_banks_19_wdata_valid, // @[:@49966.4]
  input   io_banks_19_wdata_bits, // @[:@49966.4]
  input   io_banks_20_wdata_valid, // @[:@49966.4]
  input   io_banks_20_wdata_bits, // @[:@49966.4]
  input   io_banks_21_wdata_valid, // @[:@49966.4]
  input   io_banks_21_wdata_bits, // @[:@49966.4]
  input   io_banks_22_wdata_valid, // @[:@49966.4]
  input   io_banks_22_wdata_bits, // @[:@49966.4]
  input   io_banks_23_wdata_valid, // @[:@49966.4]
  input   io_banks_23_wdata_bits, // @[:@49966.4]
  input   io_banks_24_wdata_valid, // @[:@49966.4]
  input   io_banks_24_wdata_bits, // @[:@49966.4]
  input   io_banks_25_wdata_valid, // @[:@49966.4]
  input   io_banks_25_wdata_bits, // @[:@49966.4]
  input   io_banks_26_wdata_valid, // @[:@49966.4]
  input   io_banks_26_wdata_bits, // @[:@49966.4]
  input   io_banks_27_wdata_valid, // @[:@49966.4]
  input   io_banks_27_wdata_bits, // @[:@49966.4]
  input   io_banks_28_wdata_valid, // @[:@49966.4]
  input   io_banks_28_wdata_bits, // @[:@49966.4]
  input   io_banks_29_wdata_valid, // @[:@49966.4]
  input   io_banks_29_wdata_bits, // @[:@49966.4]
  input   io_banks_30_wdata_valid, // @[:@49966.4]
  input   io_banks_30_wdata_bits, // @[:@49966.4]
  input   io_banks_31_wdata_valid, // @[:@49966.4]
  input   io_banks_31_wdata_bits, // @[:@49966.4]
  input   io_banks_32_wdata_valid, // @[:@49966.4]
  input   io_banks_32_wdata_bits, // @[:@49966.4]
  input   io_banks_33_wdata_valid, // @[:@49966.4]
  input   io_banks_33_wdata_bits, // @[:@49966.4]
  input   io_banks_34_wdata_valid, // @[:@49966.4]
  input   io_banks_34_wdata_bits, // @[:@49966.4]
  input   io_banks_35_wdata_valid, // @[:@49966.4]
  input   io_banks_35_wdata_bits, // @[:@49966.4]
  input   io_banks_36_wdata_valid, // @[:@49966.4]
  input   io_banks_36_wdata_bits, // @[:@49966.4]
  input   io_banks_37_wdata_valid, // @[:@49966.4]
  input   io_banks_37_wdata_bits, // @[:@49966.4]
  input   io_banks_38_wdata_valid, // @[:@49966.4]
  input   io_banks_38_wdata_bits, // @[:@49966.4]
  input   io_banks_39_wdata_valid, // @[:@49966.4]
  input   io_banks_39_wdata_bits, // @[:@49966.4]
  input   io_banks_40_wdata_valid, // @[:@49966.4]
  input   io_banks_40_wdata_bits, // @[:@49966.4]
  input   io_banks_41_wdata_valid, // @[:@49966.4]
  input   io_banks_41_wdata_bits, // @[:@49966.4]
  input   io_banks_42_wdata_valid, // @[:@49966.4]
  input   io_banks_42_wdata_bits, // @[:@49966.4]
  input   io_banks_43_wdata_valid, // @[:@49966.4]
  input   io_banks_43_wdata_bits, // @[:@49966.4]
  input   io_banks_44_wdata_valid, // @[:@49966.4]
  input   io_banks_44_wdata_bits, // @[:@49966.4]
  input   io_banks_45_wdata_valid, // @[:@49966.4]
  input   io_banks_45_wdata_bits, // @[:@49966.4]
  input   io_banks_46_wdata_valid, // @[:@49966.4]
  input   io_banks_46_wdata_bits, // @[:@49966.4]
  input   io_banks_47_wdata_valid, // @[:@49966.4]
  input   io_banks_47_wdata_bits, // @[:@49966.4]
  input   io_banks_48_wdata_valid, // @[:@49966.4]
  input   io_banks_48_wdata_bits, // @[:@49966.4]
  input   io_banks_49_wdata_valid, // @[:@49966.4]
  input   io_banks_49_wdata_bits, // @[:@49966.4]
  input   io_banks_50_wdata_valid, // @[:@49966.4]
  input   io_banks_50_wdata_bits, // @[:@49966.4]
  input   io_banks_51_wdata_valid, // @[:@49966.4]
  input   io_banks_51_wdata_bits, // @[:@49966.4]
  input   io_banks_52_wdata_valid, // @[:@49966.4]
  input   io_banks_52_wdata_bits, // @[:@49966.4]
  input   io_banks_53_wdata_valid, // @[:@49966.4]
  input   io_banks_53_wdata_bits, // @[:@49966.4]
  input   io_banks_54_wdata_valid, // @[:@49966.4]
  input   io_banks_54_wdata_bits, // @[:@49966.4]
  input   io_banks_55_wdata_valid, // @[:@49966.4]
  input   io_banks_55_wdata_bits, // @[:@49966.4]
  input   io_banks_56_wdata_valid, // @[:@49966.4]
  input   io_banks_56_wdata_bits, // @[:@49966.4]
  input   io_banks_57_wdata_valid, // @[:@49966.4]
  input   io_banks_57_wdata_bits, // @[:@49966.4]
  input   io_banks_58_wdata_valid, // @[:@49966.4]
  input   io_banks_58_wdata_bits, // @[:@49966.4]
  input   io_banks_59_wdata_valid, // @[:@49966.4]
  input   io_banks_59_wdata_bits, // @[:@49966.4]
  input   io_banks_60_wdata_valid, // @[:@49966.4]
  input   io_banks_60_wdata_bits, // @[:@49966.4]
  input   io_banks_61_wdata_valid, // @[:@49966.4]
  input   io_banks_61_wdata_bits, // @[:@49966.4]
  input   io_banks_62_wdata_valid, // @[:@49966.4]
  input   io_banks_62_wdata_bits, // @[:@49966.4]
  input   io_banks_63_wdata_valid, // @[:@49966.4]
  input   io_banks_63_wdata_bits // @[:@49966.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@50232.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@50232.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@50232.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@50232.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@50232.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@50242.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@50242.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@50242.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@50242.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@50242.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@50257.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@50257.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@50257.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@50257.4]
  wire  writeEn; // @[FIFO.scala 30:29:@50230.4]
  wire  readEn; // @[FIFO.scala 31:29:@50231.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@50252.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@50253.4]
  wire  _T_824; // @[FIFO.scala 45:27:@50254.4]
  wire  empty; // @[FIFO.scala 45:24:@50255.4]
  wire  full; // @[FIFO.scala 46:23:@50256.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@51423.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@51424.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@50232.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@50242.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@50257.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@50230.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@50231.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@50253.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@50254.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@50255.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@50256.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@51423.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@51424.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@51430.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@51428.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@50462.4]
  assign enqCounter_clock = clock; // @[:@50233.4]
  assign enqCounter_reset = reset; // @[:@50234.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@50240.4]
  assign deqCounter_clock = clock; // @[:@50243.4]
  assign deqCounter_reset = reset; // @[:@50244.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@50250.4]
  assign FFRAM_clock = clock; // @[:@50258.4]
  assign FFRAM_reset = reset; // @[:@50259.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@50458.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@50459.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@50460.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@50461.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@50464.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@50463.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@50467.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@50466.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@50470.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@50469.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@50473.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@50472.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@50476.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@50475.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@50479.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@50478.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@50482.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@50481.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@50485.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@50484.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@50488.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@50487.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@50491.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@50490.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@50494.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@50493.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@50497.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@50496.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@50500.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@50499.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@50503.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@50502.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@50506.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@50505.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@50509.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@50508.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@50512.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@50511.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@50515.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@50514.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@50518.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@50517.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@50521.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@50520.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@50524.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@50523.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@50527.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@50526.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@50530.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@50529.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@50533.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@50532.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@50536.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@50535.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@50539.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@50538.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@50542.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@50541.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@50545.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@50544.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@50548.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@50547.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@50551.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@50550.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@50554.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@50553.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@50557.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@50556.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@50560.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@50559.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@50563.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@50562.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@50566.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@50565.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@50569.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@50568.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@50572.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@50571.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@50575.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@50574.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@50578.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@50577.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@50581.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@50580.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@50584.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@50583.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@50587.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@50586.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@50590.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@50589.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@50593.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@50592.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@50596.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@50595.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@50599.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@50598.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@50602.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@50601.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@50605.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@50604.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@50608.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@50607.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@50611.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@50610.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@50614.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@50613.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@50617.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@50616.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@50620.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@50619.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@50623.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@50622.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@50626.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@50625.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@50629.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@50628.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@50632.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@50631.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@50635.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@50634.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@50638.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@50637.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@50641.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@50640.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@50644.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@50643.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@50647.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@50646.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@50650.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@50649.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@50653.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@50652.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@51432.2]
  input         clock, // @[:@51433.4]
  input         reset, // @[:@51434.4]
  input         io_dram_cmd_ready, // @[:@51435.4]
  output        io_dram_cmd_valid, // @[:@51435.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@51435.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@51435.4]
  input         io_dram_wdata_ready, // @[:@51435.4]
  output        io_dram_wdata_valid, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@51435.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@51435.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@51435.4]
  output        io_dram_wresp_ready, // @[:@51435.4]
  input         io_dram_wresp_valid, // @[:@51435.4]
  output        io_store_cmd_ready, // @[:@51435.4]
  input         io_store_cmd_valid, // @[:@51435.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@51435.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@51435.4]
  output        io_store_data_ready, // @[:@51435.4]
  input         io_store_data_valid, // @[:@51435.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@51435.4]
  input         io_store_data_bits_wstrb, // @[:@51435.4]
  input         io_store_wresp_ready, // @[:@51435.4]
  output        io_store_wresp_valid, // @[:@51435.4]
  output        io_store_wresp_bits // @[:@51435.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@51560.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@51560.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@51560.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@51560.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@51560.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@51560.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@51560.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@51560.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@51560.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@51560.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@51966.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@51966.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@51966.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@51966.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@51966.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@51966.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@51966.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@51966.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@51966.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@52207.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@52207.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@51963.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@51560.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@51966.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@52207.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@51963.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@51960.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@51961.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@51964.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@51996.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@51997.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@51998.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@51999.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@52000.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@52001.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@52002.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@52003.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@52004.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@52005.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@52006.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@52007.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@52008.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@52009.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@52010.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@52011.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@52012.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@52142.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@52143.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@52144.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@52145.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@52146.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@52147.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@52148.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@52149.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@52150.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@52151.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@52152.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@52153.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@52154.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@52155.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@52156.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@52157.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@52158.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@52159.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@52160.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@52161.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@52162.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@52163.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@52164.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@52165.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@52166.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@52167.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@52168.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@52169.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@52170.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@52171.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@52172.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@52173.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@52174.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@52175.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@52176.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@52177.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@52178.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@52179.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@52180.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@52181.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@52182.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@52183.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@52184.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@52185.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@52186.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@52187.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@52188.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@52189.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@52190.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@52191.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@52192.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@52193.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@52194.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@52195.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@52196.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@52197.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@52198.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@52199.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@52200.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@52201.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@52202.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@52203.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@52204.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@52205.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@52474.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@51958.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@51995.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@52475.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@52476.4]
  assign cmd_clock = clock; // @[:@51561.4]
  assign cmd_reset = reset; // @[:@51562.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@51955.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@51957.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@51956.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@51959.4]
  assign wdata_clock = clock; // @[:@51967.4]
  assign wdata_reset = reset; // @[:@51968.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@51992.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@51993.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@51994.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@52206.4]
  assign wresp_clock = clock; // @[:@52208.4]
  assign wresp_reset = reset; // @[:@52209.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@52472.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@52473.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@52477.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@52543.2]
  output        io_in_ready, // @[:@52546.4]
  input         io_in_valid, // @[:@52546.4]
  input  [63:0] io_in_bits_0_addr, // @[:@52546.4]
  input  [31:0] io_in_bits_0_size, // @[:@52546.4]
  input         io_in_bits_0_isWr, // @[:@52546.4]
  input  [31:0] io_in_bits_0_tag, // @[:@52546.4]
  input         io_out_ready, // @[:@52546.4]
  output        io_out_valid, // @[:@52546.4]
  output [63:0] io_out_bits_addr, // @[:@52546.4]
  output [31:0] io_out_bits_size, // @[:@52546.4]
  output        io_out_bits_isWr, // @[:@52546.4]
  output [31:0] io_out_bits_tag // @[:@52546.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@52548.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@52548.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@52557.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@52556.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@52562.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@52561.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@52559.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@52558.4]
endmodule
module MuxPipe_1( // @[:@52564.2]
  output        io_in_ready, // @[:@52567.4]
  input         io_in_valid, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@52567.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@52567.4]
  input         io_in_bits_0_wstrb_0, // @[:@52567.4]
  input         io_in_bits_0_wstrb_1, // @[:@52567.4]
  input         io_in_bits_0_wstrb_2, // @[:@52567.4]
  input         io_in_bits_0_wstrb_3, // @[:@52567.4]
  input         io_in_bits_0_wstrb_4, // @[:@52567.4]
  input         io_in_bits_0_wstrb_5, // @[:@52567.4]
  input         io_in_bits_0_wstrb_6, // @[:@52567.4]
  input         io_in_bits_0_wstrb_7, // @[:@52567.4]
  input         io_in_bits_0_wstrb_8, // @[:@52567.4]
  input         io_in_bits_0_wstrb_9, // @[:@52567.4]
  input         io_in_bits_0_wstrb_10, // @[:@52567.4]
  input         io_in_bits_0_wstrb_11, // @[:@52567.4]
  input         io_in_bits_0_wstrb_12, // @[:@52567.4]
  input         io_in_bits_0_wstrb_13, // @[:@52567.4]
  input         io_in_bits_0_wstrb_14, // @[:@52567.4]
  input         io_in_bits_0_wstrb_15, // @[:@52567.4]
  input         io_in_bits_0_wstrb_16, // @[:@52567.4]
  input         io_in_bits_0_wstrb_17, // @[:@52567.4]
  input         io_in_bits_0_wstrb_18, // @[:@52567.4]
  input         io_in_bits_0_wstrb_19, // @[:@52567.4]
  input         io_in_bits_0_wstrb_20, // @[:@52567.4]
  input         io_in_bits_0_wstrb_21, // @[:@52567.4]
  input         io_in_bits_0_wstrb_22, // @[:@52567.4]
  input         io_in_bits_0_wstrb_23, // @[:@52567.4]
  input         io_in_bits_0_wstrb_24, // @[:@52567.4]
  input         io_in_bits_0_wstrb_25, // @[:@52567.4]
  input         io_in_bits_0_wstrb_26, // @[:@52567.4]
  input         io_in_bits_0_wstrb_27, // @[:@52567.4]
  input         io_in_bits_0_wstrb_28, // @[:@52567.4]
  input         io_in_bits_0_wstrb_29, // @[:@52567.4]
  input         io_in_bits_0_wstrb_30, // @[:@52567.4]
  input         io_in_bits_0_wstrb_31, // @[:@52567.4]
  input         io_in_bits_0_wstrb_32, // @[:@52567.4]
  input         io_in_bits_0_wstrb_33, // @[:@52567.4]
  input         io_in_bits_0_wstrb_34, // @[:@52567.4]
  input         io_in_bits_0_wstrb_35, // @[:@52567.4]
  input         io_in_bits_0_wstrb_36, // @[:@52567.4]
  input         io_in_bits_0_wstrb_37, // @[:@52567.4]
  input         io_in_bits_0_wstrb_38, // @[:@52567.4]
  input         io_in_bits_0_wstrb_39, // @[:@52567.4]
  input         io_in_bits_0_wstrb_40, // @[:@52567.4]
  input         io_in_bits_0_wstrb_41, // @[:@52567.4]
  input         io_in_bits_0_wstrb_42, // @[:@52567.4]
  input         io_in_bits_0_wstrb_43, // @[:@52567.4]
  input         io_in_bits_0_wstrb_44, // @[:@52567.4]
  input         io_in_bits_0_wstrb_45, // @[:@52567.4]
  input         io_in_bits_0_wstrb_46, // @[:@52567.4]
  input         io_in_bits_0_wstrb_47, // @[:@52567.4]
  input         io_in_bits_0_wstrb_48, // @[:@52567.4]
  input         io_in_bits_0_wstrb_49, // @[:@52567.4]
  input         io_in_bits_0_wstrb_50, // @[:@52567.4]
  input         io_in_bits_0_wstrb_51, // @[:@52567.4]
  input         io_in_bits_0_wstrb_52, // @[:@52567.4]
  input         io_in_bits_0_wstrb_53, // @[:@52567.4]
  input         io_in_bits_0_wstrb_54, // @[:@52567.4]
  input         io_in_bits_0_wstrb_55, // @[:@52567.4]
  input         io_in_bits_0_wstrb_56, // @[:@52567.4]
  input         io_in_bits_0_wstrb_57, // @[:@52567.4]
  input         io_in_bits_0_wstrb_58, // @[:@52567.4]
  input         io_in_bits_0_wstrb_59, // @[:@52567.4]
  input         io_in_bits_0_wstrb_60, // @[:@52567.4]
  input         io_in_bits_0_wstrb_61, // @[:@52567.4]
  input         io_in_bits_0_wstrb_62, // @[:@52567.4]
  input         io_in_bits_0_wstrb_63, // @[:@52567.4]
  input         io_out_ready, // @[:@52567.4]
  output        io_out_valid, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_0, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_1, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_2, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_3, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_4, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_5, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_6, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_7, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_8, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_9, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_10, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_11, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_12, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_13, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_14, // @[:@52567.4]
  output [31:0] io_out_bits_wdata_15, // @[:@52567.4]
  output        io_out_bits_wstrb_0, // @[:@52567.4]
  output        io_out_bits_wstrb_1, // @[:@52567.4]
  output        io_out_bits_wstrb_2, // @[:@52567.4]
  output        io_out_bits_wstrb_3, // @[:@52567.4]
  output        io_out_bits_wstrb_4, // @[:@52567.4]
  output        io_out_bits_wstrb_5, // @[:@52567.4]
  output        io_out_bits_wstrb_6, // @[:@52567.4]
  output        io_out_bits_wstrb_7, // @[:@52567.4]
  output        io_out_bits_wstrb_8, // @[:@52567.4]
  output        io_out_bits_wstrb_9, // @[:@52567.4]
  output        io_out_bits_wstrb_10, // @[:@52567.4]
  output        io_out_bits_wstrb_11, // @[:@52567.4]
  output        io_out_bits_wstrb_12, // @[:@52567.4]
  output        io_out_bits_wstrb_13, // @[:@52567.4]
  output        io_out_bits_wstrb_14, // @[:@52567.4]
  output        io_out_bits_wstrb_15, // @[:@52567.4]
  output        io_out_bits_wstrb_16, // @[:@52567.4]
  output        io_out_bits_wstrb_17, // @[:@52567.4]
  output        io_out_bits_wstrb_18, // @[:@52567.4]
  output        io_out_bits_wstrb_19, // @[:@52567.4]
  output        io_out_bits_wstrb_20, // @[:@52567.4]
  output        io_out_bits_wstrb_21, // @[:@52567.4]
  output        io_out_bits_wstrb_22, // @[:@52567.4]
  output        io_out_bits_wstrb_23, // @[:@52567.4]
  output        io_out_bits_wstrb_24, // @[:@52567.4]
  output        io_out_bits_wstrb_25, // @[:@52567.4]
  output        io_out_bits_wstrb_26, // @[:@52567.4]
  output        io_out_bits_wstrb_27, // @[:@52567.4]
  output        io_out_bits_wstrb_28, // @[:@52567.4]
  output        io_out_bits_wstrb_29, // @[:@52567.4]
  output        io_out_bits_wstrb_30, // @[:@52567.4]
  output        io_out_bits_wstrb_31, // @[:@52567.4]
  output        io_out_bits_wstrb_32, // @[:@52567.4]
  output        io_out_bits_wstrb_33, // @[:@52567.4]
  output        io_out_bits_wstrb_34, // @[:@52567.4]
  output        io_out_bits_wstrb_35, // @[:@52567.4]
  output        io_out_bits_wstrb_36, // @[:@52567.4]
  output        io_out_bits_wstrb_37, // @[:@52567.4]
  output        io_out_bits_wstrb_38, // @[:@52567.4]
  output        io_out_bits_wstrb_39, // @[:@52567.4]
  output        io_out_bits_wstrb_40, // @[:@52567.4]
  output        io_out_bits_wstrb_41, // @[:@52567.4]
  output        io_out_bits_wstrb_42, // @[:@52567.4]
  output        io_out_bits_wstrb_43, // @[:@52567.4]
  output        io_out_bits_wstrb_44, // @[:@52567.4]
  output        io_out_bits_wstrb_45, // @[:@52567.4]
  output        io_out_bits_wstrb_46, // @[:@52567.4]
  output        io_out_bits_wstrb_47, // @[:@52567.4]
  output        io_out_bits_wstrb_48, // @[:@52567.4]
  output        io_out_bits_wstrb_49, // @[:@52567.4]
  output        io_out_bits_wstrb_50, // @[:@52567.4]
  output        io_out_bits_wstrb_51, // @[:@52567.4]
  output        io_out_bits_wstrb_52, // @[:@52567.4]
  output        io_out_bits_wstrb_53, // @[:@52567.4]
  output        io_out_bits_wstrb_54, // @[:@52567.4]
  output        io_out_bits_wstrb_55, // @[:@52567.4]
  output        io_out_bits_wstrb_56, // @[:@52567.4]
  output        io_out_bits_wstrb_57, // @[:@52567.4]
  output        io_out_bits_wstrb_58, // @[:@52567.4]
  output        io_out_bits_wstrb_59, // @[:@52567.4]
  output        io_out_bits_wstrb_60, // @[:@52567.4]
  output        io_out_bits_wstrb_61, // @[:@52567.4]
  output        io_out_bits_wstrb_62, // @[:@52567.4]
  output        io_out_bits_wstrb_63 // @[:@52567.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@52569.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@52569.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@52654.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@52653.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@52720.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@52721.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@52722.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@52723.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@52724.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@52725.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@52726.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@52727.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@52728.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@52729.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@52730.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@52731.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@52732.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@52733.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@52734.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@52735.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@52656.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@52657.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@52658.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@52659.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@52660.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@52661.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@52662.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@52663.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@52664.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@52665.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@52666.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@52667.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@52668.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@52669.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@52670.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@52671.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@52672.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@52673.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@52674.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@52675.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@52676.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@52677.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@52678.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@52679.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@52680.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@52681.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@52682.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@52683.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@52684.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@52685.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@52686.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@52687.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@52688.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@52689.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@52690.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@52691.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@52692.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@52693.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@52694.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@52695.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@52696.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@52697.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@52698.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@52699.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@52700.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@52701.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@52702.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@52703.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@52704.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@52705.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@52706.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@52707.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@52708.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@52709.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@52710.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@52711.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@52712.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@52713.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@52714.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@52715.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@52716.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@52717.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@52718.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@52719.4]
endmodule
module ElementCounter( // @[:@52737.2]
  input         clock, // @[:@52738.4]
  input         reset, // @[:@52739.4]
  input         io_reset, // @[:@52740.4]
  input         io_enable, // @[:@52740.4]
  output [31:0] io_out // @[:@52740.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@52742.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@52743.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@52744.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@52749.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@52745.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@52743.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@52744.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@52749.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@52745.4]
  assign io_out = count; // @[Counter.scala 47:10:@52752.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@52754.2]
  input         clock, // @[:@52755.4]
  input         reset, // @[:@52756.4]
  output        io_app_0_cmd_ready, // @[:@52757.4]
  input         io_app_0_cmd_valid, // @[:@52757.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@52757.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@52757.4]
  input         io_app_0_cmd_bits_isWr, // @[:@52757.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@52757.4]
  output        io_app_0_wdata_ready, // @[:@52757.4]
  input         io_app_0_wdata_valid, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@52757.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@52757.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@52757.4]
  input         io_app_0_rresp_ready, // @[:@52757.4]
  input         io_app_0_wresp_ready, // @[:@52757.4]
  output        io_app_0_wresp_valid, // @[:@52757.4]
  input         io_dram_cmd_ready, // @[:@52757.4]
  output        io_dram_cmd_valid, // @[:@52757.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@52757.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@52757.4]
  output        io_dram_cmd_bits_isWr, // @[:@52757.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@52757.4]
  input         io_dram_wdata_ready, // @[:@52757.4]
  output        io_dram_wdata_valid, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@52757.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@52757.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@52757.4]
  output        io_dram_rresp_ready, // @[:@52757.4]
  output        io_dram_wresp_ready, // @[:@52757.4]
  input         io_dram_wresp_valid, // @[:@52757.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@52757.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@52986.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@52986.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@52986.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@52986.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@52986.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@52993.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@52993.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@52993.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@52993.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@52993.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@53003.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@53003.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@53003.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@53003.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@53003.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@53003.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@53003.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@53003.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@53003.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@53003.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@53003.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@53003.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@53026.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@53026.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@53029.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@53029.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@53029.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@53029.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@53029.4]
  wire  _T_346; // @[package.scala 96:25:@52998.4 package.scala 96:25:@52999.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@53000.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@53002.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@53018.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@53020.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@53023.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@53032.4]
  wire [31:0] _T_365; // @[:@53036.4 :@53037.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@53038.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@53044.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@53047.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@53048.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@53235.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@53242.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@53247.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@53251.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@53252.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@53276.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@52986.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@52993.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@53003.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@53026.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@53029.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@52998.4 package.scala 96:25:@52999.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@53000.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@53002.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@53018.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@53020.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@53023.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@53032.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@53036.4 :@53037.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@53038.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@53044.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@53047.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@53048.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@53235.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@53242.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@53247.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@53251.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@53252.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@53276.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@53249.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@53255.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@53278.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@53138.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@53137.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@53136.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@53134.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@53133.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@53221.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@53205.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@53206.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@53207.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@53208.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@53209.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@53210.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@53211.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@53212.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@53213.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@53214.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@53215.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@53216.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@53217.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@53218.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@53219.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@53220.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@53141.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@53142.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@53143.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@53144.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@53145.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@53146.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@53147.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@53148.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@53149.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@53150.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@53151.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@53152.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@53153.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@53154.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@53155.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@53156.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@53157.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@53158.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@53159.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@53160.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@53161.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@53162.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@53163.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@53164.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@53165.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@53166.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@53167.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@53168.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@53169.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@53170.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@53171.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@53172.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@53173.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@53174.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@53175.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@53176.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@53177.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@53178.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@53179.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@53180.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@53181.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@53182.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@53183.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@53184.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@53185.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@53186.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@53187.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@53188.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@53189.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@53190.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@53191.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@53192.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@53193.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@53194.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@53195.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@53196.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@53197.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@53198.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@53199.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@53200.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@53201.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@53202.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@53203.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@53204.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@53282.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@53285.4]
  assign RetimeWrapper_clock = clock; // @[:@52987.4]
  assign RetimeWrapper_reset = reset; // @[:@52988.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@52990.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@52989.4]
  assign RetimeWrapper_1_clock = clock; // @[:@52994.4]
  assign RetimeWrapper_1_reset = reset; // @[:@52995.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@52997.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@52996.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@53006.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@53012.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@53011.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@53009.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@53008.4 FringeBundles.scala 115:32:@53025.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@53139.4 StreamArbiter.scala 57:23:@53245.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@53050.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@53117.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@53118.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@53119.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@53120.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@53121.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@53122.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@53123.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@53124.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@53125.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@53126.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@53127.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@53128.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@53129.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@53130.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@53131.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@53132.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@53053.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@53054.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@53055.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@53056.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@53057.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@53058.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@53059.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@53060.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@53061.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@53062.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@53063.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@53064.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@53065.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@53066.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@53067.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@53068.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@53069.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@53070.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@53071.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@53072.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@53073.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@53074.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@53075.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@53076.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@53077.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@53078.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@53079.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@53080.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@53081.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@53082.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@53083.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@53084.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@53085.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@53086.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@53087.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@53088.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@53089.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@53090.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@53091.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@53092.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@53093.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@53094.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@53095.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@53096.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@53097.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@53098.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@53099.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@53100.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@53101.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@53102.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@53103.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@53104.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@53105.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@53106.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@53107.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@53108.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@53109.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@53110.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@53111.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@53112.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@53113.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@53114.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@53115.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@53116.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@53222.4 StreamArbiter.scala 58:25:@53246.4]
  assign elementCtr_clock = clock; // @[:@53030.4]
  assign elementCtr_reset = reset; // @[:@53031.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@53034.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@53033.4]
endmodule
module Counter_72( // @[:@53287.2]
  input         clock, // @[:@53288.4]
  input         reset, // @[:@53289.4]
  input         io_reset, // @[:@53290.4]
  input         io_enable, // @[:@53290.4]
  input  [31:0] io_stride, // @[:@53290.4]
  output [31:0] io_out, // @[:@53290.4]
  output [31:0] io_next // @[:@53290.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@53292.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@53293.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@53294.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@53299.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@53295.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@53293.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@53294.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@53299.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@53295.4]
  assign io_out = count; // @[Counter.scala 25:10:@53302.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@53303.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@53305.2]
  input         clock, // @[:@53306.4]
  input         reset, // @[:@53307.4]
  output        io_in_cmd_ready, // @[:@53308.4]
  input         io_in_cmd_valid, // @[:@53308.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@53308.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@53308.4]
  input         io_in_cmd_bits_isWr, // @[:@53308.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@53308.4]
  output        io_in_wdata_ready, // @[:@53308.4]
  input         io_in_wdata_valid, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@53308.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@53308.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@53308.4]
  input         io_in_rresp_ready, // @[:@53308.4]
  input         io_in_wresp_ready, // @[:@53308.4]
  output        io_in_wresp_valid, // @[:@53308.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@53308.4]
  input         io_out_cmd_ready, // @[:@53308.4]
  output        io_out_cmd_valid, // @[:@53308.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@53308.4]
  output [31:0] io_out_cmd_bits_size, // @[:@53308.4]
  output        io_out_cmd_bits_isWr, // @[:@53308.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@53308.4]
  input         io_out_wdata_ready, // @[:@53308.4]
  output        io_out_wdata_valid, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@53308.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@53308.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@53308.4]
  output        io_out_rresp_ready, // @[:@53308.4]
  output        io_out_wresp_ready, // @[:@53308.4]
  input         io_out_wresp_valid, // @[:@53308.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@53308.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@53422.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@53422.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@53422.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@53422.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@53422.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@53422.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@53422.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@53425.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@53426.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@53427.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@53428.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@53431.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@53431.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@53432.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@53432.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@53433.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@53436.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@53443.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@53447.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@53450.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@53453.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@53464.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@53422.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@53425.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@53426.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@53427.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@53428.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@53431.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@53431.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@53432.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@53432.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@53433.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@53436.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@53443.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@53447.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@53450.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@53453.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@53464.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@53421.4 AXIProtocol.scala 38:19:@53455.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@53414.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@53311.4 AXIProtocol.scala 46:21:@53469.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@53310.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@53420.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@53419.4 AXIProtocol.scala 29:24:@53438.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@53418.4 AXIProtocol.scala 25:24:@53430.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@53416.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@53415.4 FringeBundles.scala 115:32:@53452.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@53413.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@53397.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@53398.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@53399.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@53400.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@53401.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@53402.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@53403.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@53404.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@53405.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@53406.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@53407.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@53408.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@53409.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@53410.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@53411.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@53412.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@53333.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@53334.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@53335.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@53336.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@53337.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@53338.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@53339.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@53340.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@53341.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@53342.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@53343.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@53344.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@53345.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@53346.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@53347.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@53348.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@53349.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@53350.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@53351.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@53352.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@53353.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@53354.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@53355.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@53356.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@53357.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@53358.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@53359.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@53360.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@53361.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@53362.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@53363.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@53364.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@53365.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@53366.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@53367.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@53368.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@53369.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@53370.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@53371.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@53372.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@53373.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@53374.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@53375.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@53376.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@53377.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@53378.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@53379.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@53380.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@53381.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@53382.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@53383.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@53384.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@53385.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@53386.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@53387.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@53388.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@53389.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@53390.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@53391.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@53392.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@53393.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@53394.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@53395.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@53396.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@53331.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@53312.4 AXIProtocol.scala 47:22:@53471.4]
  assign cmdSizeCounter_clock = clock; // @[:@53423.4]
  assign cmdSizeCounter_reset = reset; // @[:@53424.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@53456.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@53457.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@53458.4]
endmodule
module AXICmdIssue( // @[:@53491.2]
  input         clock, // @[:@53492.4]
  input         reset, // @[:@53493.4]
  output        io_in_cmd_ready, // @[:@53494.4]
  input         io_in_cmd_valid, // @[:@53494.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@53494.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@53494.4]
  input         io_in_cmd_bits_isWr, // @[:@53494.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@53494.4]
  output        io_in_wdata_ready, // @[:@53494.4]
  input         io_in_wdata_valid, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@53494.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@53494.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@53494.4]
  input         io_in_rresp_ready, // @[:@53494.4]
  input         io_in_wresp_ready, // @[:@53494.4]
  output        io_in_wresp_valid, // @[:@53494.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@53494.4]
  input         io_out_cmd_ready, // @[:@53494.4]
  output        io_out_cmd_valid, // @[:@53494.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@53494.4]
  output [31:0] io_out_cmd_bits_size, // @[:@53494.4]
  output        io_out_cmd_bits_isWr, // @[:@53494.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@53494.4]
  input         io_out_wdata_ready, // @[:@53494.4]
  output        io_out_wdata_valid, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@53494.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@53494.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@53494.4]
  output        io_out_wdata_bits_wlast, // @[:@53494.4]
  output        io_out_rresp_ready, // @[:@53494.4]
  output        io_out_wresp_ready, // @[:@53494.4]
  input         io_out_wresp_valid, // @[:@53494.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@53494.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@53608.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@53608.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@53608.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@53608.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@53608.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@53608.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@53608.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@53611.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@53612.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@53613.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@53614.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@53615.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@53621.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@53622.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@53617.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@53631.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@53632.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@53608.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@53612.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@53613.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@53614.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@53615.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@53621.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@53622.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@53617.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@53631.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@53632.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@53607.4 AXIProtocol.scala 81:19:@53629.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@53600.4 AXIProtocol.scala 82:21:@53630.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@53497.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@53496.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@53606.4 AXIProtocol.scala 84:20:@53634.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@53605.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@53604.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@53602.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@53601.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@53599.4 AXIProtocol.scala 86:22:@53636.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@53583.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@53584.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@53585.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@53586.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@53587.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@53588.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@53589.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@53590.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@53591.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@53592.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@53593.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@53594.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@53595.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@53596.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@53597.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@53598.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@53519.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@53520.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@53521.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@53522.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@53523.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@53524.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@53525.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@53526.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@53527.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@53528.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@53529.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@53530.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@53531.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@53532.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@53533.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@53534.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@53535.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@53536.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@53537.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@53538.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@53539.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@53540.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@53541.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@53542.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@53543.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@53544.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@53545.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@53546.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@53547.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@53548.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@53549.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@53550.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@53551.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@53552.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@53553.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@53554.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@53555.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@53556.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@53557.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@53558.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@53559.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@53560.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@53561.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@53562.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@53563.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@53564.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@53565.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@53566.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@53567.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@53568.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@53569.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@53570.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@53571.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@53572.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@53573.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@53574.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@53575.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@53576.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@53577.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@53578.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@53579.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@53580.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@53581.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@53582.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@53518.4 AXIProtocol.scala 87:27:@53637.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@53517.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@53498.4]
  assign wdataCounter_clock = clock; // @[:@53609.4]
  assign wdataCounter_reset = reset; // @[:@53610.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@53625.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@53626.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@53627.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@53639.2]
  input         clock, // @[:@53640.4]
  input         reset, // @[:@53641.4]
  input         io_enable, // @[:@53642.4]
  output        io_app_stores_0_cmd_ready, // @[:@53642.4]
  input         io_app_stores_0_cmd_valid, // @[:@53642.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@53642.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@53642.4]
  output        io_app_stores_0_data_ready, // @[:@53642.4]
  input         io_app_stores_0_data_valid, // @[:@53642.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@53642.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@53642.4]
  input         io_app_stores_0_wresp_ready, // @[:@53642.4]
  output        io_app_stores_0_wresp_valid, // @[:@53642.4]
  output        io_app_stores_0_wresp_bits, // @[:@53642.4]
  input         io_dram_cmd_ready, // @[:@53642.4]
  output        io_dram_cmd_valid, // @[:@53642.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@53642.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@53642.4]
  output        io_dram_cmd_bits_isWr, // @[:@53642.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@53642.4]
  input         io_dram_wdata_ready, // @[:@53642.4]
  output        io_dram_wdata_valid, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@53642.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@53642.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@53642.4]
  output        io_dram_wdata_bits_wlast, // @[:@53642.4]
  output        io_dram_rresp_ready, // @[:@53642.4]
  output        io_dram_wresp_ready, // @[:@53642.4]
  input         io_dram_wresp_valid, // @[:@53642.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@53642.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@54528.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@54542.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@54770.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@54885.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@54885.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@54528.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@54542.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@54770.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@54885.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@54541.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@54537.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@54532.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@54531.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@55110.4 DRAMArbiter.scala 100:23:@55113.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@55109.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@55108.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@55106.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@55105.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@55103.4 DRAMArbiter.scala 101:25:@55115.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@55087.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@55088.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@55089.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@55090.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@55091.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@55092.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@55093.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@55094.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@55095.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@55096.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@55097.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@55098.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@55099.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@55100.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@55101.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@55102.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@55023.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@55024.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@55025.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@55026.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@55027.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@55028.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@55029.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@55030.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@55031.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@55032.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@55033.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@55034.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@55035.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@55036.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@55037.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@55038.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@55039.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@55040.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@55041.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@55042.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@55043.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@55044.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@55045.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@55046.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@55047.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@55048.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@55049.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@55050.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@55051.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@55052.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@55053.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@55054.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@55055.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@55056.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@55057.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@55058.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@55059.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@55060.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@55061.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@55062.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@55063.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@55064.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@55065.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@55066.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@55067.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@55068.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@55069.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@55070.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@55071.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@55072.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@55073.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@55074.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@55075.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@55076.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@55077.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@55078.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@55079.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@55080.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@55081.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@55082.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@55083.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@55084.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@55085.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@55086.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@55022.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@55021.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@55002.4]
  assign StreamControllerStore_clock = clock; // @[:@54529.4]
  assign StreamControllerStore_reset = reset; // @[:@54530.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@54657.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@54650.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@54547.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@54540.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@54539.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@54538.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@54536.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@54535.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@54534.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@54533.4]
  assign StreamArbiter_clock = clock; // @[:@54543.4]
  assign StreamArbiter_reset = reset; // @[:@54544.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@54768.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@54767.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@54766.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@54764.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@54763.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@54761.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@54745.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@54746.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@54747.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@54748.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@54749.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@54750.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@54751.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@54752.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@54753.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@54754.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@54755.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@54756.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@54757.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@54758.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@54759.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@54760.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@54681.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@54682.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@54683.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@54684.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@54685.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@54686.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@54687.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@54688.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@54689.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@54690.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@54691.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@54692.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@54693.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@54694.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@54695.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@54696.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@54697.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@54698.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@54699.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@54700.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@54701.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@54702.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@54703.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@54704.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@54705.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@54706.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@54707.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@54708.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@54709.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@54710.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@54711.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@54712.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@54713.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@54714.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@54715.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@54716.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@54717.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@54718.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@54719.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@54720.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@54721.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@54722.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@54723.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@54724.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@54725.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@54726.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@54727.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@54728.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@54729.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@54730.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@54731.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@54732.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@54733.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@54734.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@54735.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@54736.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@54737.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@54738.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@54739.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@54740.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@54741.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@54742.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@54743.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@54744.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@54679.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@54660.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@54884.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@54877.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@54774.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@54773.4]
  assign AXICmdSplit_clock = clock; // @[:@54771.4]
  assign AXICmdSplit_reset = reset; // @[:@54772.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@54883.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@54882.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@54881.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@54879.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@54878.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@54876.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@54860.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@54861.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@54862.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@54863.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@54864.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@54865.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@54866.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@54867.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@54868.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@54869.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@54870.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@54871.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@54872.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@54873.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@54874.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@54875.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@54796.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@54797.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@54798.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@54799.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@54800.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@54801.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@54802.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@54803.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@54804.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@54805.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@54806.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@54807.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@54808.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@54809.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@54810.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@54811.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@54812.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@54813.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@54814.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@54815.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@54816.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@54817.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@54818.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@54819.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@54820.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@54821.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@54822.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@54823.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@54824.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@54825.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@54826.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@54827.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@54828.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@54829.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@54830.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@54831.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@54832.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@54833.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@54834.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@54835.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@54836.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@54837.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@54838.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@54839.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@54840.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@54841.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@54842.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@54843.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@54844.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@54845.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@54846.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@54847.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@54848.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@54849.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@54850.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@54851.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@54852.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@54853.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@54854.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@54855.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@54856.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@54857.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@54858.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@54859.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@54794.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@54775.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@54999.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@54992.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@54889.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@54888.4]
  assign AXICmdIssue_clock = clock; // @[:@54886.4]
  assign AXICmdIssue_reset = reset; // @[:@54887.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@54998.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@54997.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@54996.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@54994.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@54993.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@54991.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@54975.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@54976.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@54977.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@54978.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@54979.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@54980.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@54981.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@54982.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@54983.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@54984.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@54985.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@54986.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@54987.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@54988.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@54989.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@54990.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@54911.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@54912.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@54913.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@54914.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@54915.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@54916.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@54917.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@54918.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@54919.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@54920.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@54921.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@54922.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@54923.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@54924.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@54925.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@54926.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@54927.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@54928.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@54929.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@54930.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@54931.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@54932.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@54933.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@54934.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@54935.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@54936.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@54937.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@54938.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@54939.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@54940.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@54941.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@54942.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@54943.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@54944.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@54945.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@54946.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@54947.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@54948.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@54949.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@54950.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@54951.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@54952.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@54953.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@54954.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@54955.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@54956.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@54957.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@54958.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@54959.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@54960.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@54961.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@54962.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@54963.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@54964.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@54965.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@54966.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@54967.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@54968.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@54969.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@54970.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@54971.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@54972.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@54973.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@54974.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@54909.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@54890.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@55111.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@55104.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@55001.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@55000.4]
endmodule
module DRAMArbiter_1( // @[:@69340.2]
  input         clock, // @[:@69341.4]
  input         reset, // @[:@69342.4]
  input         io_enable, // @[:@69343.4]
  input         io_dram_cmd_ready, // @[:@69343.4]
  output        io_dram_cmd_valid, // @[:@69343.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@69343.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@69343.4]
  output        io_dram_cmd_bits_isWr, // @[:@69343.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@69343.4]
  input         io_dram_wdata_ready, // @[:@69343.4]
  output        io_dram_wdata_valid, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@69343.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@69343.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@69343.4]
  output        io_dram_wdata_bits_wlast, // @[:@69343.4]
  output        io_dram_rresp_ready, // @[:@69343.4]
  output        io_dram_wresp_ready, // @[:@69343.4]
  input         io_dram_wresp_valid, // @[:@69343.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@69343.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@70229.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@70243.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@70471.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@70586.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@70586.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@70229.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@70243.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@70471.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@70586.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@70811.4 DRAMArbiter.scala 100:23:@70814.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@70810.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@70809.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@70807.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@70806.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@70804.4 DRAMArbiter.scala 101:25:@70816.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@70788.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@70789.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@70790.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@70791.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@70792.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@70793.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@70794.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@70795.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@70796.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@70797.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@70798.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@70799.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@70800.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@70801.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@70802.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@70803.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@70724.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@70725.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@70726.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@70727.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@70728.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@70729.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@70730.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@70731.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@70732.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@70733.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@70734.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@70735.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@70736.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@70737.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@70738.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@70739.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@70740.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@70741.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@70742.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@70743.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@70744.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@70745.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@70746.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@70747.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@70748.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@70749.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@70750.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@70751.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@70752.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@70753.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@70754.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@70755.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@70756.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@70757.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@70758.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@70759.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@70760.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@70761.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@70762.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@70763.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@70764.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@70765.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@70766.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@70767.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@70768.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@70769.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@70770.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@70771.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@70772.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@70773.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@70774.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@70775.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@70776.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@70777.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@70778.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@70779.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@70780.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@70781.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@70782.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@70783.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@70784.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@70785.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@70786.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@70787.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@70723.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@70722.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@70703.4]
  assign StreamControllerStore_clock = clock; // @[:@70230.4]
  assign StreamControllerStore_reset = reset; // @[:@70231.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@70358.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@70351.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@70248.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@70241.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@70240.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@70239.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@70237.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@70236.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@70235.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@70234.4]
  assign StreamArbiter_clock = clock; // @[:@70244.4]
  assign StreamArbiter_reset = reset; // @[:@70245.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@70469.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@70468.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@70467.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@70465.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@70464.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@70462.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@70446.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@70447.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@70448.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@70449.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@70450.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@70451.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@70452.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@70453.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@70454.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@70455.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@70456.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@70457.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@70458.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@70459.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@70460.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@70461.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@70382.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@70383.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@70384.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@70385.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@70386.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@70387.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@70388.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@70389.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@70390.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@70391.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@70392.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@70393.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@70394.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@70395.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@70396.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@70397.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@70398.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@70399.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@70400.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@70401.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@70402.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@70403.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@70404.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@70405.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@70406.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@70407.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@70408.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@70409.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@70410.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@70411.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@70412.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@70413.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@70414.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@70415.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@70416.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@70417.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@70418.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@70419.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@70420.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@70421.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@70422.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@70423.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@70424.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@70425.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@70426.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@70427.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@70428.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@70429.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@70430.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@70431.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@70432.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@70433.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@70434.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@70435.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@70436.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@70437.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@70438.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@70439.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@70440.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@70441.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@70442.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@70443.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@70444.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@70445.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@70380.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@70361.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@70585.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@70578.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@70475.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@70474.4]
  assign AXICmdSplit_clock = clock; // @[:@70472.4]
  assign AXICmdSplit_reset = reset; // @[:@70473.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@70584.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@70583.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@70582.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@70580.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@70579.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@70577.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@70561.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@70562.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@70563.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@70564.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@70565.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@70566.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@70567.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@70568.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@70569.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@70570.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@70571.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@70572.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@70573.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@70574.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@70575.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@70576.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@70497.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@70498.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@70499.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@70500.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@70501.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@70502.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@70503.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@70504.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@70505.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@70506.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@70507.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@70508.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@70509.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@70510.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@70511.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@70512.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@70513.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@70514.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@70515.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@70516.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@70517.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@70518.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@70519.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@70520.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@70521.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@70522.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@70523.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@70524.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@70525.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@70526.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@70527.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@70528.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@70529.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@70530.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@70531.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@70532.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@70533.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@70534.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@70535.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@70536.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@70537.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@70538.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@70539.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@70540.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@70541.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@70542.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@70543.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@70544.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@70545.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@70546.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@70547.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@70548.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@70549.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@70550.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@70551.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@70552.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@70553.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@70554.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@70555.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@70556.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@70557.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@70558.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@70559.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@70560.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@70495.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@70476.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@70700.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@70693.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@70590.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@70589.4]
  assign AXICmdIssue_clock = clock; // @[:@70587.4]
  assign AXICmdIssue_reset = reset; // @[:@70588.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@70699.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@70698.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@70697.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@70695.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@70694.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@70692.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@70676.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@70677.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@70678.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@70679.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@70680.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@70681.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@70682.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@70683.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@70684.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@70685.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@70686.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@70687.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@70688.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@70689.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@70690.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@70691.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@70612.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@70613.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@70614.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@70615.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@70616.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@70617.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@70618.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@70619.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@70620.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@70621.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@70622.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@70623.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@70624.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@70625.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@70626.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@70627.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@70628.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@70629.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@70630.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@70631.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@70632.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@70633.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@70634.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@70635.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@70636.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@70637.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@70638.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@70639.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@70640.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@70641.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@70642.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@70643.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@70644.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@70645.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@70646.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@70647.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@70648.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@70649.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@70650.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@70651.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@70652.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@70653.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@70654.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@70655.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@70656.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@70657.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@70658.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@70659.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@70660.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@70661.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@70662.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@70663.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@70664.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@70665.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@70666.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@70667.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@70668.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@70669.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@70670.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@70671.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@70672.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@70673.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@70674.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@70675.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@70610.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@70591.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@70812.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@70805.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@70702.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@70701.4]
endmodule
module DRAMHeap( // @[:@101448.2]
  input         io_accel_0_req_valid, // @[:@101451.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@101451.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@101451.4]
  output        io_accel_0_resp_valid, // @[:@101451.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@101451.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@101451.4]
  output        io_host_0_req_valid, // @[:@101451.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@101451.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@101451.4]
  input         io_host_0_resp_valid, // @[:@101451.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@101451.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@101451.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@101458.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@101460.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@101459.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@101455.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@101454.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@101453.4]
endmodule
module FringeFF( // @[:@101494.2]
  input         clock, // @[:@101495.4]
  input         reset, // @[:@101496.4]
  input  [63:0] io_in, // @[:@101497.4]
  input         io_reset, // @[:@101497.4]
  output [63:0] io_out, // @[:@101497.4]
  input         io_enable // @[:@101497.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@101500.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@101500.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@101500.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@101500.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@101500.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@101505.4 package.scala 96:25:@101506.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@101511.6]
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@101500.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@101505.4 package.scala 96:25:@101506.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@101511.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@101517.4]
  assign RetimeWrapper_clock = clock; // @[:@101501.4]
  assign RetimeWrapper_reset = reset; // @[:@101502.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@101504.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@101503.4]
endmodule
module MuxN( // @[:@130133.2]
  input  [63:0] io_ins_0, // @[:@130136.4]
  input  [63:0] io_ins_1, // @[:@130136.4]
  input  [63:0] io_ins_2, // @[:@130136.4]
  input  [63:0] io_ins_3, // @[:@130136.4]
  input  [63:0] io_ins_4, // @[:@130136.4]
  input  [63:0] io_ins_5, // @[:@130136.4]
  input  [63:0] io_ins_6, // @[:@130136.4]
  input  [63:0] io_ins_7, // @[:@130136.4]
  input  [63:0] io_ins_8, // @[:@130136.4]
  input  [63:0] io_ins_9, // @[:@130136.4]
  input  [63:0] io_ins_10, // @[:@130136.4]
  input  [63:0] io_ins_11, // @[:@130136.4]
  input  [63:0] io_ins_12, // @[:@130136.4]
  input  [63:0] io_ins_13, // @[:@130136.4]
  input  [63:0] io_ins_14, // @[:@130136.4]
  input  [63:0] io_ins_15, // @[:@130136.4]
  input  [63:0] io_ins_16, // @[:@130136.4]
  input  [63:0] io_ins_17, // @[:@130136.4]
  input  [63:0] io_ins_18, // @[:@130136.4]
  input  [63:0] io_ins_19, // @[:@130136.4]
  input  [63:0] io_ins_20, // @[:@130136.4]
  input  [63:0] io_ins_21, // @[:@130136.4]
  input  [63:0] io_ins_22, // @[:@130136.4]
  input  [63:0] io_ins_23, // @[:@130136.4]
  input  [63:0] io_ins_24, // @[:@130136.4]
  input  [63:0] io_ins_25, // @[:@130136.4]
  input  [63:0] io_ins_26, // @[:@130136.4]
  input  [63:0] io_ins_27, // @[:@130136.4]
  input  [63:0] io_ins_28, // @[:@130136.4]
  input  [63:0] io_ins_29, // @[:@130136.4]
  input  [63:0] io_ins_30, // @[:@130136.4]
  input  [63:0] io_ins_31, // @[:@130136.4]
  input  [63:0] io_ins_32, // @[:@130136.4]
  input  [63:0] io_ins_33, // @[:@130136.4]
  input  [63:0] io_ins_34, // @[:@130136.4]
  input  [63:0] io_ins_35, // @[:@130136.4]
  input  [63:0] io_ins_36, // @[:@130136.4]
  input  [63:0] io_ins_37, // @[:@130136.4]
  input  [63:0] io_ins_38, // @[:@130136.4]
  input  [63:0] io_ins_39, // @[:@130136.4]
  input  [63:0] io_ins_40, // @[:@130136.4]
  input  [63:0] io_ins_41, // @[:@130136.4]
  input  [63:0] io_ins_42, // @[:@130136.4]
  input  [63:0] io_ins_43, // @[:@130136.4]
  input  [63:0] io_ins_44, // @[:@130136.4]
  input  [63:0] io_ins_45, // @[:@130136.4]
  input  [63:0] io_ins_46, // @[:@130136.4]
  input  [63:0] io_ins_47, // @[:@130136.4]
  input  [63:0] io_ins_48, // @[:@130136.4]
  input  [63:0] io_ins_49, // @[:@130136.4]
  input  [63:0] io_ins_50, // @[:@130136.4]
  input  [63:0] io_ins_51, // @[:@130136.4]
  input  [63:0] io_ins_52, // @[:@130136.4]
  input  [63:0] io_ins_53, // @[:@130136.4]
  input  [63:0] io_ins_54, // @[:@130136.4]
  input  [63:0] io_ins_55, // @[:@130136.4]
  input  [63:0] io_ins_56, // @[:@130136.4]
  input  [63:0] io_ins_57, // @[:@130136.4]
  input  [63:0] io_ins_58, // @[:@130136.4]
  input  [63:0] io_ins_59, // @[:@130136.4]
  input  [63:0] io_ins_60, // @[:@130136.4]
  input  [63:0] io_ins_61, // @[:@130136.4]
  input  [63:0] io_ins_62, // @[:@130136.4]
  input  [63:0] io_ins_63, // @[:@130136.4]
  input  [63:0] io_ins_64, // @[:@130136.4]
  input  [63:0] io_ins_65, // @[:@130136.4]
  input  [63:0] io_ins_66, // @[:@130136.4]
  input  [63:0] io_ins_67, // @[:@130136.4]
  input  [63:0] io_ins_68, // @[:@130136.4]
  input  [63:0] io_ins_69, // @[:@130136.4]
  input  [63:0] io_ins_70, // @[:@130136.4]
  input  [63:0] io_ins_71, // @[:@130136.4]
  input  [63:0] io_ins_72, // @[:@130136.4]
  input  [63:0] io_ins_73, // @[:@130136.4]
  input  [63:0] io_ins_74, // @[:@130136.4]
  input  [63:0] io_ins_75, // @[:@130136.4]
  input  [63:0] io_ins_76, // @[:@130136.4]
  input  [63:0] io_ins_77, // @[:@130136.4]
  input  [63:0] io_ins_78, // @[:@130136.4]
  input  [63:0] io_ins_79, // @[:@130136.4]
  input  [63:0] io_ins_80, // @[:@130136.4]
  input  [63:0] io_ins_81, // @[:@130136.4]
  input  [63:0] io_ins_82, // @[:@130136.4]
  input  [63:0] io_ins_83, // @[:@130136.4]
  input  [63:0] io_ins_84, // @[:@130136.4]
  input  [63:0] io_ins_85, // @[:@130136.4]
  input  [63:0] io_ins_86, // @[:@130136.4]
  input  [63:0] io_ins_87, // @[:@130136.4]
  input  [63:0] io_ins_88, // @[:@130136.4]
  input  [63:0] io_ins_89, // @[:@130136.4]
  input  [63:0] io_ins_90, // @[:@130136.4]
  input  [63:0] io_ins_91, // @[:@130136.4]
  input  [63:0] io_ins_92, // @[:@130136.4]
  input  [63:0] io_ins_93, // @[:@130136.4]
  input  [63:0] io_ins_94, // @[:@130136.4]
  input  [63:0] io_ins_95, // @[:@130136.4]
  input  [63:0] io_ins_96, // @[:@130136.4]
  input  [63:0] io_ins_97, // @[:@130136.4]
  input  [63:0] io_ins_98, // @[:@130136.4]
  input  [63:0] io_ins_99, // @[:@130136.4]
  input  [63:0] io_ins_100, // @[:@130136.4]
  input  [63:0] io_ins_101, // @[:@130136.4]
  input  [63:0] io_ins_102, // @[:@130136.4]
  input  [63:0] io_ins_103, // @[:@130136.4]
  input  [63:0] io_ins_104, // @[:@130136.4]
  input  [63:0] io_ins_105, // @[:@130136.4]
  input  [63:0] io_ins_106, // @[:@130136.4]
  input  [63:0] io_ins_107, // @[:@130136.4]
  input  [63:0] io_ins_108, // @[:@130136.4]
  input  [63:0] io_ins_109, // @[:@130136.4]
  input  [63:0] io_ins_110, // @[:@130136.4]
  input  [63:0] io_ins_111, // @[:@130136.4]
  input  [63:0] io_ins_112, // @[:@130136.4]
  input  [63:0] io_ins_113, // @[:@130136.4]
  input  [63:0] io_ins_114, // @[:@130136.4]
  input  [63:0] io_ins_115, // @[:@130136.4]
  input  [63:0] io_ins_116, // @[:@130136.4]
  input  [63:0] io_ins_117, // @[:@130136.4]
  input  [63:0] io_ins_118, // @[:@130136.4]
  input  [63:0] io_ins_119, // @[:@130136.4]
  input  [63:0] io_ins_120, // @[:@130136.4]
  input  [63:0] io_ins_121, // @[:@130136.4]
  input  [63:0] io_ins_122, // @[:@130136.4]
  input  [63:0] io_ins_123, // @[:@130136.4]
  input  [63:0] io_ins_124, // @[:@130136.4]
  input  [63:0] io_ins_125, // @[:@130136.4]
  input  [63:0] io_ins_126, // @[:@130136.4]
  input  [63:0] io_ins_127, // @[:@130136.4]
  input  [63:0] io_ins_128, // @[:@130136.4]
  input  [63:0] io_ins_129, // @[:@130136.4]
  input  [63:0] io_ins_130, // @[:@130136.4]
  input  [63:0] io_ins_131, // @[:@130136.4]
  input  [63:0] io_ins_132, // @[:@130136.4]
  input  [63:0] io_ins_133, // @[:@130136.4]
  input  [63:0] io_ins_134, // @[:@130136.4]
  input  [63:0] io_ins_135, // @[:@130136.4]
  input  [63:0] io_ins_136, // @[:@130136.4]
  input  [63:0] io_ins_137, // @[:@130136.4]
  input  [63:0] io_ins_138, // @[:@130136.4]
  input  [63:0] io_ins_139, // @[:@130136.4]
  input  [63:0] io_ins_140, // @[:@130136.4]
  input  [63:0] io_ins_141, // @[:@130136.4]
  input  [63:0] io_ins_142, // @[:@130136.4]
  input  [63:0] io_ins_143, // @[:@130136.4]
  input  [63:0] io_ins_144, // @[:@130136.4]
  input  [63:0] io_ins_145, // @[:@130136.4]
  input  [63:0] io_ins_146, // @[:@130136.4]
  input  [63:0] io_ins_147, // @[:@130136.4]
  input  [63:0] io_ins_148, // @[:@130136.4]
  input  [63:0] io_ins_149, // @[:@130136.4]
  input  [63:0] io_ins_150, // @[:@130136.4]
  input  [63:0] io_ins_151, // @[:@130136.4]
  input  [63:0] io_ins_152, // @[:@130136.4]
  input  [63:0] io_ins_153, // @[:@130136.4]
  input  [63:0] io_ins_154, // @[:@130136.4]
  input  [63:0] io_ins_155, // @[:@130136.4]
  input  [63:0] io_ins_156, // @[:@130136.4]
  input  [63:0] io_ins_157, // @[:@130136.4]
  input  [63:0] io_ins_158, // @[:@130136.4]
  input  [63:0] io_ins_159, // @[:@130136.4]
  input  [63:0] io_ins_160, // @[:@130136.4]
  input  [63:0] io_ins_161, // @[:@130136.4]
  input  [63:0] io_ins_162, // @[:@130136.4]
  input  [63:0] io_ins_163, // @[:@130136.4]
  input  [63:0] io_ins_164, // @[:@130136.4]
  input  [63:0] io_ins_165, // @[:@130136.4]
  input  [63:0] io_ins_166, // @[:@130136.4]
  input  [63:0] io_ins_167, // @[:@130136.4]
  input  [63:0] io_ins_168, // @[:@130136.4]
  input  [63:0] io_ins_169, // @[:@130136.4]
  input  [63:0] io_ins_170, // @[:@130136.4]
  input  [63:0] io_ins_171, // @[:@130136.4]
  input  [63:0] io_ins_172, // @[:@130136.4]
  input  [63:0] io_ins_173, // @[:@130136.4]
  input  [63:0] io_ins_174, // @[:@130136.4]
  input  [63:0] io_ins_175, // @[:@130136.4]
  input  [63:0] io_ins_176, // @[:@130136.4]
  input  [63:0] io_ins_177, // @[:@130136.4]
  input  [63:0] io_ins_178, // @[:@130136.4]
  input  [63:0] io_ins_179, // @[:@130136.4]
  input  [63:0] io_ins_180, // @[:@130136.4]
  input  [63:0] io_ins_181, // @[:@130136.4]
  input  [63:0] io_ins_182, // @[:@130136.4]
  input  [63:0] io_ins_183, // @[:@130136.4]
  input  [63:0] io_ins_184, // @[:@130136.4]
  input  [63:0] io_ins_185, // @[:@130136.4]
  input  [63:0] io_ins_186, // @[:@130136.4]
  input  [63:0] io_ins_187, // @[:@130136.4]
  input  [63:0] io_ins_188, // @[:@130136.4]
  input  [63:0] io_ins_189, // @[:@130136.4]
  input  [63:0] io_ins_190, // @[:@130136.4]
  input  [63:0] io_ins_191, // @[:@130136.4]
  input  [63:0] io_ins_192, // @[:@130136.4]
  input  [63:0] io_ins_193, // @[:@130136.4]
  input  [63:0] io_ins_194, // @[:@130136.4]
  input  [63:0] io_ins_195, // @[:@130136.4]
  input  [63:0] io_ins_196, // @[:@130136.4]
  input  [63:0] io_ins_197, // @[:@130136.4]
  input  [63:0] io_ins_198, // @[:@130136.4]
  input  [63:0] io_ins_199, // @[:@130136.4]
  input  [63:0] io_ins_200, // @[:@130136.4]
  input  [63:0] io_ins_201, // @[:@130136.4]
  input  [63:0] io_ins_202, // @[:@130136.4]
  input  [63:0] io_ins_203, // @[:@130136.4]
  input  [63:0] io_ins_204, // @[:@130136.4]
  input  [63:0] io_ins_205, // @[:@130136.4]
  input  [63:0] io_ins_206, // @[:@130136.4]
  input  [63:0] io_ins_207, // @[:@130136.4]
  input  [63:0] io_ins_208, // @[:@130136.4]
  input  [63:0] io_ins_209, // @[:@130136.4]
  input  [63:0] io_ins_210, // @[:@130136.4]
  input  [63:0] io_ins_211, // @[:@130136.4]
  input  [63:0] io_ins_212, // @[:@130136.4]
  input  [63:0] io_ins_213, // @[:@130136.4]
  input  [63:0] io_ins_214, // @[:@130136.4]
  input  [63:0] io_ins_215, // @[:@130136.4]
  input  [63:0] io_ins_216, // @[:@130136.4]
  input  [63:0] io_ins_217, // @[:@130136.4]
  input  [63:0] io_ins_218, // @[:@130136.4]
  input  [63:0] io_ins_219, // @[:@130136.4]
  input  [63:0] io_ins_220, // @[:@130136.4]
  input  [63:0] io_ins_221, // @[:@130136.4]
  input  [63:0] io_ins_222, // @[:@130136.4]
  input  [63:0] io_ins_223, // @[:@130136.4]
  input  [63:0] io_ins_224, // @[:@130136.4]
  input  [63:0] io_ins_225, // @[:@130136.4]
  input  [63:0] io_ins_226, // @[:@130136.4]
  input  [63:0] io_ins_227, // @[:@130136.4]
  input  [63:0] io_ins_228, // @[:@130136.4]
  input  [63:0] io_ins_229, // @[:@130136.4]
  input  [63:0] io_ins_230, // @[:@130136.4]
  input  [63:0] io_ins_231, // @[:@130136.4]
  input  [63:0] io_ins_232, // @[:@130136.4]
  input  [63:0] io_ins_233, // @[:@130136.4]
  input  [63:0] io_ins_234, // @[:@130136.4]
  input  [63:0] io_ins_235, // @[:@130136.4]
  input  [63:0] io_ins_236, // @[:@130136.4]
  input  [63:0] io_ins_237, // @[:@130136.4]
  input  [63:0] io_ins_238, // @[:@130136.4]
  input  [63:0] io_ins_239, // @[:@130136.4]
  input  [63:0] io_ins_240, // @[:@130136.4]
  input  [63:0] io_ins_241, // @[:@130136.4]
  input  [63:0] io_ins_242, // @[:@130136.4]
  input  [63:0] io_ins_243, // @[:@130136.4]
  input  [63:0] io_ins_244, // @[:@130136.4]
  input  [63:0] io_ins_245, // @[:@130136.4]
  input  [63:0] io_ins_246, // @[:@130136.4]
  input  [63:0] io_ins_247, // @[:@130136.4]
  input  [63:0] io_ins_248, // @[:@130136.4]
  input  [63:0] io_ins_249, // @[:@130136.4]
  input  [63:0] io_ins_250, // @[:@130136.4]
  input  [63:0] io_ins_251, // @[:@130136.4]
  input  [63:0] io_ins_252, // @[:@130136.4]
  input  [63:0] io_ins_253, // @[:@130136.4]
  input  [63:0] io_ins_254, // @[:@130136.4]
  input  [63:0] io_ins_255, // @[:@130136.4]
  input  [63:0] io_ins_256, // @[:@130136.4]
  input  [63:0] io_ins_257, // @[:@130136.4]
  input  [63:0] io_ins_258, // @[:@130136.4]
  input  [63:0] io_ins_259, // @[:@130136.4]
  input  [63:0] io_ins_260, // @[:@130136.4]
  input  [63:0] io_ins_261, // @[:@130136.4]
  input  [63:0] io_ins_262, // @[:@130136.4]
  input  [63:0] io_ins_263, // @[:@130136.4]
  input  [63:0] io_ins_264, // @[:@130136.4]
  input  [63:0] io_ins_265, // @[:@130136.4]
  input  [63:0] io_ins_266, // @[:@130136.4]
  input  [63:0] io_ins_267, // @[:@130136.4]
  input  [63:0] io_ins_268, // @[:@130136.4]
  input  [63:0] io_ins_269, // @[:@130136.4]
  input  [63:0] io_ins_270, // @[:@130136.4]
  input  [63:0] io_ins_271, // @[:@130136.4]
  input  [63:0] io_ins_272, // @[:@130136.4]
  input  [63:0] io_ins_273, // @[:@130136.4]
  input  [63:0] io_ins_274, // @[:@130136.4]
  input  [63:0] io_ins_275, // @[:@130136.4]
  input  [63:0] io_ins_276, // @[:@130136.4]
  input  [63:0] io_ins_277, // @[:@130136.4]
  input  [63:0] io_ins_278, // @[:@130136.4]
  input  [63:0] io_ins_279, // @[:@130136.4]
  input  [63:0] io_ins_280, // @[:@130136.4]
  input  [63:0] io_ins_281, // @[:@130136.4]
  input  [63:0] io_ins_282, // @[:@130136.4]
  input  [63:0] io_ins_283, // @[:@130136.4]
  input  [63:0] io_ins_284, // @[:@130136.4]
  input  [63:0] io_ins_285, // @[:@130136.4]
  input  [63:0] io_ins_286, // @[:@130136.4]
  input  [63:0] io_ins_287, // @[:@130136.4]
  input  [63:0] io_ins_288, // @[:@130136.4]
  input  [63:0] io_ins_289, // @[:@130136.4]
  input  [63:0] io_ins_290, // @[:@130136.4]
  input  [63:0] io_ins_291, // @[:@130136.4]
  input  [63:0] io_ins_292, // @[:@130136.4]
  input  [63:0] io_ins_293, // @[:@130136.4]
  input  [63:0] io_ins_294, // @[:@130136.4]
  input  [63:0] io_ins_295, // @[:@130136.4]
  input  [63:0] io_ins_296, // @[:@130136.4]
  input  [63:0] io_ins_297, // @[:@130136.4]
  input  [63:0] io_ins_298, // @[:@130136.4]
  input  [63:0] io_ins_299, // @[:@130136.4]
  input  [63:0] io_ins_300, // @[:@130136.4]
  input  [63:0] io_ins_301, // @[:@130136.4]
  input  [63:0] io_ins_302, // @[:@130136.4]
  input  [63:0] io_ins_303, // @[:@130136.4]
  input  [63:0] io_ins_304, // @[:@130136.4]
  input  [63:0] io_ins_305, // @[:@130136.4]
  input  [63:0] io_ins_306, // @[:@130136.4]
  input  [63:0] io_ins_307, // @[:@130136.4]
  input  [63:0] io_ins_308, // @[:@130136.4]
  input  [63:0] io_ins_309, // @[:@130136.4]
  input  [63:0] io_ins_310, // @[:@130136.4]
  input  [63:0] io_ins_311, // @[:@130136.4]
  input  [63:0] io_ins_312, // @[:@130136.4]
  input  [63:0] io_ins_313, // @[:@130136.4]
  input  [63:0] io_ins_314, // @[:@130136.4]
  input  [63:0] io_ins_315, // @[:@130136.4]
  input  [63:0] io_ins_316, // @[:@130136.4]
  input  [63:0] io_ins_317, // @[:@130136.4]
  input  [63:0] io_ins_318, // @[:@130136.4]
  input  [63:0] io_ins_319, // @[:@130136.4]
  input  [63:0] io_ins_320, // @[:@130136.4]
  input  [63:0] io_ins_321, // @[:@130136.4]
  input  [63:0] io_ins_322, // @[:@130136.4]
  input  [63:0] io_ins_323, // @[:@130136.4]
  input  [63:0] io_ins_324, // @[:@130136.4]
  input  [63:0] io_ins_325, // @[:@130136.4]
  input  [63:0] io_ins_326, // @[:@130136.4]
  input  [63:0] io_ins_327, // @[:@130136.4]
  input  [63:0] io_ins_328, // @[:@130136.4]
  input  [63:0] io_ins_329, // @[:@130136.4]
  input  [63:0] io_ins_330, // @[:@130136.4]
  input  [63:0] io_ins_331, // @[:@130136.4]
  input  [63:0] io_ins_332, // @[:@130136.4]
  input  [63:0] io_ins_333, // @[:@130136.4]
  input  [63:0] io_ins_334, // @[:@130136.4]
  input  [63:0] io_ins_335, // @[:@130136.4]
  input  [63:0] io_ins_336, // @[:@130136.4]
  input  [63:0] io_ins_337, // @[:@130136.4]
  input  [63:0] io_ins_338, // @[:@130136.4]
  input  [63:0] io_ins_339, // @[:@130136.4]
  input  [63:0] io_ins_340, // @[:@130136.4]
  input  [63:0] io_ins_341, // @[:@130136.4]
  input  [63:0] io_ins_342, // @[:@130136.4]
  input  [63:0] io_ins_343, // @[:@130136.4]
  input  [63:0] io_ins_344, // @[:@130136.4]
  input  [63:0] io_ins_345, // @[:@130136.4]
  input  [63:0] io_ins_346, // @[:@130136.4]
  input  [63:0] io_ins_347, // @[:@130136.4]
  input  [63:0] io_ins_348, // @[:@130136.4]
  input  [63:0] io_ins_349, // @[:@130136.4]
  input  [63:0] io_ins_350, // @[:@130136.4]
  input  [63:0] io_ins_351, // @[:@130136.4]
  input  [63:0] io_ins_352, // @[:@130136.4]
  input  [63:0] io_ins_353, // @[:@130136.4]
  input  [63:0] io_ins_354, // @[:@130136.4]
  input  [63:0] io_ins_355, // @[:@130136.4]
  input  [63:0] io_ins_356, // @[:@130136.4]
  input  [63:0] io_ins_357, // @[:@130136.4]
  input  [63:0] io_ins_358, // @[:@130136.4]
  input  [63:0] io_ins_359, // @[:@130136.4]
  input  [63:0] io_ins_360, // @[:@130136.4]
  input  [63:0] io_ins_361, // @[:@130136.4]
  input  [63:0] io_ins_362, // @[:@130136.4]
  input  [63:0] io_ins_363, // @[:@130136.4]
  input  [63:0] io_ins_364, // @[:@130136.4]
  input  [63:0] io_ins_365, // @[:@130136.4]
  input  [63:0] io_ins_366, // @[:@130136.4]
  input  [63:0] io_ins_367, // @[:@130136.4]
  input  [63:0] io_ins_368, // @[:@130136.4]
  input  [63:0] io_ins_369, // @[:@130136.4]
  input  [63:0] io_ins_370, // @[:@130136.4]
  input  [63:0] io_ins_371, // @[:@130136.4]
  input  [63:0] io_ins_372, // @[:@130136.4]
  input  [63:0] io_ins_373, // @[:@130136.4]
  input  [63:0] io_ins_374, // @[:@130136.4]
  input  [63:0] io_ins_375, // @[:@130136.4]
  input  [63:0] io_ins_376, // @[:@130136.4]
  input  [63:0] io_ins_377, // @[:@130136.4]
  input  [63:0] io_ins_378, // @[:@130136.4]
  input  [63:0] io_ins_379, // @[:@130136.4]
  input  [63:0] io_ins_380, // @[:@130136.4]
  input  [63:0] io_ins_381, // @[:@130136.4]
  input  [63:0] io_ins_382, // @[:@130136.4]
  input  [63:0] io_ins_383, // @[:@130136.4]
  input  [63:0] io_ins_384, // @[:@130136.4]
  input  [63:0] io_ins_385, // @[:@130136.4]
  input  [63:0] io_ins_386, // @[:@130136.4]
  input  [63:0] io_ins_387, // @[:@130136.4]
  input  [63:0] io_ins_388, // @[:@130136.4]
  input  [63:0] io_ins_389, // @[:@130136.4]
  input  [63:0] io_ins_390, // @[:@130136.4]
  input  [63:0] io_ins_391, // @[:@130136.4]
  input  [63:0] io_ins_392, // @[:@130136.4]
  input  [63:0] io_ins_393, // @[:@130136.4]
  input  [63:0] io_ins_394, // @[:@130136.4]
  input  [63:0] io_ins_395, // @[:@130136.4]
  input  [63:0] io_ins_396, // @[:@130136.4]
  input  [63:0] io_ins_397, // @[:@130136.4]
  input  [63:0] io_ins_398, // @[:@130136.4]
  input  [63:0] io_ins_399, // @[:@130136.4]
  input  [63:0] io_ins_400, // @[:@130136.4]
  input  [63:0] io_ins_401, // @[:@130136.4]
  input  [63:0] io_ins_402, // @[:@130136.4]
  input  [63:0] io_ins_403, // @[:@130136.4]
  input  [63:0] io_ins_404, // @[:@130136.4]
  input  [63:0] io_ins_405, // @[:@130136.4]
  input  [63:0] io_ins_406, // @[:@130136.4]
  input  [63:0] io_ins_407, // @[:@130136.4]
  input  [63:0] io_ins_408, // @[:@130136.4]
  input  [63:0] io_ins_409, // @[:@130136.4]
  input  [63:0] io_ins_410, // @[:@130136.4]
  input  [63:0] io_ins_411, // @[:@130136.4]
  input  [63:0] io_ins_412, // @[:@130136.4]
  input  [63:0] io_ins_413, // @[:@130136.4]
  input  [63:0] io_ins_414, // @[:@130136.4]
  input  [63:0] io_ins_415, // @[:@130136.4]
  input  [63:0] io_ins_416, // @[:@130136.4]
  input  [63:0] io_ins_417, // @[:@130136.4]
  input  [63:0] io_ins_418, // @[:@130136.4]
  input  [63:0] io_ins_419, // @[:@130136.4]
  input  [63:0] io_ins_420, // @[:@130136.4]
  input  [63:0] io_ins_421, // @[:@130136.4]
  input  [63:0] io_ins_422, // @[:@130136.4]
  input  [63:0] io_ins_423, // @[:@130136.4]
  input  [63:0] io_ins_424, // @[:@130136.4]
  input  [63:0] io_ins_425, // @[:@130136.4]
  input  [63:0] io_ins_426, // @[:@130136.4]
  input  [63:0] io_ins_427, // @[:@130136.4]
  input  [63:0] io_ins_428, // @[:@130136.4]
  input  [63:0] io_ins_429, // @[:@130136.4]
  input  [63:0] io_ins_430, // @[:@130136.4]
  input  [63:0] io_ins_431, // @[:@130136.4]
  input  [63:0] io_ins_432, // @[:@130136.4]
  input  [63:0] io_ins_433, // @[:@130136.4]
  input  [63:0] io_ins_434, // @[:@130136.4]
  input  [63:0] io_ins_435, // @[:@130136.4]
  input  [63:0] io_ins_436, // @[:@130136.4]
  input  [63:0] io_ins_437, // @[:@130136.4]
  input  [63:0] io_ins_438, // @[:@130136.4]
  input  [63:0] io_ins_439, // @[:@130136.4]
  input  [63:0] io_ins_440, // @[:@130136.4]
  input  [63:0] io_ins_441, // @[:@130136.4]
  input  [63:0] io_ins_442, // @[:@130136.4]
  input  [63:0] io_ins_443, // @[:@130136.4]
  input  [63:0] io_ins_444, // @[:@130136.4]
  input  [63:0] io_ins_445, // @[:@130136.4]
  input  [63:0] io_ins_446, // @[:@130136.4]
  input  [63:0] io_ins_447, // @[:@130136.4]
  input  [63:0] io_ins_448, // @[:@130136.4]
  input  [63:0] io_ins_449, // @[:@130136.4]
  input  [63:0] io_ins_450, // @[:@130136.4]
  input  [63:0] io_ins_451, // @[:@130136.4]
  input  [63:0] io_ins_452, // @[:@130136.4]
  input  [63:0] io_ins_453, // @[:@130136.4]
  input  [63:0] io_ins_454, // @[:@130136.4]
  input  [63:0] io_ins_455, // @[:@130136.4]
  input  [63:0] io_ins_456, // @[:@130136.4]
  input  [63:0] io_ins_457, // @[:@130136.4]
  input  [63:0] io_ins_458, // @[:@130136.4]
  input  [63:0] io_ins_459, // @[:@130136.4]
  input  [63:0] io_ins_460, // @[:@130136.4]
  input  [63:0] io_ins_461, // @[:@130136.4]
  input  [63:0] io_ins_462, // @[:@130136.4]
  input  [63:0] io_ins_463, // @[:@130136.4]
  input  [63:0] io_ins_464, // @[:@130136.4]
  input  [63:0] io_ins_465, // @[:@130136.4]
  input  [63:0] io_ins_466, // @[:@130136.4]
  input  [63:0] io_ins_467, // @[:@130136.4]
  input  [63:0] io_ins_468, // @[:@130136.4]
  input  [63:0] io_ins_469, // @[:@130136.4]
  input  [63:0] io_ins_470, // @[:@130136.4]
  input  [63:0] io_ins_471, // @[:@130136.4]
  input  [63:0] io_ins_472, // @[:@130136.4]
  input  [63:0] io_ins_473, // @[:@130136.4]
  input  [63:0] io_ins_474, // @[:@130136.4]
  input  [63:0] io_ins_475, // @[:@130136.4]
  input  [63:0] io_ins_476, // @[:@130136.4]
  input  [63:0] io_ins_477, // @[:@130136.4]
  input  [63:0] io_ins_478, // @[:@130136.4]
  input  [63:0] io_ins_479, // @[:@130136.4]
  input  [63:0] io_ins_480, // @[:@130136.4]
  input  [63:0] io_ins_481, // @[:@130136.4]
  input  [63:0] io_ins_482, // @[:@130136.4]
  input  [63:0] io_ins_483, // @[:@130136.4]
  input  [63:0] io_ins_484, // @[:@130136.4]
  input  [63:0] io_ins_485, // @[:@130136.4]
  input  [63:0] io_ins_486, // @[:@130136.4]
  input  [63:0] io_ins_487, // @[:@130136.4]
  input  [63:0] io_ins_488, // @[:@130136.4]
  input  [63:0] io_ins_489, // @[:@130136.4]
  input  [63:0] io_ins_490, // @[:@130136.4]
  input  [63:0] io_ins_491, // @[:@130136.4]
  input  [63:0] io_ins_492, // @[:@130136.4]
  input  [63:0] io_ins_493, // @[:@130136.4]
  input  [63:0] io_ins_494, // @[:@130136.4]
  input  [63:0] io_ins_495, // @[:@130136.4]
  input  [63:0] io_ins_496, // @[:@130136.4]
  input  [63:0] io_ins_497, // @[:@130136.4]
  input  [63:0] io_ins_498, // @[:@130136.4]
  input  [63:0] io_ins_499, // @[:@130136.4]
  input  [63:0] io_ins_500, // @[:@130136.4]
  input  [63:0] io_ins_501, // @[:@130136.4]
  input  [63:0] io_ins_502, // @[:@130136.4]
  input  [8:0]  io_sel, // @[:@130136.4]
  output [63:0] io_out // @[:@130136.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@130138.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@130138.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@130138.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@130138.4]
endmodule
module RegFile( // @[:@130140.2]
  input         clock, // @[:@130141.4]
  input         reset, // @[:@130142.4]
  input  [31:0] io_raddr, // @[:@130143.4]
  input         io_wen, // @[:@130143.4]
  input  [31:0] io_waddr, // @[:@130143.4]
  input  [63:0] io_wdata, // @[:@130143.4]
  output [63:0] io_rdata, // @[:@130143.4]
  input         io_reset, // @[:@130143.4]
  output [63:0] io_argIns_0, // @[:@130143.4]
  output [63:0] io_argIns_1, // @[:@130143.4]
  output [63:0] io_argIns_2, // @[:@130143.4]
  output [63:0] io_argIns_3, // @[:@130143.4]
  input         io_argOuts_0_valid, // @[:@130143.4]
  input  [63:0] io_argOuts_0_bits, // @[:@130143.4]
  input         io_argOuts_1_valid, // @[:@130143.4]
  input  [63:0] io_argOuts_1_bits // @[:@130143.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@132153.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@132153.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@132153.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@132153.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@132153.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@132153.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@132165.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@132165.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@132165.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@132165.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@132165.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@132165.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@132184.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@132184.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@132184.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@132184.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@132184.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@132184.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@132196.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@132196.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@132196.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@132196.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@132196.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@132196.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@132208.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@132208.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@132208.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@132208.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@132208.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@132208.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@132222.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@132222.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@132222.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@132222.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@132222.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@132222.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@132236.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@132236.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@132236.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@132236.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@132236.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@132236.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@132250.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@132250.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@132250.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@132250.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@132250.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@132250.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@132264.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@132264.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@132264.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@132264.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@132264.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@132264.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@132278.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@132278.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@132278.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@132278.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@132278.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@132278.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@132292.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@132292.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@132292.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@132292.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@132292.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@132292.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@132306.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@132306.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@132306.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@132306.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@132306.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@132306.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@132320.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@132320.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@132320.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@132320.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@132320.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@132320.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@132334.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@132334.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@132334.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@132334.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@132334.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@132334.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@132348.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@132348.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@132348.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@132348.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@132348.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@132348.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@132362.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@132362.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@132362.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@132362.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@132362.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@132362.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@132376.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@132376.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@132376.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@132376.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@132376.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@132376.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@132390.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@132390.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@132390.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@132390.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@132390.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@132390.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@132404.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@132404.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@132404.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@132404.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@132404.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@132404.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@132418.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@132418.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@132418.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@132418.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@132418.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@132418.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@132432.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@132432.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@132432.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@132432.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@132432.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@132432.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@132446.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@132446.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@132446.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@132446.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@132446.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@132446.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@132460.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@132460.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@132460.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@132460.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@132460.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@132460.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@132474.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@132474.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@132474.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@132474.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@132474.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@132474.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@132488.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@132488.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@132488.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@132488.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@132488.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@132488.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@132502.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@132502.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@132502.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@132502.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@132502.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@132502.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@132516.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@132516.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@132516.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@132516.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@132516.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@132516.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@132530.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@132530.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@132530.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@132530.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@132530.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@132530.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@132544.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@132544.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@132544.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@132544.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@132544.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@132544.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@132558.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@132558.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@132558.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@132558.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@132558.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@132558.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@132572.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@132572.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@132572.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@132572.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@132572.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@132572.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@132586.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@132586.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@132586.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@132586.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@132586.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@132586.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@132600.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@132600.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@132600.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@132600.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@132600.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@132600.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@132614.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@132614.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@132614.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@132614.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@132614.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@132614.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@132628.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@132628.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@132628.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@132628.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@132628.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@132628.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@132642.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@132642.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@132642.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@132642.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@132642.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@132642.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@132656.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@132656.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@132656.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@132656.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@132656.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@132656.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@132670.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@132670.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@132670.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@132670.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@132670.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@132670.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@132684.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@132684.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@132684.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@132684.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@132684.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@132684.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@132698.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@132698.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@132698.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@132698.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@132698.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@132698.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@132712.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@132712.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@132712.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@132712.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@132712.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@132712.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@132726.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@132726.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@132726.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@132726.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@132726.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@132726.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@132740.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@132740.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@132740.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@132740.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@132740.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@132740.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@132754.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@132754.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@132754.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@132768.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@132768.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@132768.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@132768.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@132768.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@132768.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@132782.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@132782.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@132782.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@132782.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@132782.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@132782.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@132796.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@132796.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@132796.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@132796.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@132796.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@132796.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@132810.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@132810.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@132810.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@132810.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@132810.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@132810.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@132824.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@132824.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@132824.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@132824.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@132824.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@132824.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@132838.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@132838.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@132838.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@132838.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@132838.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@132838.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@132852.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@132852.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@132852.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@132852.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@132852.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@132852.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@132866.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@132866.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@132866.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@132866.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@132866.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@132866.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@132880.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@132880.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@132880.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@132880.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@132880.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@132880.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@132894.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@132894.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@132894.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@132894.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@132894.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@132894.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@132908.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@132908.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@132908.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@132908.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@132908.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@132908.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@132922.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@132922.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@132922.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@132922.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@132922.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@132922.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@132936.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@132936.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@132936.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@132936.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@132936.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@132936.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@132950.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@132950.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@132950.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@132950.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@132950.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@132950.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@132964.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@132964.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@132964.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@132964.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@132964.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@132964.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@132978.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@132978.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@132978.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@132978.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@132978.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@132978.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@132992.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@132992.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@132992.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@132992.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@132992.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@132992.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@133006.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@133006.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@133006.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@133006.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@133006.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@133006.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@133020.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@133020.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@133020.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@133020.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@133020.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@133020.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@133034.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@133034.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@133034.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@133034.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@133034.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@133034.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@133048.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@133048.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@133048.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@133048.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@133048.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@133048.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@133062.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@133062.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@133062.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@133062.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@133062.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@133062.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@133076.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@133076.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@133076.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@133076.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@133076.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@133076.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@133090.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@133090.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@133090.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@133090.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@133090.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@133090.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@133104.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@133104.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@133104.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@133104.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@133104.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@133104.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@133118.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@133118.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@133118.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@133118.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@133118.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@133118.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@133132.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@133132.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@133132.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@133132.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@133132.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@133132.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@133146.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@133146.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@133146.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@133146.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@133146.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@133146.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@133160.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@133160.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@133160.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@133160.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@133160.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@133160.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@133174.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@133174.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@133174.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@133174.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@133174.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@133174.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@133188.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@133188.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@133188.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@133188.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@133188.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@133188.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@133202.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@133202.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@133202.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@133202.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@133202.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@133202.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@133216.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@133216.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@133216.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@133216.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@133216.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@133216.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@133230.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@133230.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@133230.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@133230.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@133230.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@133230.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@133244.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@133244.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@133244.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@133244.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@133244.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@133244.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@133258.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@133258.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@133258.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@133258.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@133258.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@133258.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@133272.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@133272.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@133272.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@133272.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@133272.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@133272.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@133286.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@133286.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@133286.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@133286.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@133286.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@133286.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@133300.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@133300.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@133300.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@133300.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@133300.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@133300.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@133314.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@133314.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@133314.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@133314.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@133314.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@133314.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@133328.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@133328.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@133328.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@133328.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@133328.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@133328.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@133342.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@133342.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@133342.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@133342.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@133342.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@133342.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@133356.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@133356.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@133356.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@133356.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@133356.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@133356.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@133370.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@133370.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@133370.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@133370.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@133370.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@133370.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@133384.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@133384.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@133384.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@133384.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@133384.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@133384.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@133398.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@133398.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@133398.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@133398.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@133398.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@133398.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@133412.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@133412.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@133412.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@133412.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@133412.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@133412.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@133426.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@133426.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@133426.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@133426.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@133426.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@133426.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@133440.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@133440.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@133440.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@133440.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@133440.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@133440.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@133454.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@133454.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@133454.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@133454.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@133454.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@133454.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@133468.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@133468.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@133468.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@133468.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@133468.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@133468.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@133482.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@133482.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@133482.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@133482.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@133482.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@133482.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@133496.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@133496.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@133496.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@133496.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@133496.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@133496.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@133510.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@133510.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@133510.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@133510.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@133510.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@133510.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@133524.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@133524.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@133524.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@133524.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@133524.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@133524.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@133538.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@133538.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@133538.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@133538.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@133538.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@133538.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@133552.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@133552.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@133552.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@133552.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@133552.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@133552.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@133566.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@133566.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@133566.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@133566.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@133566.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@133566.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@133580.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@133580.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@133580.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@133580.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@133580.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@133580.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@133594.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@133594.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@133594.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@133594.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@133594.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@133594.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@133608.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@133608.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@133608.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@133608.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@133608.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@133608.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@133622.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@133622.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@133622.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@133622.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@133622.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@133622.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@133636.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@133636.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@133636.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@133636.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@133636.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@133636.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@133650.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@133650.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@133650.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@133650.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@133650.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@133650.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@133664.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@133664.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@133664.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@133664.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@133664.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@133664.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@133678.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@133678.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@133678.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@133678.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@133678.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@133678.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@133692.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@133692.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@133692.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@133692.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@133692.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@133692.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@133706.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@133706.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@133706.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@133706.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@133706.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@133706.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@133720.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@133720.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@133720.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@133720.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@133720.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@133720.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@133734.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@133734.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@133734.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@133734.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@133734.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@133734.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@133748.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@133748.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@133748.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@133748.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@133748.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@133748.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@133762.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@133762.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@133762.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@133762.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@133762.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@133762.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@133776.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@133776.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@133776.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@133776.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@133776.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@133776.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@133790.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@133790.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@133790.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@133790.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@133790.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@133790.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@133804.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@133804.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@133804.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@133804.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@133804.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@133804.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@133818.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@133818.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@133818.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@133818.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@133818.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@133818.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@133832.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@133832.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@133832.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@133832.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@133832.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@133832.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@133846.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@133846.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@133846.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@133846.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@133846.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@133846.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@133860.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@133860.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@133860.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@133860.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@133860.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@133860.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@133874.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@133874.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@133874.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@133874.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@133874.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@133874.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@133888.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@133888.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@133888.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@133888.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@133888.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@133888.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@133902.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@133902.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@133902.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@133902.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@133902.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@133902.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@133916.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@133916.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@133916.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@133916.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@133916.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@133916.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@133930.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@133930.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@133930.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@133930.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@133930.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@133930.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@133944.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@133944.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@133944.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@133944.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@133944.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@133944.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@133958.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@133958.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@133958.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@133958.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@133958.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@133958.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@133972.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@133972.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@133972.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@133972.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@133972.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@133972.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@133986.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@133986.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@133986.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@133986.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@133986.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@133986.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@134000.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@134000.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@134000.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@134000.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@134000.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@134000.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@134014.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@134014.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@134014.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@134014.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@134014.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@134014.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@134028.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@134028.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@134028.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@134028.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@134028.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@134028.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@134042.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@134042.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@134042.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@134042.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@134042.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@134042.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@134056.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@134056.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@134056.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@134056.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@134056.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@134056.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@134070.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@134070.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@134070.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@134070.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@134070.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@134070.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@134084.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@134084.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@134084.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@134084.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@134084.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@134084.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@134098.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@134098.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@134098.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@134098.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@134098.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@134098.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@134112.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@134112.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@134112.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@134112.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@134112.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@134112.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@134126.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@134126.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@134126.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@134126.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@134126.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@134126.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@134140.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@134140.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@134140.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@134140.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@134140.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@134140.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@134154.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@134154.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@134154.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@134154.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@134154.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@134154.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@134168.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@134168.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@134168.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@134168.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@134168.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@134168.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@134182.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@134182.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@134182.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@134182.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@134182.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@134182.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@134196.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@134196.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@134196.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@134196.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@134196.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@134196.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@134210.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@134210.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@134210.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@134210.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@134210.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@134210.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@134224.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@134224.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@134224.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@134224.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@134224.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@134224.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@134238.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@134238.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@134238.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@134238.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@134238.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@134238.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@134252.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@134252.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@134252.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@134252.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@134252.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@134252.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@134266.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@134266.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@134266.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@134266.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@134266.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@134266.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@134280.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@134280.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@134280.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@134280.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@134280.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@134280.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@134294.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@134294.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@134294.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@134294.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@134294.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@134294.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@134308.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@134308.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@134308.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@134308.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@134308.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@134308.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@134322.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@134322.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@134322.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@134322.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@134322.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@134322.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@134336.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@134336.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@134336.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@134336.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@134336.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@134336.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@134350.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@134350.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@134350.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@134350.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@134350.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@134350.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@134364.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@134364.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@134364.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@134364.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@134364.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@134364.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@134378.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@134378.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@134378.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@134378.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@134378.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@134378.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@134392.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@134392.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@134392.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@134392.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@134392.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@134392.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@134406.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@134406.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@134406.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@134406.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@134406.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@134406.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@134420.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@134420.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@134420.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@134420.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@134420.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@134420.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@134434.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@134434.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@134434.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@134434.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@134434.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@134434.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@134448.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@134448.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@134448.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@134448.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@134448.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@134448.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@134462.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@134462.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@134462.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@134462.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@134462.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@134462.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@134476.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@134476.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@134476.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@134476.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@134476.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@134476.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@134490.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@134490.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@134490.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@134490.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@134490.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@134490.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@134504.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@134504.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@134504.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@134504.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@134504.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@134504.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@134518.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@134518.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@134518.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@134518.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@134518.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@134518.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@134532.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@134532.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@134532.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@134532.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@134532.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@134532.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@134546.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@134546.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@134546.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@134546.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@134546.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@134546.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@134560.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@134560.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@134560.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@134560.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@134560.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@134560.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@134574.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@134574.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@134574.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@134574.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@134574.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@134574.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@134588.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@134588.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@134588.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@134588.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@134588.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@134588.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@134602.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@134602.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@134602.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@134602.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@134602.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@134602.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@134616.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@134616.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@134616.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@134616.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@134616.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@134616.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@134630.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@134630.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@134630.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@134630.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@134630.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@134630.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@134644.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@134644.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@134644.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@134644.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@134644.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@134644.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@134658.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@134658.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@134658.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@134658.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@134658.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@134658.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@134672.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@134672.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@134672.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@134672.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@134672.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@134672.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@134686.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@134686.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@134686.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@134686.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@134686.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@134686.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@134700.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@134700.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@134700.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@134700.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@134700.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@134700.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@134714.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@134714.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@134714.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@134714.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@134714.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@134714.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@134728.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@134728.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@134728.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@134728.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@134728.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@134728.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@134742.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@134742.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@134742.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@134742.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@134742.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@134742.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@134756.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@134756.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@134756.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@134756.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@134756.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@134756.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@134770.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@134770.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@134770.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@134770.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@134770.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@134770.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@134784.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@134784.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@134784.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@134784.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@134784.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@134784.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@134798.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@134798.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@134798.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@134798.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@134798.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@134798.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@134812.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@134812.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@134812.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@134812.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@134812.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@134812.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@134826.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@134826.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@134826.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@134826.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@134826.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@134826.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@134840.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@134840.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@134840.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@134840.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@134840.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@134840.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@134854.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@134854.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@134854.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@134854.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@134854.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@134854.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@134868.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@134868.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@134868.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@134868.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@134868.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@134868.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@134882.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@134882.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@134882.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@134882.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@134882.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@134882.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@134896.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@134896.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@134896.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@134896.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@134896.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@134896.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@134910.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@134910.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@134910.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@134910.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@134910.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@134910.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@134924.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@134924.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@134924.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@134924.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@134924.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@134924.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@134938.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@134938.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@134938.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@134938.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@134938.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@134938.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@134952.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@134952.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@134952.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@134952.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@134952.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@134952.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@134966.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@134966.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@134966.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@134966.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@134966.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@134966.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@134980.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@134980.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@134980.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@134980.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@134980.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@134980.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@134994.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@134994.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@134994.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@134994.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@134994.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@134994.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@135008.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@135008.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@135008.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@135008.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@135008.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@135008.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@135022.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@135022.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@135022.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@135022.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@135022.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@135022.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@135036.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@135036.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@135036.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@135036.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@135036.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@135036.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@135050.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@135050.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@135050.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@135050.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@135050.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@135050.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@135064.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@135064.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@135064.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@135064.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@135064.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@135064.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@135078.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@135078.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@135078.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@135078.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@135078.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@135078.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@135092.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@135092.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@135092.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@135092.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@135092.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@135092.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@135106.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@135106.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@135106.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@135106.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@135106.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@135106.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@135120.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@135120.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@135120.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@135120.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@135120.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@135120.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@135134.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@135134.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@135134.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@135134.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@135134.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@135134.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@135148.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@135148.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@135148.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@135148.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@135148.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@135148.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@135162.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@135162.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@135162.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@135162.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@135162.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@135162.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@135176.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@135176.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@135176.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@135176.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@135176.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@135176.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@135190.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@135190.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@135190.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@135190.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@135190.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@135190.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@135204.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@135204.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@135204.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@135204.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@135204.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@135204.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@135218.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@135218.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@135218.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@135218.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@135218.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@135218.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@135232.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@135232.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@135232.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@135232.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@135232.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@135232.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@135246.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@135246.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@135246.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@135246.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@135246.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@135246.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@135260.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@135260.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@135260.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@135260.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@135260.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@135260.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@135274.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@135274.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@135274.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@135274.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@135274.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@135274.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@135288.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@135288.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@135288.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@135288.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@135288.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@135288.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@135302.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@135302.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@135302.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@135302.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@135302.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@135302.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@135316.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@135316.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@135316.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@135316.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@135316.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@135316.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@135330.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@135330.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@135330.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@135330.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@135330.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@135330.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@135344.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@135344.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@135344.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@135344.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@135344.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@135344.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@135358.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@135358.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@135358.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@135358.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@135358.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@135358.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@135372.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@135372.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@135372.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@135372.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@135372.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@135372.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@135386.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@135386.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@135386.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@135386.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@135386.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@135386.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@135400.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@135400.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@135400.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@135400.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@135400.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@135400.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@135414.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@135414.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@135414.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@135414.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@135414.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@135414.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@135428.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@135428.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@135428.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@135428.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@135428.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@135428.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@135442.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@135442.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@135442.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@135442.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@135442.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@135442.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@135456.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@135456.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@135456.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@135456.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@135456.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@135456.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@135470.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@135470.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@135470.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@135470.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@135470.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@135470.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@135484.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@135484.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@135484.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@135484.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@135484.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@135484.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@135498.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@135498.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@135498.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@135498.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@135498.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@135498.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@135512.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@135512.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@135512.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@135512.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@135512.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@135512.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@135526.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@135526.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@135526.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@135526.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@135526.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@135526.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@135540.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@135540.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@135540.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@135540.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@135540.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@135540.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@135554.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@135554.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@135554.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@135554.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@135554.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@135554.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@135568.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@135568.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@135568.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@135568.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@135568.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@135568.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@135582.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@135582.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@135582.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@135582.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@135582.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@135582.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@135596.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@135596.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@135596.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@135596.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@135596.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@135596.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@135610.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@135610.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@135610.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@135610.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@135610.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@135610.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@135624.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@135624.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@135624.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@135624.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@135624.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@135624.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@135638.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@135638.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@135638.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@135638.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@135638.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@135638.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@135652.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@135652.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@135652.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@135652.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@135652.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@135652.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@135666.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@135666.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@135666.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@135666.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@135666.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@135666.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@135680.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@135680.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@135680.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@135680.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@135680.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@135680.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@135694.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@135694.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@135694.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@135694.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@135694.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@135694.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@135708.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@135708.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@135708.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@135708.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@135708.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@135708.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@135722.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@135722.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@135722.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@135722.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@135722.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@135722.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@135736.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@135736.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@135736.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@135736.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@135736.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@135736.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@135750.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@135750.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@135750.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@135750.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@135750.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@135750.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@135764.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@135764.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@135764.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@135764.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@135764.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@135764.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@135778.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@135778.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@135778.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@135778.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@135778.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@135778.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@135792.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@135792.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@135792.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@135792.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@135792.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@135792.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@135806.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@135806.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@135806.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@135806.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@135806.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@135806.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@135820.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@135820.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@135820.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@135820.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@135820.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@135820.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@135834.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@135834.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@135834.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@135834.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@135834.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@135834.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@135848.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@135848.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@135848.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@135848.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@135848.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@135848.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@135862.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@135862.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@135862.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@135862.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@135862.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@135862.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@135876.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@135876.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@135876.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@135876.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@135876.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@135876.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@135890.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@135890.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@135890.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@135890.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@135890.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@135890.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@135904.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@135904.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@135904.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@135904.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@135904.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@135904.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@135918.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@135918.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@135918.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@135918.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@135918.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@135918.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@135932.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@135932.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@135932.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@135932.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@135932.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@135932.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@135946.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@135946.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@135946.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@135946.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@135946.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@135946.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@135960.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@135960.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@135960.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@135960.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@135960.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@135960.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@135974.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@135974.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@135974.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@135974.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@135974.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@135974.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@135988.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@135988.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@135988.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@135988.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@135988.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@135988.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@136002.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@136002.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@136002.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@136002.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@136002.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@136002.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@136016.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@136016.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@136016.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@136016.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@136016.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@136016.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@136030.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@136030.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@136030.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@136030.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@136030.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@136030.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@136044.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@136044.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@136044.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@136044.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@136044.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@136044.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@136058.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@136058.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@136058.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@136058.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@136058.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@136058.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@136072.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@136072.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@136072.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@136072.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@136072.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@136072.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@136086.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@136086.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@136086.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@136086.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@136086.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@136086.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@136100.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@136100.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@136100.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@136100.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@136100.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@136100.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@136114.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@136114.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@136114.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@136114.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@136114.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@136114.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@136128.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@136128.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@136128.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@136128.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@136128.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@136128.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@136142.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@136142.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@136142.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@136142.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@136142.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@136142.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@136156.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@136156.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@136156.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@136156.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@136156.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@136156.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@136170.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@136170.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@136170.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@136170.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@136170.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@136170.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@136184.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@136184.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@136184.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@136184.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@136184.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@136184.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@136198.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@136198.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@136198.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@136198.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@136198.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@136198.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@136212.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@136212.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@136212.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@136212.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@136212.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@136212.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@136226.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@136226.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@136226.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@136226.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@136226.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@136226.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@136240.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@136240.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@136240.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@136240.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@136240.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@136240.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@136254.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@136254.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@136254.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@136254.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@136254.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@136254.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@136268.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@136268.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@136268.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@136268.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@136268.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@136268.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@136282.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@136282.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@136282.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@136282.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@136282.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@136282.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@136296.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@136296.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@136296.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@136296.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@136296.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@136296.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@136310.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@136310.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@136310.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@136310.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@136310.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@136310.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@136324.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@136324.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@136324.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@136324.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@136324.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@136324.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@136338.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@136338.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@136338.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@136338.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@136338.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@136338.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@136352.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@136352.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@136352.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@136352.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@136352.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@136352.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@136366.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@136366.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@136366.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@136366.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@136366.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@136366.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@136380.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@136380.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@136380.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@136380.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@136380.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@136380.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@136394.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@136394.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@136394.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@136394.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@136394.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@136394.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@136408.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@136408.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@136408.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@136408.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@136408.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@136408.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@136422.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@136422.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@136422.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@136422.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@136422.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@136422.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@136436.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@136436.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@136436.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@136436.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@136436.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@136436.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@136450.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@136450.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@136450.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@136450.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@136450.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@136450.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@136464.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@136464.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@136464.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@136464.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@136464.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@136464.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@136478.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@136478.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@136478.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@136478.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@136478.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@136478.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@136492.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@136492.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@136492.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@136492.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@136492.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@136492.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@136506.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@136506.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@136506.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@136506.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@136506.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@136506.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@136520.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@136520.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@136520.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@136520.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@136520.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@136520.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@136534.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@136534.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@136534.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@136534.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@136534.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@136534.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@136548.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@136548.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@136548.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@136548.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@136548.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@136548.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@136562.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@136562.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@136562.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@136562.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@136562.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@136562.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@136576.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@136576.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@136576.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@136576.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@136576.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@136576.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@136590.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@136590.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@136590.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@136590.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@136590.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@136590.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@136604.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@136604.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@136604.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@136604.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@136604.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@136604.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@136618.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@136618.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@136618.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@136618.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@136618.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@136618.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@136632.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@136632.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@136632.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@136632.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@136632.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@136632.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@136646.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@136646.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@136646.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@136646.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@136646.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@136646.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@136660.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@136660.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@136660.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@136660.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@136660.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@136660.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@136674.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@136674.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@136674.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@136674.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@136674.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@136674.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@136688.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@136688.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@136688.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@136688.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@136688.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@136688.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@136702.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@136702.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@136702.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@136702.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@136702.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@136702.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@136716.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@136716.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@136716.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@136716.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@136716.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@136716.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@136730.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@136730.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@136730.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@136730.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@136730.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@136730.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@136744.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@136744.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@136744.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@136744.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@136744.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@136744.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@136758.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@136758.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@136758.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@136758.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@136758.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@136758.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@136772.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@136772.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@136772.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@136772.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@136772.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@136772.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@136786.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@136786.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@136786.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@136786.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@136786.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@136786.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@136800.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@136800.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@136800.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@136800.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@136800.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@136800.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@136814.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@136814.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@136814.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@136814.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@136814.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@136814.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@136828.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@136828.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@136828.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@136828.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@136828.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@136828.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@136842.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@136842.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@136842.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@136842.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@136842.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@136842.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@136856.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@136856.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@136856.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@136856.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@136856.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@136856.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@136870.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@136870.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@136870.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@136870.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@136870.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@136870.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@136884.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@136884.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@136884.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@136884.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@136884.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@136884.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@136898.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@136898.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@136898.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@136898.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@136898.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@136898.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@136912.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@136912.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@136912.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@136912.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@136912.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@136912.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@136926.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@136926.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@136926.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@136926.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@136926.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@136926.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@136940.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@136940.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@136940.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@136940.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@136940.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@136940.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@136954.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@136954.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@136954.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@136954.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@136954.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@136954.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@136968.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@136968.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@136968.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@136968.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@136968.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@136968.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@136982.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@136982.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@136982.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@136982.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@136982.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@136982.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@136996.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@136996.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@136996.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@136996.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@136996.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@136996.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@137010.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@137010.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@137010.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@137010.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@137010.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@137010.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@137024.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@137024.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@137024.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@137024.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@137024.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@137024.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@137038.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@137038.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@137038.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@137038.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@137038.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@137038.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@137052.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@137052.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@137052.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@137052.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@137052.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@137052.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@137066.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@137066.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@137066.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@137066.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@137066.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@137066.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@137080.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@137080.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@137080.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@137080.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@137080.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@137080.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@137094.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@137094.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@137094.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@137094.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@137094.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@137094.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@137108.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@137108.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@137108.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@137108.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@137108.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@137108.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@137122.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@137122.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@137122.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@137122.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@137122.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@137122.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@137136.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@137136.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@137136.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@137136.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@137136.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@137136.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@137150.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@137150.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@137150.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@137150.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@137150.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@137150.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@137164.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@137164.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@137164.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@137164.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@137164.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@137164.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@137178.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@137178.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@137178.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@137178.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@137178.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@137178.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@137192.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@137192.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@137192.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@137192.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@137192.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@137192.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@137206.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@137206.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@137206.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@137206.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@137206.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@137206.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@137220.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@137220.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@137220.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@137220.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@137220.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@137220.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@137234.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@137234.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@137234.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@137234.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@137234.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@137234.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@137248.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@137248.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@137248.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@137248.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@137248.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@137248.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@137262.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@137262.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@137262.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@137262.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@137262.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@137262.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@137276.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@137276.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@137276.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@137276.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@137276.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@137276.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@137290.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@137290.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@137290.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@137290.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@137290.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@137290.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@137304.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@137304.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@137304.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@137304.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@137304.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@137304.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@137318.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@137318.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@137318.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@137318.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@137318.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@137318.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@137332.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@137332.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@137332.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@137332.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@137332.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@137332.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@137346.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@137346.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@137346.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@137346.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@137346.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@137346.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@137360.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@137360.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@137360.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@137360.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@137360.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@137360.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@137374.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@137374.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@137374.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@137374.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@137374.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@137374.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@137388.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@137388.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@137388.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@137388.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@137388.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@137388.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@137402.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@137402.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@137402.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@137402.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@137402.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@137402.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@137416.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@137416.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@137416.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@137416.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@137416.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@137416.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@137430.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@137430.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@137430.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@137430.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@137430.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@137430.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@137444.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@137444.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@137444.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@137444.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@137444.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@137444.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@137458.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@137458.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@137458.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@137458.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@137458.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@137458.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@137472.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@137472.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@137472.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@137472.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@137472.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@137472.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@137486.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@137486.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@137486.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@137486.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@137486.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@137486.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@137500.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@137500.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@137500.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@137500.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@137500.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@137500.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@137514.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@137514.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@137514.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@137514.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@137514.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@137514.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@137528.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@137528.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@137528.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@137528.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@137528.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@137528.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@137542.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@137542.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@137542.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@137542.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@137542.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@137542.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@137556.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@137556.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@137556.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@137556.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@137556.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@137556.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@137570.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@137570.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@137570.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@137570.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@137570.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@137570.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@137584.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@137584.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@137584.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@137584.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@137584.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@137584.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@137598.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@137598.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@137598.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@137598.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@137598.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@137598.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@137612.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@137612.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@137612.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@137612.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@137612.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@137612.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@137626.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@137626.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@137626.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@137626.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@137626.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@137626.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@137640.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@137640.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@137640.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@137640.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@137640.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@137640.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@137654.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@137654.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@137654.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@137654.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@137654.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@137654.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@137668.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@137668.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@137668.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@137668.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@137668.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@137668.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@137682.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@137682.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@137682.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@137682.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@137682.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@137682.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@137696.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@137696.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@137696.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@137696.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@137696.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@137696.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@137710.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@137710.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@137710.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@137710.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@137710.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@137710.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@137724.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@137724.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@137724.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@137724.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@137724.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@137724.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@137738.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@137738.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@137738.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@137738.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@137738.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@137738.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@137752.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@137752.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@137752.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@137752.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@137752.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@137752.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@137766.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@137766.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@137766.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@137766.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@137766.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@137766.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@137780.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@137780.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@137780.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@137780.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@137780.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@137780.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@137794.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@137794.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@137794.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@137794.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@137794.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@137794.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@137808.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@137808.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@137808.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@137808.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@137808.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@137808.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@137822.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@137822.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@137822.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@137822.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@137822.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@137822.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@137836.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@137836.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@137836.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@137836.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@137836.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@137836.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@137850.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@137850.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@137850.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@137850.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@137850.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@137850.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@137864.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@137864.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@137864.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@137864.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@137864.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@137864.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@137878.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@137878.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@137878.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@137878.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@137878.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@137878.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@137892.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@137892.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@137892.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@137892.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@137892.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@137892.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@137906.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@137906.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@137906.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@137906.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@137906.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@137906.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@137920.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@137920.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@137920.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@137920.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@137920.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@137920.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@137934.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@137934.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@137934.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@137934.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@137934.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@137934.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@137948.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@137948.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@137948.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@137948.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@137948.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@137948.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@137962.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@137962.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@137962.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@137962.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@137962.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@137962.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@137976.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@137976.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@137976.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@137976.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@137976.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@137976.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@137990.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@137990.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@137990.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@137990.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@137990.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@137990.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@138004.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@138004.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@138004.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@138004.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@138004.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@138004.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@138018.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@138018.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@138018.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@138018.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@138018.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@138018.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@138032.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@138032.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@138032.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@138032.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@138032.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@138032.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@138046.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@138046.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@138046.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@138046.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@138046.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@138046.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@138060.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@138060.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@138060.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@138060.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@138060.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@138060.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@138074.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@138074.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@138074.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@138074.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@138074.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@138074.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@138088.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@138088.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@138088.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@138088.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@138088.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@138088.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@138102.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@138102.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@138102.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@138102.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@138102.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@138102.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@138116.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@138116.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@138116.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@138116.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@138116.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@138116.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@138130.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@138130.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@138130.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@138130.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@138130.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@138130.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@138144.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@138144.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@138144.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@138144.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@138144.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@138144.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@138158.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@138158.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@138158.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@138158.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@138158.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@138158.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@138172.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@138172.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@138172.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@138172.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@138172.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@138172.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@138186.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@138186.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@138186.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@138186.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@138186.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@138186.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@138200.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@138200.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@138200.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@138200.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@138200.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@138200.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@138214.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@138214.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@138214.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@138214.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@138214.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@138214.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@138228.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@138228.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@138228.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@138228.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@138228.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@138228.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@138242.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@138242.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@138242.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@138242.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@138242.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@138242.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@138256.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@138256.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@138256.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@138256.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@138256.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@138256.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@138270.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@138270.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@138270.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@138270.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@138270.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@138270.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@138284.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@138284.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@138284.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@138284.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@138284.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@138284.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@138298.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@138298.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@138298.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@138298.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@138298.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@138298.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@138312.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@138312.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@138312.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@138312.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@138312.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@138312.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@138326.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@138326.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@138326.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@138326.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@138326.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@138326.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@138340.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@138340.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@138340.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@138340.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@138340.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@138340.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@138354.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@138354.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@138354.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@138354.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@138354.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@138354.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@138368.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@138368.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@138368.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@138368.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@138368.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@138368.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@138382.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@138382.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@138382.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@138382.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@138382.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@138382.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@138396.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@138396.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@138396.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@138396.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@138396.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@138396.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@138410.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@138410.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@138410.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@138410.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@138410.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@138410.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@138424.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@138424.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@138424.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@138424.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@138424.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@138424.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@138438.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@138438.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@138438.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@138438.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@138438.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@138438.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@138452.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@138452.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@138452.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@138452.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@138452.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@138452.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@138466.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@138466.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@138466.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@138466.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@138466.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@138466.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@138480.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@138480.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@138480.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@138480.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@138480.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@138480.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@138494.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@138494.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@138494.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@138494.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@138494.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@138494.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@138508.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@138508.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@138508.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@138508.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@138508.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@138508.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@138522.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@138522.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@138522.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@138522.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@138522.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@138522.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@138536.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@138536.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@138536.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@138536.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@138536.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@138536.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@138550.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@138550.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@138550.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@138550.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@138550.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@138550.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@138564.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@138564.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@138564.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@138564.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@138564.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@138564.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@138578.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@138578.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@138578.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@138578.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@138578.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@138578.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@138592.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@138592.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@138592.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@138592.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@138592.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@138592.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@138606.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@138606.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@138606.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@138606.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@138606.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@138606.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@138620.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@138620.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@138620.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@138620.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@138620.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@138620.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@138634.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@138634.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@138634.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@138634.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@138634.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@138634.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@138648.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@138648.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@138648.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@138648.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@138648.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@138648.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@138662.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@138662.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@138662.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@138662.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@138662.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@138662.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@138676.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@138676.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@138676.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@138676.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@138676.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@138676.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@138690.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@138690.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@138690.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@138690.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@138690.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@138690.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@138704.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@138704.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@138704.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@138704.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@138704.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@138704.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@138718.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@138718.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@138718.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@138718.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@138718.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@138718.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@138732.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@138732.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@138732.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@138732.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@138732.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@138732.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@138746.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@138746.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@138746.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@138746.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@138746.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@138746.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@138760.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@138760.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@138760.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@138760.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@138760.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@138760.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@138774.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@138774.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@138774.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@138774.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@138774.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@138774.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@138788.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@138788.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@138788.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@138788.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@138788.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@138788.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@138802.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@138802.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@138802.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@138802.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@138802.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@138802.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@138816.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@138816.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@138816.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@138816.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@138816.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@138816.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@138830.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@138830.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@138830.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@138830.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@138830.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@138830.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@138844.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@138844.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@138844.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@138844.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@138844.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@138844.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@138858.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@138858.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@138858.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@138858.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@138858.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@138858.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@138872.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@138872.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@138872.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@138872.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@138872.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@138872.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@138886.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@138886.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@138886.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@138886.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@138886.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@138886.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@138900.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@138900.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@138900.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@138900.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@138900.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@138900.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@138914.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@138914.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@138914.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@138914.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@138914.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@138914.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@138928.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@138928.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@138928.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@138928.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@138928.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@138928.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@138942.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@138942.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@138942.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@138942.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@138942.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@138942.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@138956.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@138956.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@138956.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@138956.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@138956.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@138956.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@138970.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@138970.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@138970.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@138970.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@138970.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@138970.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@138984.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@138984.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@138984.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@138984.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@138984.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@138984.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@138998.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@138998.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@138998.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@138998.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@138998.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@138998.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@139012.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@139012.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@139012.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@139012.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@139012.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@139012.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@139026.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@139026.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@139026.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@139026.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@139026.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@139026.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@139040.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@139040.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@139040.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@139040.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@139040.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@139040.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@139054.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@139054.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@139054.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@139054.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@139054.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@139054.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@139068.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@139068.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@139068.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@139068.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@139068.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@139068.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@139082.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@139082.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@139082.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@139082.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@139082.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@139082.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@139096.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@139096.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@139096.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@139096.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@139096.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@139096.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@139110.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@139110.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@139110.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@139110.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@139110.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@139110.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@139124.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@139124.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@139124.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@139124.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@139124.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@139124.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@139138.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@139138.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@139138.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@139138.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@139138.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@139138.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@139152.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@139152.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@139152.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@139152.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@139152.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@139152.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@139166.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@139166.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@139166.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@139166.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@139166.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@139166.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@139180.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@139180.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@139180.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@139180.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@139180.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@139180.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@139194.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@139194.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@139194.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@132156.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@132168.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@132169.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@132187.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@132199.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@132211.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@132212.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@132153.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@132165.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@132184.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@132196.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@132208.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@132222.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@132236.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@132250.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@132264.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@132278.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@132292.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@132306.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@132320.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@132334.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@132348.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@132362.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@132376.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@132390.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@132404.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@132418.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@132432.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@132446.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@132460.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@132474.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@132488.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@132502.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@132516.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@132530.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@132544.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@132558.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@132572.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@132586.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@132600.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@132614.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@132628.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@132642.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@132656.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@132670.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@132684.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@132698.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@132712.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@132726.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@132740.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@132754.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@132768.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@132782.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@132796.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@132810.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@132824.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@132838.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@132852.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@132866.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@132880.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@132894.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@132908.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@132922.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@132936.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@132950.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@132964.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@132978.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@132992.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@133006.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@133020.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@133034.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@133048.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@133062.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@133076.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@133090.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@133104.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@133118.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@133132.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@133146.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@133160.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@133174.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@133188.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@133202.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@133216.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@133230.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@133244.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@133258.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@133272.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@133286.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@133300.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@133314.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@133328.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@133342.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@133356.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@133370.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@133384.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@133398.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@133412.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@133426.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@133440.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@133454.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@133468.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@133482.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@133496.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@133510.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@133524.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@133538.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@133552.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@133566.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@133580.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@133594.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@133608.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@133622.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@133636.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@133650.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@133664.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@133678.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@133692.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@133706.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@133720.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@133734.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@133748.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@133762.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@133776.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@133790.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@133804.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@133818.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@133832.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@133846.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@133860.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@133874.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@133888.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@133902.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@133916.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@133930.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@133944.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@133958.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@133972.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@133986.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@134000.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@134014.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@134028.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@134042.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@134056.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@134070.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@134084.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@134098.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@134112.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@134126.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@134140.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@134154.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@134168.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@134182.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@134196.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@134210.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@134224.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@134238.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@134252.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@134266.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@134280.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@134294.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@134308.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@134322.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@134336.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@134350.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@134364.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@134378.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@134392.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@134406.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@134420.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@134434.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@134448.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@134462.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@134476.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@134490.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@134504.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@134518.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@134532.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@134546.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@134560.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@134574.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@134588.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@134602.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@134616.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@134630.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@134644.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@134658.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@134672.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@134686.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@134700.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@134714.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@134728.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@134742.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@134756.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@134770.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@134784.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@134798.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@134812.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@134826.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@134840.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@134854.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@134868.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@134882.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@134896.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@134910.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@134924.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@134938.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@134952.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@134966.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@134980.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@134994.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@135008.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@135022.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@135036.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@135050.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@135064.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@135078.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@135092.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@135106.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@135120.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@135134.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@135148.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@135162.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@135176.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@135190.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@135204.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@135218.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@135232.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@135246.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@135260.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@135274.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@135288.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@135302.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@135316.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@135330.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@135344.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@135358.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@135372.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@135386.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@135400.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@135414.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@135428.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@135442.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@135456.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@135470.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@135484.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@135498.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@135512.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@135526.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@135540.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@135554.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@135568.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@135582.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@135596.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@135610.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@135624.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@135638.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@135652.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@135666.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@135680.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@135694.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@135708.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@135722.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@135736.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@135750.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@135764.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@135778.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@135792.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@135806.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@135820.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@135834.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@135848.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@135862.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@135876.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@135890.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@135904.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@135918.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@135932.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@135946.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@135960.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@135974.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@135988.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@136002.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@136016.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@136030.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@136044.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@136058.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@136072.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@136086.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@136100.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@136114.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@136128.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@136142.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@136156.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@136170.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@136184.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@136198.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@136212.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@136226.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@136240.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@136254.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@136268.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@136282.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@136296.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@136310.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@136324.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@136338.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@136352.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@136366.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@136380.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@136394.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@136408.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@136422.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@136436.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@136450.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@136464.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@136478.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@136492.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@136506.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@136520.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@136534.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@136548.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@136562.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@136576.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@136590.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@136604.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@136618.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@136632.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@136646.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@136660.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@136674.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@136688.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@136702.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@136716.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@136730.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@136744.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@136758.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@136772.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@136786.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@136800.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@136814.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@136828.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@136842.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@136856.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@136870.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@136884.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@136898.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@136912.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@136926.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@136940.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@136954.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@136968.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@136982.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@136996.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@137010.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@137024.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@137038.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@137052.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@137066.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@137080.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@137094.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@137108.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@137122.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@137136.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@137150.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@137164.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@137178.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@137192.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@137206.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@137220.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@137234.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@137248.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@137262.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@137276.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@137290.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@137304.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@137318.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@137332.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@137346.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@137360.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@137374.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@137388.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@137402.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@137416.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@137430.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@137444.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@137458.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@137472.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@137486.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@137500.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@137514.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@137528.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@137542.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@137556.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@137570.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@137584.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@137598.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@137612.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@137626.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@137640.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@137654.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@137668.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@137682.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@137696.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@137710.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@137724.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@137738.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@137752.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@137766.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@137780.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@137794.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@137808.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@137822.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@137836.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@137850.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@137864.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@137878.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@137892.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@137906.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@137920.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@137934.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@137948.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@137962.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@137976.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@137990.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@138004.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@138018.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@138032.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@138046.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@138060.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@138074.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@138088.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@138102.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@138116.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@138130.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@138144.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@138158.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@138172.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@138186.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@138200.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@138214.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@138228.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@138242.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@138256.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@138270.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@138284.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@138298.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@138312.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@138326.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@138340.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@138354.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@138368.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@138382.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@138396.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@138410.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@138424.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@138438.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@138452.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@138466.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@138480.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@138494.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@138508.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@138522.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@138536.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@138550.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@138564.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@138578.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@138592.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@138606.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@138620.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@138634.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@138648.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@138662.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@138676.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@138690.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@138704.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@138718.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@138732.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@138746.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@138760.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@138774.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@138788.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@138802.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@138816.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@138830.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@138844.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@138858.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@138872.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@138886.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@138900.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@138914.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@138928.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@138942.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@138956.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@138970.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@138984.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@138998.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@139012.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@139026.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@139040.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@139054.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@139068.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@139082.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@139096.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@139110.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@139124.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@139138.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@139152.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@139166.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@139180.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@139194.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@132156.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@132168.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@132169.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@132187.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@132199.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@132211.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@132212.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@140205.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@140211.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@140212.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@140213.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@140214.4]
  assign regs_0_clock = clock; // @[:@132154.4]
  assign regs_0_reset = reset; // @[:@132155.4 RegFile.scala 82:16:@132161.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@132159.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@132163.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@132158.4]
  assign regs_1_clock = clock; // @[:@132166.4]
  assign regs_1_reset = reset; // @[:@132167.4 RegFile.scala 70:16:@132179.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@132177.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@132182.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@132173.4]
  assign regs_2_clock = clock; // @[:@132185.4]
  assign regs_2_reset = reset; // @[:@132186.4 RegFile.scala 82:16:@132192.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@132190.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@132194.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@132189.4]
  assign regs_3_clock = clock; // @[:@132197.4]
  assign regs_3_reset = reset; // @[:@132198.4 RegFile.scala 82:16:@132204.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@132202.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@132206.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@132201.4]
  assign regs_4_clock = clock; // @[:@132209.4]
  assign regs_4_reset = io_reset; // @[:@132210.4 RegFile.scala 76:16:@132217.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@132216.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@132220.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@132214.4]
  assign regs_5_clock = clock; // @[:@132223.4]
  assign regs_5_reset = io_reset; // @[:@132224.4 RegFile.scala 76:16:@132231.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@132230.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@132234.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@132228.4]
  assign regs_6_clock = clock; // @[:@132237.4]
  assign regs_6_reset = io_reset; // @[:@132238.4 RegFile.scala 76:16:@132245.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@132244.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@132248.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@132242.4]
  assign regs_7_clock = clock; // @[:@132251.4]
  assign regs_7_reset = io_reset; // @[:@132252.4 RegFile.scala 76:16:@132259.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@132258.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@132262.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@132256.4]
  assign regs_8_clock = clock; // @[:@132265.4]
  assign regs_8_reset = io_reset; // @[:@132266.4 RegFile.scala 76:16:@132273.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@132272.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@132276.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@132270.4]
  assign regs_9_clock = clock; // @[:@132279.4]
  assign regs_9_reset = io_reset; // @[:@132280.4 RegFile.scala 76:16:@132287.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@132286.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@132290.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@132284.4]
  assign regs_10_clock = clock; // @[:@132293.4]
  assign regs_10_reset = io_reset; // @[:@132294.4 RegFile.scala 76:16:@132301.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@132300.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@132304.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@132298.4]
  assign regs_11_clock = clock; // @[:@132307.4]
  assign regs_11_reset = io_reset; // @[:@132308.4 RegFile.scala 76:16:@132315.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@132314.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@132318.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@132312.4]
  assign regs_12_clock = clock; // @[:@132321.4]
  assign regs_12_reset = io_reset; // @[:@132322.4 RegFile.scala 76:16:@132329.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@132328.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@132332.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@132326.4]
  assign regs_13_clock = clock; // @[:@132335.4]
  assign regs_13_reset = io_reset; // @[:@132336.4 RegFile.scala 76:16:@132343.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@132342.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@132346.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@132340.4]
  assign regs_14_clock = clock; // @[:@132349.4]
  assign regs_14_reset = io_reset; // @[:@132350.4 RegFile.scala 76:16:@132357.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@132356.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@132360.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@132354.4]
  assign regs_15_clock = clock; // @[:@132363.4]
  assign regs_15_reset = io_reset; // @[:@132364.4 RegFile.scala 76:16:@132371.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@132370.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@132374.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@132368.4]
  assign regs_16_clock = clock; // @[:@132377.4]
  assign regs_16_reset = io_reset; // @[:@132378.4 RegFile.scala 76:16:@132385.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@132384.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@132388.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@132382.4]
  assign regs_17_clock = clock; // @[:@132391.4]
  assign regs_17_reset = io_reset; // @[:@132392.4 RegFile.scala 76:16:@132399.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@132398.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@132402.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@132396.4]
  assign regs_18_clock = clock; // @[:@132405.4]
  assign regs_18_reset = io_reset; // @[:@132406.4 RegFile.scala 76:16:@132413.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@132412.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@132416.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@132410.4]
  assign regs_19_clock = clock; // @[:@132419.4]
  assign regs_19_reset = io_reset; // @[:@132420.4 RegFile.scala 76:16:@132427.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@132426.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@132430.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@132424.4]
  assign regs_20_clock = clock; // @[:@132433.4]
  assign regs_20_reset = io_reset; // @[:@132434.4 RegFile.scala 76:16:@132441.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@132440.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@132444.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@132438.4]
  assign regs_21_clock = clock; // @[:@132447.4]
  assign regs_21_reset = io_reset; // @[:@132448.4 RegFile.scala 76:16:@132455.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@132454.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@132458.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@132452.4]
  assign regs_22_clock = clock; // @[:@132461.4]
  assign regs_22_reset = io_reset; // @[:@132462.4 RegFile.scala 76:16:@132469.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@132468.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@132472.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@132466.4]
  assign regs_23_clock = clock; // @[:@132475.4]
  assign regs_23_reset = io_reset; // @[:@132476.4 RegFile.scala 76:16:@132483.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@132482.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@132486.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@132480.4]
  assign regs_24_clock = clock; // @[:@132489.4]
  assign regs_24_reset = io_reset; // @[:@132490.4 RegFile.scala 76:16:@132497.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@132496.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@132500.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@132494.4]
  assign regs_25_clock = clock; // @[:@132503.4]
  assign regs_25_reset = io_reset; // @[:@132504.4 RegFile.scala 76:16:@132511.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@132510.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@132514.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@132508.4]
  assign regs_26_clock = clock; // @[:@132517.4]
  assign regs_26_reset = io_reset; // @[:@132518.4 RegFile.scala 76:16:@132525.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@132524.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@132528.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@132522.4]
  assign regs_27_clock = clock; // @[:@132531.4]
  assign regs_27_reset = io_reset; // @[:@132532.4 RegFile.scala 76:16:@132539.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@132538.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@132542.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@132536.4]
  assign regs_28_clock = clock; // @[:@132545.4]
  assign regs_28_reset = io_reset; // @[:@132546.4 RegFile.scala 76:16:@132553.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@132552.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@132556.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@132550.4]
  assign regs_29_clock = clock; // @[:@132559.4]
  assign regs_29_reset = io_reset; // @[:@132560.4 RegFile.scala 76:16:@132567.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@132566.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@132570.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@132564.4]
  assign regs_30_clock = clock; // @[:@132573.4]
  assign regs_30_reset = io_reset; // @[:@132574.4 RegFile.scala 76:16:@132581.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@132580.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@132584.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@132578.4]
  assign regs_31_clock = clock; // @[:@132587.4]
  assign regs_31_reset = io_reset; // @[:@132588.4 RegFile.scala 76:16:@132595.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@132594.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@132598.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@132592.4]
  assign regs_32_clock = clock; // @[:@132601.4]
  assign regs_32_reset = io_reset; // @[:@132602.4 RegFile.scala 76:16:@132609.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@132608.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@132612.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@132606.4]
  assign regs_33_clock = clock; // @[:@132615.4]
  assign regs_33_reset = io_reset; // @[:@132616.4 RegFile.scala 76:16:@132623.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@132622.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@132626.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@132620.4]
  assign regs_34_clock = clock; // @[:@132629.4]
  assign regs_34_reset = io_reset; // @[:@132630.4 RegFile.scala 76:16:@132637.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@132636.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@132640.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@132634.4]
  assign regs_35_clock = clock; // @[:@132643.4]
  assign regs_35_reset = io_reset; // @[:@132644.4 RegFile.scala 76:16:@132651.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@132650.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@132654.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@132648.4]
  assign regs_36_clock = clock; // @[:@132657.4]
  assign regs_36_reset = io_reset; // @[:@132658.4 RegFile.scala 76:16:@132665.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@132664.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@132668.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@132662.4]
  assign regs_37_clock = clock; // @[:@132671.4]
  assign regs_37_reset = io_reset; // @[:@132672.4 RegFile.scala 76:16:@132679.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@132678.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@132682.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@132676.4]
  assign regs_38_clock = clock; // @[:@132685.4]
  assign regs_38_reset = io_reset; // @[:@132686.4 RegFile.scala 76:16:@132693.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@132692.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@132696.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@132690.4]
  assign regs_39_clock = clock; // @[:@132699.4]
  assign regs_39_reset = io_reset; // @[:@132700.4 RegFile.scala 76:16:@132707.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@132706.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@132710.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@132704.4]
  assign regs_40_clock = clock; // @[:@132713.4]
  assign regs_40_reset = io_reset; // @[:@132714.4 RegFile.scala 76:16:@132721.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@132720.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@132724.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@132718.4]
  assign regs_41_clock = clock; // @[:@132727.4]
  assign regs_41_reset = io_reset; // @[:@132728.4 RegFile.scala 76:16:@132735.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@132734.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@132738.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@132732.4]
  assign regs_42_clock = clock; // @[:@132741.4]
  assign regs_42_reset = io_reset; // @[:@132742.4 RegFile.scala 76:16:@132749.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@132748.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@132752.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@132746.4]
  assign regs_43_clock = clock; // @[:@132755.4]
  assign regs_43_reset = io_reset; // @[:@132756.4 RegFile.scala 76:16:@132763.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@132762.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@132766.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@132760.4]
  assign regs_44_clock = clock; // @[:@132769.4]
  assign regs_44_reset = io_reset; // @[:@132770.4 RegFile.scala 76:16:@132777.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@132776.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@132780.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@132774.4]
  assign regs_45_clock = clock; // @[:@132783.4]
  assign regs_45_reset = io_reset; // @[:@132784.4 RegFile.scala 76:16:@132791.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@132790.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@132794.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@132788.4]
  assign regs_46_clock = clock; // @[:@132797.4]
  assign regs_46_reset = io_reset; // @[:@132798.4 RegFile.scala 76:16:@132805.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@132804.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@132808.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@132802.4]
  assign regs_47_clock = clock; // @[:@132811.4]
  assign regs_47_reset = io_reset; // @[:@132812.4 RegFile.scala 76:16:@132819.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@132818.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@132822.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@132816.4]
  assign regs_48_clock = clock; // @[:@132825.4]
  assign regs_48_reset = io_reset; // @[:@132826.4 RegFile.scala 76:16:@132833.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@132832.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@132836.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@132830.4]
  assign regs_49_clock = clock; // @[:@132839.4]
  assign regs_49_reset = io_reset; // @[:@132840.4 RegFile.scala 76:16:@132847.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@132846.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@132850.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@132844.4]
  assign regs_50_clock = clock; // @[:@132853.4]
  assign regs_50_reset = io_reset; // @[:@132854.4 RegFile.scala 76:16:@132861.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@132860.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@132864.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@132858.4]
  assign regs_51_clock = clock; // @[:@132867.4]
  assign regs_51_reset = io_reset; // @[:@132868.4 RegFile.scala 76:16:@132875.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@132874.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@132878.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@132872.4]
  assign regs_52_clock = clock; // @[:@132881.4]
  assign regs_52_reset = io_reset; // @[:@132882.4 RegFile.scala 76:16:@132889.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@132888.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@132892.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@132886.4]
  assign regs_53_clock = clock; // @[:@132895.4]
  assign regs_53_reset = io_reset; // @[:@132896.4 RegFile.scala 76:16:@132903.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@132902.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@132906.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@132900.4]
  assign regs_54_clock = clock; // @[:@132909.4]
  assign regs_54_reset = io_reset; // @[:@132910.4 RegFile.scala 76:16:@132917.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@132916.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@132920.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@132914.4]
  assign regs_55_clock = clock; // @[:@132923.4]
  assign regs_55_reset = io_reset; // @[:@132924.4 RegFile.scala 76:16:@132931.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@132930.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@132934.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@132928.4]
  assign regs_56_clock = clock; // @[:@132937.4]
  assign regs_56_reset = io_reset; // @[:@132938.4 RegFile.scala 76:16:@132945.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@132944.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@132948.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@132942.4]
  assign regs_57_clock = clock; // @[:@132951.4]
  assign regs_57_reset = io_reset; // @[:@132952.4 RegFile.scala 76:16:@132959.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@132958.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@132962.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@132956.4]
  assign regs_58_clock = clock; // @[:@132965.4]
  assign regs_58_reset = io_reset; // @[:@132966.4 RegFile.scala 76:16:@132973.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@132972.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@132976.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@132970.4]
  assign regs_59_clock = clock; // @[:@132979.4]
  assign regs_59_reset = io_reset; // @[:@132980.4 RegFile.scala 76:16:@132987.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@132986.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@132990.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@132984.4]
  assign regs_60_clock = clock; // @[:@132993.4]
  assign regs_60_reset = io_reset; // @[:@132994.4 RegFile.scala 76:16:@133001.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@133000.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@133004.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@132998.4]
  assign regs_61_clock = clock; // @[:@133007.4]
  assign regs_61_reset = io_reset; // @[:@133008.4 RegFile.scala 76:16:@133015.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@133014.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@133018.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@133012.4]
  assign regs_62_clock = clock; // @[:@133021.4]
  assign regs_62_reset = io_reset; // @[:@133022.4 RegFile.scala 76:16:@133029.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@133028.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@133032.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@133026.4]
  assign regs_63_clock = clock; // @[:@133035.4]
  assign regs_63_reset = io_reset; // @[:@133036.4 RegFile.scala 76:16:@133043.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@133042.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@133046.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@133040.4]
  assign regs_64_clock = clock; // @[:@133049.4]
  assign regs_64_reset = io_reset; // @[:@133050.4 RegFile.scala 76:16:@133057.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@133056.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@133060.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@133054.4]
  assign regs_65_clock = clock; // @[:@133063.4]
  assign regs_65_reset = io_reset; // @[:@133064.4 RegFile.scala 76:16:@133071.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@133070.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@133074.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@133068.4]
  assign regs_66_clock = clock; // @[:@133077.4]
  assign regs_66_reset = io_reset; // @[:@133078.4 RegFile.scala 76:16:@133085.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@133084.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@133088.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@133082.4]
  assign regs_67_clock = clock; // @[:@133091.4]
  assign regs_67_reset = io_reset; // @[:@133092.4 RegFile.scala 76:16:@133099.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@133098.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@133102.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@133096.4]
  assign regs_68_clock = clock; // @[:@133105.4]
  assign regs_68_reset = io_reset; // @[:@133106.4 RegFile.scala 76:16:@133113.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@133112.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@133116.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@133110.4]
  assign regs_69_clock = clock; // @[:@133119.4]
  assign regs_69_reset = io_reset; // @[:@133120.4 RegFile.scala 76:16:@133127.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@133126.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@133130.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@133124.4]
  assign regs_70_clock = clock; // @[:@133133.4]
  assign regs_70_reset = io_reset; // @[:@133134.4 RegFile.scala 76:16:@133141.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@133140.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@133144.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@133138.4]
  assign regs_71_clock = clock; // @[:@133147.4]
  assign regs_71_reset = io_reset; // @[:@133148.4 RegFile.scala 76:16:@133155.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@133154.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@133158.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@133152.4]
  assign regs_72_clock = clock; // @[:@133161.4]
  assign regs_72_reset = io_reset; // @[:@133162.4 RegFile.scala 76:16:@133169.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@133168.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@133172.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@133166.4]
  assign regs_73_clock = clock; // @[:@133175.4]
  assign regs_73_reset = io_reset; // @[:@133176.4 RegFile.scala 76:16:@133183.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@133182.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@133186.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@133180.4]
  assign regs_74_clock = clock; // @[:@133189.4]
  assign regs_74_reset = io_reset; // @[:@133190.4 RegFile.scala 76:16:@133197.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@133196.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@133200.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@133194.4]
  assign regs_75_clock = clock; // @[:@133203.4]
  assign regs_75_reset = io_reset; // @[:@133204.4 RegFile.scala 76:16:@133211.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@133210.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@133214.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@133208.4]
  assign regs_76_clock = clock; // @[:@133217.4]
  assign regs_76_reset = io_reset; // @[:@133218.4 RegFile.scala 76:16:@133225.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@133224.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@133228.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@133222.4]
  assign regs_77_clock = clock; // @[:@133231.4]
  assign regs_77_reset = io_reset; // @[:@133232.4 RegFile.scala 76:16:@133239.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@133238.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@133242.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@133236.4]
  assign regs_78_clock = clock; // @[:@133245.4]
  assign regs_78_reset = io_reset; // @[:@133246.4 RegFile.scala 76:16:@133253.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@133252.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@133256.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@133250.4]
  assign regs_79_clock = clock; // @[:@133259.4]
  assign regs_79_reset = io_reset; // @[:@133260.4 RegFile.scala 76:16:@133267.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@133266.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@133270.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@133264.4]
  assign regs_80_clock = clock; // @[:@133273.4]
  assign regs_80_reset = io_reset; // @[:@133274.4 RegFile.scala 76:16:@133281.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@133280.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@133284.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@133278.4]
  assign regs_81_clock = clock; // @[:@133287.4]
  assign regs_81_reset = io_reset; // @[:@133288.4 RegFile.scala 76:16:@133295.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@133294.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@133298.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@133292.4]
  assign regs_82_clock = clock; // @[:@133301.4]
  assign regs_82_reset = io_reset; // @[:@133302.4 RegFile.scala 76:16:@133309.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@133308.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@133312.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@133306.4]
  assign regs_83_clock = clock; // @[:@133315.4]
  assign regs_83_reset = io_reset; // @[:@133316.4 RegFile.scala 76:16:@133323.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@133322.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@133326.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@133320.4]
  assign regs_84_clock = clock; // @[:@133329.4]
  assign regs_84_reset = io_reset; // @[:@133330.4 RegFile.scala 76:16:@133337.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@133336.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@133340.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@133334.4]
  assign regs_85_clock = clock; // @[:@133343.4]
  assign regs_85_reset = io_reset; // @[:@133344.4 RegFile.scala 76:16:@133351.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@133350.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@133354.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@133348.4]
  assign regs_86_clock = clock; // @[:@133357.4]
  assign regs_86_reset = io_reset; // @[:@133358.4 RegFile.scala 76:16:@133365.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@133364.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@133368.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@133362.4]
  assign regs_87_clock = clock; // @[:@133371.4]
  assign regs_87_reset = io_reset; // @[:@133372.4 RegFile.scala 76:16:@133379.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@133378.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@133382.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@133376.4]
  assign regs_88_clock = clock; // @[:@133385.4]
  assign regs_88_reset = io_reset; // @[:@133386.4 RegFile.scala 76:16:@133393.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@133392.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@133396.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@133390.4]
  assign regs_89_clock = clock; // @[:@133399.4]
  assign regs_89_reset = io_reset; // @[:@133400.4 RegFile.scala 76:16:@133407.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@133406.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@133410.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@133404.4]
  assign regs_90_clock = clock; // @[:@133413.4]
  assign regs_90_reset = io_reset; // @[:@133414.4 RegFile.scala 76:16:@133421.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@133420.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@133424.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@133418.4]
  assign regs_91_clock = clock; // @[:@133427.4]
  assign regs_91_reset = io_reset; // @[:@133428.4 RegFile.scala 76:16:@133435.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@133434.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@133438.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@133432.4]
  assign regs_92_clock = clock; // @[:@133441.4]
  assign regs_92_reset = io_reset; // @[:@133442.4 RegFile.scala 76:16:@133449.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@133448.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@133452.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@133446.4]
  assign regs_93_clock = clock; // @[:@133455.4]
  assign regs_93_reset = io_reset; // @[:@133456.4 RegFile.scala 76:16:@133463.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@133462.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@133466.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@133460.4]
  assign regs_94_clock = clock; // @[:@133469.4]
  assign regs_94_reset = io_reset; // @[:@133470.4 RegFile.scala 76:16:@133477.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@133476.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@133480.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@133474.4]
  assign regs_95_clock = clock; // @[:@133483.4]
  assign regs_95_reset = io_reset; // @[:@133484.4 RegFile.scala 76:16:@133491.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@133490.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@133494.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@133488.4]
  assign regs_96_clock = clock; // @[:@133497.4]
  assign regs_96_reset = io_reset; // @[:@133498.4 RegFile.scala 76:16:@133505.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@133504.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@133508.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@133502.4]
  assign regs_97_clock = clock; // @[:@133511.4]
  assign regs_97_reset = io_reset; // @[:@133512.4 RegFile.scala 76:16:@133519.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@133518.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@133522.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@133516.4]
  assign regs_98_clock = clock; // @[:@133525.4]
  assign regs_98_reset = io_reset; // @[:@133526.4 RegFile.scala 76:16:@133533.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@133532.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@133536.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@133530.4]
  assign regs_99_clock = clock; // @[:@133539.4]
  assign regs_99_reset = io_reset; // @[:@133540.4 RegFile.scala 76:16:@133547.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@133546.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@133550.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@133544.4]
  assign regs_100_clock = clock; // @[:@133553.4]
  assign regs_100_reset = io_reset; // @[:@133554.4 RegFile.scala 76:16:@133561.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@133560.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@133564.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@133558.4]
  assign regs_101_clock = clock; // @[:@133567.4]
  assign regs_101_reset = io_reset; // @[:@133568.4 RegFile.scala 76:16:@133575.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@133574.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@133578.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@133572.4]
  assign regs_102_clock = clock; // @[:@133581.4]
  assign regs_102_reset = io_reset; // @[:@133582.4 RegFile.scala 76:16:@133589.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@133588.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@133592.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@133586.4]
  assign regs_103_clock = clock; // @[:@133595.4]
  assign regs_103_reset = io_reset; // @[:@133596.4 RegFile.scala 76:16:@133603.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@133602.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@133606.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@133600.4]
  assign regs_104_clock = clock; // @[:@133609.4]
  assign regs_104_reset = io_reset; // @[:@133610.4 RegFile.scala 76:16:@133617.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@133616.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@133620.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@133614.4]
  assign regs_105_clock = clock; // @[:@133623.4]
  assign regs_105_reset = io_reset; // @[:@133624.4 RegFile.scala 76:16:@133631.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@133630.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@133634.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@133628.4]
  assign regs_106_clock = clock; // @[:@133637.4]
  assign regs_106_reset = io_reset; // @[:@133638.4 RegFile.scala 76:16:@133645.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@133644.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@133648.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@133642.4]
  assign regs_107_clock = clock; // @[:@133651.4]
  assign regs_107_reset = io_reset; // @[:@133652.4 RegFile.scala 76:16:@133659.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@133658.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@133662.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@133656.4]
  assign regs_108_clock = clock; // @[:@133665.4]
  assign regs_108_reset = io_reset; // @[:@133666.4 RegFile.scala 76:16:@133673.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@133672.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@133676.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@133670.4]
  assign regs_109_clock = clock; // @[:@133679.4]
  assign regs_109_reset = io_reset; // @[:@133680.4 RegFile.scala 76:16:@133687.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@133686.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@133690.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@133684.4]
  assign regs_110_clock = clock; // @[:@133693.4]
  assign regs_110_reset = io_reset; // @[:@133694.4 RegFile.scala 76:16:@133701.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@133700.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@133704.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@133698.4]
  assign regs_111_clock = clock; // @[:@133707.4]
  assign regs_111_reset = io_reset; // @[:@133708.4 RegFile.scala 76:16:@133715.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@133714.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@133718.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@133712.4]
  assign regs_112_clock = clock; // @[:@133721.4]
  assign regs_112_reset = io_reset; // @[:@133722.4 RegFile.scala 76:16:@133729.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@133728.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@133732.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@133726.4]
  assign regs_113_clock = clock; // @[:@133735.4]
  assign regs_113_reset = io_reset; // @[:@133736.4 RegFile.scala 76:16:@133743.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@133742.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@133746.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@133740.4]
  assign regs_114_clock = clock; // @[:@133749.4]
  assign regs_114_reset = io_reset; // @[:@133750.4 RegFile.scala 76:16:@133757.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@133756.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@133760.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@133754.4]
  assign regs_115_clock = clock; // @[:@133763.4]
  assign regs_115_reset = io_reset; // @[:@133764.4 RegFile.scala 76:16:@133771.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@133770.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@133774.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@133768.4]
  assign regs_116_clock = clock; // @[:@133777.4]
  assign regs_116_reset = io_reset; // @[:@133778.4 RegFile.scala 76:16:@133785.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@133784.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@133788.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@133782.4]
  assign regs_117_clock = clock; // @[:@133791.4]
  assign regs_117_reset = io_reset; // @[:@133792.4 RegFile.scala 76:16:@133799.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@133798.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@133802.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@133796.4]
  assign regs_118_clock = clock; // @[:@133805.4]
  assign regs_118_reset = io_reset; // @[:@133806.4 RegFile.scala 76:16:@133813.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@133812.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@133816.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@133810.4]
  assign regs_119_clock = clock; // @[:@133819.4]
  assign regs_119_reset = io_reset; // @[:@133820.4 RegFile.scala 76:16:@133827.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@133826.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@133830.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@133824.4]
  assign regs_120_clock = clock; // @[:@133833.4]
  assign regs_120_reset = io_reset; // @[:@133834.4 RegFile.scala 76:16:@133841.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@133840.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@133844.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@133838.4]
  assign regs_121_clock = clock; // @[:@133847.4]
  assign regs_121_reset = io_reset; // @[:@133848.4 RegFile.scala 76:16:@133855.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@133854.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@133858.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@133852.4]
  assign regs_122_clock = clock; // @[:@133861.4]
  assign regs_122_reset = io_reset; // @[:@133862.4 RegFile.scala 76:16:@133869.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@133868.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@133872.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@133866.4]
  assign regs_123_clock = clock; // @[:@133875.4]
  assign regs_123_reset = io_reset; // @[:@133876.4 RegFile.scala 76:16:@133883.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@133882.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@133886.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@133880.4]
  assign regs_124_clock = clock; // @[:@133889.4]
  assign regs_124_reset = io_reset; // @[:@133890.4 RegFile.scala 76:16:@133897.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@133896.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@133900.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@133894.4]
  assign regs_125_clock = clock; // @[:@133903.4]
  assign regs_125_reset = io_reset; // @[:@133904.4 RegFile.scala 76:16:@133911.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@133910.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@133914.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@133908.4]
  assign regs_126_clock = clock; // @[:@133917.4]
  assign regs_126_reset = io_reset; // @[:@133918.4 RegFile.scala 76:16:@133925.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@133924.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@133928.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@133922.4]
  assign regs_127_clock = clock; // @[:@133931.4]
  assign regs_127_reset = io_reset; // @[:@133932.4 RegFile.scala 76:16:@133939.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@133938.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@133942.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@133936.4]
  assign regs_128_clock = clock; // @[:@133945.4]
  assign regs_128_reset = io_reset; // @[:@133946.4 RegFile.scala 76:16:@133953.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@133952.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@133956.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@133950.4]
  assign regs_129_clock = clock; // @[:@133959.4]
  assign regs_129_reset = io_reset; // @[:@133960.4 RegFile.scala 76:16:@133967.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@133966.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@133970.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@133964.4]
  assign regs_130_clock = clock; // @[:@133973.4]
  assign regs_130_reset = io_reset; // @[:@133974.4 RegFile.scala 76:16:@133981.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@133980.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@133984.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@133978.4]
  assign regs_131_clock = clock; // @[:@133987.4]
  assign regs_131_reset = io_reset; // @[:@133988.4 RegFile.scala 76:16:@133995.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@133994.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@133998.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@133992.4]
  assign regs_132_clock = clock; // @[:@134001.4]
  assign regs_132_reset = io_reset; // @[:@134002.4 RegFile.scala 76:16:@134009.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@134008.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@134012.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@134006.4]
  assign regs_133_clock = clock; // @[:@134015.4]
  assign regs_133_reset = io_reset; // @[:@134016.4 RegFile.scala 76:16:@134023.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@134022.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@134026.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@134020.4]
  assign regs_134_clock = clock; // @[:@134029.4]
  assign regs_134_reset = io_reset; // @[:@134030.4 RegFile.scala 76:16:@134037.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@134036.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@134040.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@134034.4]
  assign regs_135_clock = clock; // @[:@134043.4]
  assign regs_135_reset = io_reset; // @[:@134044.4 RegFile.scala 76:16:@134051.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@134050.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@134054.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@134048.4]
  assign regs_136_clock = clock; // @[:@134057.4]
  assign regs_136_reset = io_reset; // @[:@134058.4 RegFile.scala 76:16:@134065.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@134064.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@134068.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@134062.4]
  assign regs_137_clock = clock; // @[:@134071.4]
  assign regs_137_reset = io_reset; // @[:@134072.4 RegFile.scala 76:16:@134079.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@134078.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@134082.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@134076.4]
  assign regs_138_clock = clock; // @[:@134085.4]
  assign regs_138_reset = io_reset; // @[:@134086.4 RegFile.scala 76:16:@134093.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@134092.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@134096.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@134090.4]
  assign regs_139_clock = clock; // @[:@134099.4]
  assign regs_139_reset = io_reset; // @[:@134100.4 RegFile.scala 76:16:@134107.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@134106.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@134110.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@134104.4]
  assign regs_140_clock = clock; // @[:@134113.4]
  assign regs_140_reset = io_reset; // @[:@134114.4 RegFile.scala 76:16:@134121.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@134120.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@134124.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@134118.4]
  assign regs_141_clock = clock; // @[:@134127.4]
  assign regs_141_reset = io_reset; // @[:@134128.4 RegFile.scala 76:16:@134135.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@134134.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@134138.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@134132.4]
  assign regs_142_clock = clock; // @[:@134141.4]
  assign regs_142_reset = io_reset; // @[:@134142.4 RegFile.scala 76:16:@134149.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@134148.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@134152.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@134146.4]
  assign regs_143_clock = clock; // @[:@134155.4]
  assign regs_143_reset = io_reset; // @[:@134156.4 RegFile.scala 76:16:@134163.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@134162.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@134166.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@134160.4]
  assign regs_144_clock = clock; // @[:@134169.4]
  assign regs_144_reset = io_reset; // @[:@134170.4 RegFile.scala 76:16:@134177.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@134176.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@134180.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@134174.4]
  assign regs_145_clock = clock; // @[:@134183.4]
  assign regs_145_reset = io_reset; // @[:@134184.4 RegFile.scala 76:16:@134191.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@134190.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@134194.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@134188.4]
  assign regs_146_clock = clock; // @[:@134197.4]
  assign regs_146_reset = io_reset; // @[:@134198.4 RegFile.scala 76:16:@134205.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@134204.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@134208.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@134202.4]
  assign regs_147_clock = clock; // @[:@134211.4]
  assign regs_147_reset = io_reset; // @[:@134212.4 RegFile.scala 76:16:@134219.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@134218.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@134222.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@134216.4]
  assign regs_148_clock = clock; // @[:@134225.4]
  assign regs_148_reset = io_reset; // @[:@134226.4 RegFile.scala 76:16:@134233.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@134232.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@134236.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@134230.4]
  assign regs_149_clock = clock; // @[:@134239.4]
  assign regs_149_reset = io_reset; // @[:@134240.4 RegFile.scala 76:16:@134247.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@134246.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@134250.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@134244.4]
  assign regs_150_clock = clock; // @[:@134253.4]
  assign regs_150_reset = io_reset; // @[:@134254.4 RegFile.scala 76:16:@134261.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@134260.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@134264.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@134258.4]
  assign regs_151_clock = clock; // @[:@134267.4]
  assign regs_151_reset = io_reset; // @[:@134268.4 RegFile.scala 76:16:@134275.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@134274.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@134278.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@134272.4]
  assign regs_152_clock = clock; // @[:@134281.4]
  assign regs_152_reset = io_reset; // @[:@134282.4 RegFile.scala 76:16:@134289.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@134288.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@134292.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@134286.4]
  assign regs_153_clock = clock; // @[:@134295.4]
  assign regs_153_reset = io_reset; // @[:@134296.4 RegFile.scala 76:16:@134303.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@134302.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@134306.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@134300.4]
  assign regs_154_clock = clock; // @[:@134309.4]
  assign regs_154_reset = io_reset; // @[:@134310.4 RegFile.scala 76:16:@134317.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@134316.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@134320.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@134314.4]
  assign regs_155_clock = clock; // @[:@134323.4]
  assign regs_155_reset = io_reset; // @[:@134324.4 RegFile.scala 76:16:@134331.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@134330.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@134334.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@134328.4]
  assign regs_156_clock = clock; // @[:@134337.4]
  assign regs_156_reset = io_reset; // @[:@134338.4 RegFile.scala 76:16:@134345.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@134344.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@134348.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@134342.4]
  assign regs_157_clock = clock; // @[:@134351.4]
  assign regs_157_reset = io_reset; // @[:@134352.4 RegFile.scala 76:16:@134359.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@134358.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@134362.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@134356.4]
  assign regs_158_clock = clock; // @[:@134365.4]
  assign regs_158_reset = io_reset; // @[:@134366.4 RegFile.scala 76:16:@134373.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@134372.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@134376.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@134370.4]
  assign regs_159_clock = clock; // @[:@134379.4]
  assign regs_159_reset = io_reset; // @[:@134380.4 RegFile.scala 76:16:@134387.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@134386.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@134390.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@134384.4]
  assign regs_160_clock = clock; // @[:@134393.4]
  assign regs_160_reset = io_reset; // @[:@134394.4 RegFile.scala 76:16:@134401.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@134400.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@134404.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@134398.4]
  assign regs_161_clock = clock; // @[:@134407.4]
  assign regs_161_reset = io_reset; // @[:@134408.4 RegFile.scala 76:16:@134415.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@134414.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@134418.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@134412.4]
  assign regs_162_clock = clock; // @[:@134421.4]
  assign regs_162_reset = io_reset; // @[:@134422.4 RegFile.scala 76:16:@134429.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@134428.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@134432.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@134426.4]
  assign regs_163_clock = clock; // @[:@134435.4]
  assign regs_163_reset = io_reset; // @[:@134436.4 RegFile.scala 76:16:@134443.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@134442.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@134446.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@134440.4]
  assign regs_164_clock = clock; // @[:@134449.4]
  assign regs_164_reset = io_reset; // @[:@134450.4 RegFile.scala 76:16:@134457.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@134456.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@134460.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@134454.4]
  assign regs_165_clock = clock; // @[:@134463.4]
  assign regs_165_reset = io_reset; // @[:@134464.4 RegFile.scala 76:16:@134471.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@134470.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@134474.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@134468.4]
  assign regs_166_clock = clock; // @[:@134477.4]
  assign regs_166_reset = io_reset; // @[:@134478.4 RegFile.scala 76:16:@134485.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@134484.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@134488.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@134482.4]
  assign regs_167_clock = clock; // @[:@134491.4]
  assign regs_167_reset = io_reset; // @[:@134492.4 RegFile.scala 76:16:@134499.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@134498.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@134502.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@134496.4]
  assign regs_168_clock = clock; // @[:@134505.4]
  assign regs_168_reset = io_reset; // @[:@134506.4 RegFile.scala 76:16:@134513.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@134512.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@134516.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@134510.4]
  assign regs_169_clock = clock; // @[:@134519.4]
  assign regs_169_reset = io_reset; // @[:@134520.4 RegFile.scala 76:16:@134527.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@134526.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@134530.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@134524.4]
  assign regs_170_clock = clock; // @[:@134533.4]
  assign regs_170_reset = io_reset; // @[:@134534.4 RegFile.scala 76:16:@134541.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@134540.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@134544.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@134538.4]
  assign regs_171_clock = clock; // @[:@134547.4]
  assign regs_171_reset = io_reset; // @[:@134548.4 RegFile.scala 76:16:@134555.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@134554.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@134558.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@134552.4]
  assign regs_172_clock = clock; // @[:@134561.4]
  assign regs_172_reset = io_reset; // @[:@134562.4 RegFile.scala 76:16:@134569.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@134568.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@134572.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@134566.4]
  assign regs_173_clock = clock; // @[:@134575.4]
  assign regs_173_reset = io_reset; // @[:@134576.4 RegFile.scala 76:16:@134583.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@134582.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@134586.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@134580.4]
  assign regs_174_clock = clock; // @[:@134589.4]
  assign regs_174_reset = io_reset; // @[:@134590.4 RegFile.scala 76:16:@134597.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@134596.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@134600.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@134594.4]
  assign regs_175_clock = clock; // @[:@134603.4]
  assign regs_175_reset = io_reset; // @[:@134604.4 RegFile.scala 76:16:@134611.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@134610.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@134614.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@134608.4]
  assign regs_176_clock = clock; // @[:@134617.4]
  assign regs_176_reset = io_reset; // @[:@134618.4 RegFile.scala 76:16:@134625.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@134624.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@134628.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@134622.4]
  assign regs_177_clock = clock; // @[:@134631.4]
  assign regs_177_reset = io_reset; // @[:@134632.4 RegFile.scala 76:16:@134639.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@134638.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@134642.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@134636.4]
  assign regs_178_clock = clock; // @[:@134645.4]
  assign regs_178_reset = io_reset; // @[:@134646.4 RegFile.scala 76:16:@134653.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@134652.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@134656.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@134650.4]
  assign regs_179_clock = clock; // @[:@134659.4]
  assign regs_179_reset = io_reset; // @[:@134660.4 RegFile.scala 76:16:@134667.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@134666.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@134670.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@134664.4]
  assign regs_180_clock = clock; // @[:@134673.4]
  assign regs_180_reset = io_reset; // @[:@134674.4 RegFile.scala 76:16:@134681.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@134680.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@134684.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@134678.4]
  assign regs_181_clock = clock; // @[:@134687.4]
  assign regs_181_reset = io_reset; // @[:@134688.4 RegFile.scala 76:16:@134695.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@134694.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@134698.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@134692.4]
  assign regs_182_clock = clock; // @[:@134701.4]
  assign regs_182_reset = io_reset; // @[:@134702.4 RegFile.scala 76:16:@134709.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@134708.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@134712.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@134706.4]
  assign regs_183_clock = clock; // @[:@134715.4]
  assign regs_183_reset = io_reset; // @[:@134716.4 RegFile.scala 76:16:@134723.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@134722.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@134726.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@134720.4]
  assign regs_184_clock = clock; // @[:@134729.4]
  assign regs_184_reset = io_reset; // @[:@134730.4 RegFile.scala 76:16:@134737.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@134736.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@134740.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@134734.4]
  assign regs_185_clock = clock; // @[:@134743.4]
  assign regs_185_reset = io_reset; // @[:@134744.4 RegFile.scala 76:16:@134751.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@134750.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@134754.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@134748.4]
  assign regs_186_clock = clock; // @[:@134757.4]
  assign regs_186_reset = io_reset; // @[:@134758.4 RegFile.scala 76:16:@134765.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@134764.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@134768.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@134762.4]
  assign regs_187_clock = clock; // @[:@134771.4]
  assign regs_187_reset = io_reset; // @[:@134772.4 RegFile.scala 76:16:@134779.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@134778.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@134782.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@134776.4]
  assign regs_188_clock = clock; // @[:@134785.4]
  assign regs_188_reset = io_reset; // @[:@134786.4 RegFile.scala 76:16:@134793.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@134792.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@134796.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@134790.4]
  assign regs_189_clock = clock; // @[:@134799.4]
  assign regs_189_reset = io_reset; // @[:@134800.4 RegFile.scala 76:16:@134807.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@134806.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@134810.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@134804.4]
  assign regs_190_clock = clock; // @[:@134813.4]
  assign regs_190_reset = io_reset; // @[:@134814.4 RegFile.scala 76:16:@134821.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@134820.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@134824.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@134818.4]
  assign regs_191_clock = clock; // @[:@134827.4]
  assign regs_191_reset = io_reset; // @[:@134828.4 RegFile.scala 76:16:@134835.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@134834.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@134838.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@134832.4]
  assign regs_192_clock = clock; // @[:@134841.4]
  assign regs_192_reset = io_reset; // @[:@134842.4 RegFile.scala 76:16:@134849.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@134848.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@134852.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@134846.4]
  assign regs_193_clock = clock; // @[:@134855.4]
  assign regs_193_reset = io_reset; // @[:@134856.4 RegFile.scala 76:16:@134863.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@134862.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@134866.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@134860.4]
  assign regs_194_clock = clock; // @[:@134869.4]
  assign regs_194_reset = io_reset; // @[:@134870.4 RegFile.scala 76:16:@134877.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@134876.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@134880.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@134874.4]
  assign regs_195_clock = clock; // @[:@134883.4]
  assign regs_195_reset = io_reset; // @[:@134884.4 RegFile.scala 76:16:@134891.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@134890.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@134894.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@134888.4]
  assign regs_196_clock = clock; // @[:@134897.4]
  assign regs_196_reset = io_reset; // @[:@134898.4 RegFile.scala 76:16:@134905.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@134904.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@134908.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@134902.4]
  assign regs_197_clock = clock; // @[:@134911.4]
  assign regs_197_reset = io_reset; // @[:@134912.4 RegFile.scala 76:16:@134919.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@134918.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@134922.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@134916.4]
  assign regs_198_clock = clock; // @[:@134925.4]
  assign regs_198_reset = io_reset; // @[:@134926.4 RegFile.scala 76:16:@134933.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@134932.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@134936.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@134930.4]
  assign regs_199_clock = clock; // @[:@134939.4]
  assign regs_199_reset = io_reset; // @[:@134940.4 RegFile.scala 76:16:@134947.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@134946.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@134950.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@134944.4]
  assign regs_200_clock = clock; // @[:@134953.4]
  assign regs_200_reset = io_reset; // @[:@134954.4 RegFile.scala 76:16:@134961.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@134960.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@134964.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@134958.4]
  assign regs_201_clock = clock; // @[:@134967.4]
  assign regs_201_reset = io_reset; // @[:@134968.4 RegFile.scala 76:16:@134975.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@134974.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@134978.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@134972.4]
  assign regs_202_clock = clock; // @[:@134981.4]
  assign regs_202_reset = io_reset; // @[:@134982.4 RegFile.scala 76:16:@134989.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@134988.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@134992.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@134986.4]
  assign regs_203_clock = clock; // @[:@134995.4]
  assign regs_203_reset = io_reset; // @[:@134996.4 RegFile.scala 76:16:@135003.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@135002.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@135006.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@135000.4]
  assign regs_204_clock = clock; // @[:@135009.4]
  assign regs_204_reset = io_reset; // @[:@135010.4 RegFile.scala 76:16:@135017.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@135016.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@135020.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@135014.4]
  assign regs_205_clock = clock; // @[:@135023.4]
  assign regs_205_reset = io_reset; // @[:@135024.4 RegFile.scala 76:16:@135031.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@135030.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@135034.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@135028.4]
  assign regs_206_clock = clock; // @[:@135037.4]
  assign regs_206_reset = io_reset; // @[:@135038.4 RegFile.scala 76:16:@135045.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@135044.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@135048.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@135042.4]
  assign regs_207_clock = clock; // @[:@135051.4]
  assign regs_207_reset = io_reset; // @[:@135052.4 RegFile.scala 76:16:@135059.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@135058.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@135062.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@135056.4]
  assign regs_208_clock = clock; // @[:@135065.4]
  assign regs_208_reset = io_reset; // @[:@135066.4 RegFile.scala 76:16:@135073.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@135072.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@135076.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@135070.4]
  assign regs_209_clock = clock; // @[:@135079.4]
  assign regs_209_reset = io_reset; // @[:@135080.4 RegFile.scala 76:16:@135087.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@135086.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@135090.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@135084.4]
  assign regs_210_clock = clock; // @[:@135093.4]
  assign regs_210_reset = io_reset; // @[:@135094.4 RegFile.scala 76:16:@135101.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@135100.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@135104.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@135098.4]
  assign regs_211_clock = clock; // @[:@135107.4]
  assign regs_211_reset = io_reset; // @[:@135108.4 RegFile.scala 76:16:@135115.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@135114.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@135118.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@135112.4]
  assign regs_212_clock = clock; // @[:@135121.4]
  assign regs_212_reset = io_reset; // @[:@135122.4 RegFile.scala 76:16:@135129.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@135128.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@135132.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@135126.4]
  assign regs_213_clock = clock; // @[:@135135.4]
  assign regs_213_reset = io_reset; // @[:@135136.4 RegFile.scala 76:16:@135143.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@135142.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@135146.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@135140.4]
  assign regs_214_clock = clock; // @[:@135149.4]
  assign regs_214_reset = io_reset; // @[:@135150.4 RegFile.scala 76:16:@135157.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@135156.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@135160.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@135154.4]
  assign regs_215_clock = clock; // @[:@135163.4]
  assign regs_215_reset = io_reset; // @[:@135164.4 RegFile.scala 76:16:@135171.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@135170.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@135174.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@135168.4]
  assign regs_216_clock = clock; // @[:@135177.4]
  assign regs_216_reset = io_reset; // @[:@135178.4 RegFile.scala 76:16:@135185.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@135184.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@135188.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@135182.4]
  assign regs_217_clock = clock; // @[:@135191.4]
  assign regs_217_reset = io_reset; // @[:@135192.4 RegFile.scala 76:16:@135199.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@135198.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@135202.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@135196.4]
  assign regs_218_clock = clock; // @[:@135205.4]
  assign regs_218_reset = io_reset; // @[:@135206.4 RegFile.scala 76:16:@135213.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@135212.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@135216.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@135210.4]
  assign regs_219_clock = clock; // @[:@135219.4]
  assign regs_219_reset = io_reset; // @[:@135220.4 RegFile.scala 76:16:@135227.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@135226.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@135230.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@135224.4]
  assign regs_220_clock = clock; // @[:@135233.4]
  assign regs_220_reset = io_reset; // @[:@135234.4 RegFile.scala 76:16:@135241.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@135240.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@135244.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@135238.4]
  assign regs_221_clock = clock; // @[:@135247.4]
  assign regs_221_reset = io_reset; // @[:@135248.4 RegFile.scala 76:16:@135255.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@135254.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@135258.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@135252.4]
  assign regs_222_clock = clock; // @[:@135261.4]
  assign regs_222_reset = io_reset; // @[:@135262.4 RegFile.scala 76:16:@135269.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@135268.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@135272.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@135266.4]
  assign regs_223_clock = clock; // @[:@135275.4]
  assign regs_223_reset = io_reset; // @[:@135276.4 RegFile.scala 76:16:@135283.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@135282.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@135286.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@135280.4]
  assign regs_224_clock = clock; // @[:@135289.4]
  assign regs_224_reset = io_reset; // @[:@135290.4 RegFile.scala 76:16:@135297.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@135296.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@135300.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@135294.4]
  assign regs_225_clock = clock; // @[:@135303.4]
  assign regs_225_reset = io_reset; // @[:@135304.4 RegFile.scala 76:16:@135311.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@135310.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@135314.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@135308.4]
  assign regs_226_clock = clock; // @[:@135317.4]
  assign regs_226_reset = io_reset; // @[:@135318.4 RegFile.scala 76:16:@135325.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@135324.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@135328.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@135322.4]
  assign regs_227_clock = clock; // @[:@135331.4]
  assign regs_227_reset = io_reset; // @[:@135332.4 RegFile.scala 76:16:@135339.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@135338.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@135342.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@135336.4]
  assign regs_228_clock = clock; // @[:@135345.4]
  assign regs_228_reset = io_reset; // @[:@135346.4 RegFile.scala 76:16:@135353.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@135352.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@135356.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@135350.4]
  assign regs_229_clock = clock; // @[:@135359.4]
  assign regs_229_reset = io_reset; // @[:@135360.4 RegFile.scala 76:16:@135367.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@135366.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@135370.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@135364.4]
  assign regs_230_clock = clock; // @[:@135373.4]
  assign regs_230_reset = io_reset; // @[:@135374.4 RegFile.scala 76:16:@135381.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@135380.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@135384.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@135378.4]
  assign regs_231_clock = clock; // @[:@135387.4]
  assign regs_231_reset = io_reset; // @[:@135388.4 RegFile.scala 76:16:@135395.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@135394.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@135398.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@135392.4]
  assign regs_232_clock = clock; // @[:@135401.4]
  assign regs_232_reset = io_reset; // @[:@135402.4 RegFile.scala 76:16:@135409.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@135408.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@135412.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@135406.4]
  assign regs_233_clock = clock; // @[:@135415.4]
  assign regs_233_reset = io_reset; // @[:@135416.4 RegFile.scala 76:16:@135423.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@135422.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@135426.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@135420.4]
  assign regs_234_clock = clock; // @[:@135429.4]
  assign regs_234_reset = io_reset; // @[:@135430.4 RegFile.scala 76:16:@135437.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@135436.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@135440.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@135434.4]
  assign regs_235_clock = clock; // @[:@135443.4]
  assign regs_235_reset = io_reset; // @[:@135444.4 RegFile.scala 76:16:@135451.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@135450.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@135454.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@135448.4]
  assign regs_236_clock = clock; // @[:@135457.4]
  assign regs_236_reset = io_reset; // @[:@135458.4 RegFile.scala 76:16:@135465.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@135464.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@135468.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@135462.4]
  assign regs_237_clock = clock; // @[:@135471.4]
  assign regs_237_reset = io_reset; // @[:@135472.4 RegFile.scala 76:16:@135479.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@135478.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@135482.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@135476.4]
  assign regs_238_clock = clock; // @[:@135485.4]
  assign regs_238_reset = io_reset; // @[:@135486.4 RegFile.scala 76:16:@135493.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@135492.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@135496.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@135490.4]
  assign regs_239_clock = clock; // @[:@135499.4]
  assign regs_239_reset = io_reset; // @[:@135500.4 RegFile.scala 76:16:@135507.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@135506.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@135510.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@135504.4]
  assign regs_240_clock = clock; // @[:@135513.4]
  assign regs_240_reset = io_reset; // @[:@135514.4 RegFile.scala 76:16:@135521.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@135520.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@135524.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@135518.4]
  assign regs_241_clock = clock; // @[:@135527.4]
  assign regs_241_reset = io_reset; // @[:@135528.4 RegFile.scala 76:16:@135535.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@135534.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@135538.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@135532.4]
  assign regs_242_clock = clock; // @[:@135541.4]
  assign regs_242_reset = io_reset; // @[:@135542.4 RegFile.scala 76:16:@135549.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@135548.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@135552.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@135546.4]
  assign regs_243_clock = clock; // @[:@135555.4]
  assign regs_243_reset = io_reset; // @[:@135556.4 RegFile.scala 76:16:@135563.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@135562.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@135566.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@135560.4]
  assign regs_244_clock = clock; // @[:@135569.4]
  assign regs_244_reset = io_reset; // @[:@135570.4 RegFile.scala 76:16:@135577.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@135576.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@135580.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@135574.4]
  assign regs_245_clock = clock; // @[:@135583.4]
  assign regs_245_reset = io_reset; // @[:@135584.4 RegFile.scala 76:16:@135591.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@135590.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@135594.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@135588.4]
  assign regs_246_clock = clock; // @[:@135597.4]
  assign regs_246_reset = io_reset; // @[:@135598.4 RegFile.scala 76:16:@135605.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@135604.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@135608.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@135602.4]
  assign regs_247_clock = clock; // @[:@135611.4]
  assign regs_247_reset = io_reset; // @[:@135612.4 RegFile.scala 76:16:@135619.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@135618.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@135622.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@135616.4]
  assign regs_248_clock = clock; // @[:@135625.4]
  assign regs_248_reset = io_reset; // @[:@135626.4 RegFile.scala 76:16:@135633.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@135632.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@135636.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@135630.4]
  assign regs_249_clock = clock; // @[:@135639.4]
  assign regs_249_reset = io_reset; // @[:@135640.4 RegFile.scala 76:16:@135647.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@135646.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@135650.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@135644.4]
  assign regs_250_clock = clock; // @[:@135653.4]
  assign regs_250_reset = io_reset; // @[:@135654.4 RegFile.scala 76:16:@135661.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@135660.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@135664.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@135658.4]
  assign regs_251_clock = clock; // @[:@135667.4]
  assign regs_251_reset = io_reset; // @[:@135668.4 RegFile.scala 76:16:@135675.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@135674.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@135678.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@135672.4]
  assign regs_252_clock = clock; // @[:@135681.4]
  assign regs_252_reset = io_reset; // @[:@135682.4 RegFile.scala 76:16:@135689.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@135688.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@135692.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@135686.4]
  assign regs_253_clock = clock; // @[:@135695.4]
  assign regs_253_reset = io_reset; // @[:@135696.4 RegFile.scala 76:16:@135703.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@135702.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@135706.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@135700.4]
  assign regs_254_clock = clock; // @[:@135709.4]
  assign regs_254_reset = io_reset; // @[:@135710.4 RegFile.scala 76:16:@135717.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@135716.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@135720.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@135714.4]
  assign regs_255_clock = clock; // @[:@135723.4]
  assign regs_255_reset = io_reset; // @[:@135724.4 RegFile.scala 76:16:@135731.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@135730.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@135734.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@135728.4]
  assign regs_256_clock = clock; // @[:@135737.4]
  assign regs_256_reset = io_reset; // @[:@135738.4 RegFile.scala 76:16:@135745.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@135744.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@135748.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@135742.4]
  assign regs_257_clock = clock; // @[:@135751.4]
  assign regs_257_reset = io_reset; // @[:@135752.4 RegFile.scala 76:16:@135759.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@135758.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@135762.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@135756.4]
  assign regs_258_clock = clock; // @[:@135765.4]
  assign regs_258_reset = io_reset; // @[:@135766.4 RegFile.scala 76:16:@135773.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@135772.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@135776.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@135770.4]
  assign regs_259_clock = clock; // @[:@135779.4]
  assign regs_259_reset = io_reset; // @[:@135780.4 RegFile.scala 76:16:@135787.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@135786.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@135790.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@135784.4]
  assign regs_260_clock = clock; // @[:@135793.4]
  assign regs_260_reset = io_reset; // @[:@135794.4 RegFile.scala 76:16:@135801.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@135800.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@135804.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@135798.4]
  assign regs_261_clock = clock; // @[:@135807.4]
  assign regs_261_reset = io_reset; // @[:@135808.4 RegFile.scala 76:16:@135815.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@135814.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@135818.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@135812.4]
  assign regs_262_clock = clock; // @[:@135821.4]
  assign regs_262_reset = io_reset; // @[:@135822.4 RegFile.scala 76:16:@135829.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@135828.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@135832.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@135826.4]
  assign regs_263_clock = clock; // @[:@135835.4]
  assign regs_263_reset = io_reset; // @[:@135836.4 RegFile.scala 76:16:@135843.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@135842.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@135846.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@135840.4]
  assign regs_264_clock = clock; // @[:@135849.4]
  assign regs_264_reset = io_reset; // @[:@135850.4 RegFile.scala 76:16:@135857.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@135856.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@135860.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@135854.4]
  assign regs_265_clock = clock; // @[:@135863.4]
  assign regs_265_reset = io_reset; // @[:@135864.4 RegFile.scala 76:16:@135871.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@135870.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@135874.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@135868.4]
  assign regs_266_clock = clock; // @[:@135877.4]
  assign regs_266_reset = io_reset; // @[:@135878.4 RegFile.scala 76:16:@135885.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@135884.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@135888.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@135882.4]
  assign regs_267_clock = clock; // @[:@135891.4]
  assign regs_267_reset = io_reset; // @[:@135892.4 RegFile.scala 76:16:@135899.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@135898.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@135902.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@135896.4]
  assign regs_268_clock = clock; // @[:@135905.4]
  assign regs_268_reset = io_reset; // @[:@135906.4 RegFile.scala 76:16:@135913.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@135912.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@135916.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@135910.4]
  assign regs_269_clock = clock; // @[:@135919.4]
  assign regs_269_reset = io_reset; // @[:@135920.4 RegFile.scala 76:16:@135927.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@135926.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@135930.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@135924.4]
  assign regs_270_clock = clock; // @[:@135933.4]
  assign regs_270_reset = io_reset; // @[:@135934.4 RegFile.scala 76:16:@135941.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@135940.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@135944.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@135938.4]
  assign regs_271_clock = clock; // @[:@135947.4]
  assign regs_271_reset = io_reset; // @[:@135948.4 RegFile.scala 76:16:@135955.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@135954.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@135958.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@135952.4]
  assign regs_272_clock = clock; // @[:@135961.4]
  assign regs_272_reset = io_reset; // @[:@135962.4 RegFile.scala 76:16:@135969.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@135968.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@135972.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@135966.4]
  assign regs_273_clock = clock; // @[:@135975.4]
  assign regs_273_reset = io_reset; // @[:@135976.4 RegFile.scala 76:16:@135983.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@135982.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@135986.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@135980.4]
  assign regs_274_clock = clock; // @[:@135989.4]
  assign regs_274_reset = io_reset; // @[:@135990.4 RegFile.scala 76:16:@135997.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@135996.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@136000.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@135994.4]
  assign regs_275_clock = clock; // @[:@136003.4]
  assign regs_275_reset = io_reset; // @[:@136004.4 RegFile.scala 76:16:@136011.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@136010.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@136014.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@136008.4]
  assign regs_276_clock = clock; // @[:@136017.4]
  assign regs_276_reset = io_reset; // @[:@136018.4 RegFile.scala 76:16:@136025.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@136024.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@136028.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@136022.4]
  assign regs_277_clock = clock; // @[:@136031.4]
  assign regs_277_reset = io_reset; // @[:@136032.4 RegFile.scala 76:16:@136039.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@136038.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@136042.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@136036.4]
  assign regs_278_clock = clock; // @[:@136045.4]
  assign regs_278_reset = io_reset; // @[:@136046.4 RegFile.scala 76:16:@136053.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@136052.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@136056.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@136050.4]
  assign regs_279_clock = clock; // @[:@136059.4]
  assign regs_279_reset = io_reset; // @[:@136060.4 RegFile.scala 76:16:@136067.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@136066.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@136070.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@136064.4]
  assign regs_280_clock = clock; // @[:@136073.4]
  assign regs_280_reset = io_reset; // @[:@136074.4 RegFile.scala 76:16:@136081.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@136080.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@136084.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@136078.4]
  assign regs_281_clock = clock; // @[:@136087.4]
  assign regs_281_reset = io_reset; // @[:@136088.4 RegFile.scala 76:16:@136095.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@136094.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@136098.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@136092.4]
  assign regs_282_clock = clock; // @[:@136101.4]
  assign regs_282_reset = io_reset; // @[:@136102.4 RegFile.scala 76:16:@136109.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@136108.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@136112.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@136106.4]
  assign regs_283_clock = clock; // @[:@136115.4]
  assign regs_283_reset = io_reset; // @[:@136116.4 RegFile.scala 76:16:@136123.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@136122.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@136126.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@136120.4]
  assign regs_284_clock = clock; // @[:@136129.4]
  assign regs_284_reset = io_reset; // @[:@136130.4 RegFile.scala 76:16:@136137.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@136136.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@136140.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@136134.4]
  assign regs_285_clock = clock; // @[:@136143.4]
  assign regs_285_reset = io_reset; // @[:@136144.4 RegFile.scala 76:16:@136151.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@136150.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@136154.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@136148.4]
  assign regs_286_clock = clock; // @[:@136157.4]
  assign regs_286_reset = io_reset; // @[:@136158.4 RegFile.scala 76:16:@136165.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@136164.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@136168.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@136162.4]
  assign regs_287_clock = clock; // @[:@136171.4]
  assign regs_287_reset = io_reset; // @[:@136172.4 RegFile.scala 76:16:@136179.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@136178.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@136182.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@136176.4]
  assign regs_288_clock = clock; // @[:@136185.4]
  assign regs_288_reset = io_reset; // @[:@136186.4 RegFile.scala 76:16:@136193.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@136192.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@136196.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@136190.4]
  assign regs_289_clock = clock; // @[:@136199.4]
  assign regs_289_reset = io_reset; // @[:@136200.4 RegFile.scala 76:16:@136207.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@136206.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@136210.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@136204.4]
  assign regs_290_clock = clock; // @[:@136213.4]
  assign regs_290_reset = io_reset; // @[:@136214.4 RegFile.scala 76:16:@136221.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@136220.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@136224.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@136218.4]
  assign regs_291_clock = clock; // @[:@136227.4]
  assign regs_291_reset = io_reset; // @[:@136228.4 RegFile.scala 76:16:@136235.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@136234.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@136238.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@136232.4]
  assign regs_292_clock = clock; // @[:@136241.4]
  assign regs_292_reset = io_reset; // @[:@136242.4 RegFile.scala 76:16:@136249.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@136248.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@136252.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@136246.4]
  assign regs_293_clock = clock; // @[:@136255.4]
  assign regs_293_reset = io_reset; // @[:@136256.4 RegFile.scala 76:16:@136263.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@136262.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@136266.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@136260.4]
  assign regs_294_clock = clock; // @[:@136269.4]
  assign regs_294_reset = io_reset; // @[:@136270.4 RegFile.scala 76:16:@136277.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@136276.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@136280.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@136274.4]
  assign regs_295_clock = clock; // @[:@136283.4]
  assign regs_295_reset = io_reset; // @[:@136284.4 RegFile.scala 76:16:@136291.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@136290.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@136294.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@136288.4]
  assign regs_296_clock = clock; // @[:@136297.4]
  assign regs_296_reset = io_reset; // @[:@136298.4 RegFile.scala 76:16:@136305.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@136304.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@136308.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@136302.4]
  assign regs_297_clock = clock; // @[:@136311.4]
  assign regs_297_reset = io_reset; // @[:@136312.4 RegFile.scala 76:16:@136319.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@136318.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@136322.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@136316.4]
  assign regs_298_clock = clock; // @[:@136325.4]
  assign regs_298_reset = io_reset; // @[:@136326.4 RegFile.scala 76:16:@136333.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@136332.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@136336.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@136330.4]
  assign regs_299_clock = clock; // @[:@136339.4]
  assign regs_299_reset = io_reset; // @[:@136340.4 RegFile.scala 76:16:@136347.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@136346.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@136350.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@136344.4]
  assign regs_300_clock = clock; // @[:@136353.4]
  assign regs_300_reset = io_reset; // @[:@136354.4 RegFile.scala 76:16:@136361.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@136360.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@136364.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@136358.4]
  assign regs_301_clock = clock; // @[:@136367.4]
  assign regs_301_reset = io_reset; // @[:@136368.4 RegFile.scala 76:16:@136375.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@136374.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@136378.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@136372.4]
  assign regs_302_clock = clock; // @[:@136381.4]
  assign regs_302_reset = io_reset; // @[:@136382.4 RegFile.scala 76:16:@136389.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@136388.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@136392.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@136386.4]
  assign regs_303_clock = clock; // @[:@136395.4]
  assign regs_303_reset = io_reset; // @[:@136396.4 RegFile.scala 76:16:@136403.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@136402.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@136406.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@136400.4]
  assign regs_304_clock = clock; // @[:@136409.4]
  assign regs_304_reset = io_reset; // @[:@136410.4 RegFile.scala 76:16:@136417.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@136416.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@136420.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@136414.4]
  assign regs_305_clock = clock; // @[:@136423.4]
  assign regs_305_reset = io_reset; // @[:@136424.4 RegFile.scala 76:16:@136431.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@136430.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@136434.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@136428.4]
  assign regs_306_clock = clock; // @[:@136437.4]
  assign regs_306_reset = io_reset; // @[:@136438.4 RegFile.scala 76:16:@136445.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@136444.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@136448.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@136442.4]
  assign regs_307_clock = clock; // @[:@136451.4]
  assign regs_307_reset = io_reset; // @[:@136452.4 RegFile.scala 76:16:@136459.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@136458.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@136462.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@136456.4]
  assign regs_308_clock = clock; // @[:@136465.4]
  assign regs_308_reset = io_reset; // @[:@136466.4 RegFile.scala 76:16:@136473.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@136472.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@136476.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@136470.4]
  assign regs_309_clock = clock; // @[:@136479.4]
  assign regs_309_reset = io_reset; // @[:@136480.4 RegFile.scala 76:16:@136487.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@136486.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@136490.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@136484.4]
  assign regs_310_clock = clock; // @[:@136493.4]
  assign regs_310_reset = io_reset; // @[:@136494.4 RegFile.scala 76:16:@136501.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@136500.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@136504.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@136498.4]
  assign regs_311_clock = clock; // @[:@136507.4]
  assign regs_311_reset = io_reset; // @[:@136508.4 RegFile.scala 76:16:@136515.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@136514.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@136518.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@136512.4]
  assign regs_312_clock = clock; // @[:@136521.4]
  assign regs_312_reset = io_reset; // @[:@136522.4 RegFile.scala 76:16:@136529.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@136528.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@136532.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@136526.4]
  assign regs_313_clock = clock; // @[:@136535.4]
  assign regs_313_reset = io_reset; // @[:@136536.4 RegFile.scala 76:16:@136543.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@136542.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@136546.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@136540.4]
  assign regs_314_clock = clock; // @[:@136549.4]
  assign regs_314_reset = io_reset; // @[:@136550.4 RegFile.scala 76:16:@136557.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@136556.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@136560.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@136554.4]
  assign regs_315_clock = clock; // @[:@136563.4]
  assign regs_315_reset = io_reset; // @[:@136564.4 RegFile.scala 76:16:@136571.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@136570.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@136574.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@136568.4]
  assign regs_316_clock = clock; // @[:@136577.4]
  assign regs_316_reset = io_reset; // @[:@136578.4 RegFile.scala 76:16:@136585.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@136584.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@136588.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@136582.4]
  assign regs_317_clock = clock; // @[:@136591.4]
  assign regs_317_reset = io_reset; // @[:@136592.4 RegFile.scala 76:16:@136599.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@136598.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@136602.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@136596.4]
  assign regs_318_clock = clock; // @[:@136605.4]
  assign regs_318_reset = io_reset; // @[:@136606.4 RegFile.scala 76:16:@136613.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@136612.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@136616.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@136610.4]
  assign regs_319_clock = clock; // @[:@136619.4]
  assign regs_319_reset = io_reset; // @[:@136620.4 RegFile.scala 76:16:@136627.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@136626.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@136630.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@136624.4]
  assign regs_320_clock = clock; // @[:@136633.4]
  assign regs_320_reset = io_reset; // @[:@136634.4 RegFile.scala 76:16:@136641.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@136640.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@136644.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@136638.4]
  assign regs_321_clock = clock; // @[:@136647.4]
  assign regs_321_reset = io_reset; // @[:@136648.4 RegFile.scala 76:16:@136655.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@136654.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@136658.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@136652.4]
  assign regs_322_clock = clock; // @[:@136661.4]
  assign regs_322_reset = io_reset; // @[:@136662.4 RegFile.scala 76:16:@136669.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@136668.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@136672.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@136666.4]
  assign regs_323_clock = clock; // @[:@136675.4]
  assign regs_323_reset = io_reset; // @[:@136676.4 RegFile.scala 76:16:@136683.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@136682.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@136686.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@136680.4]
  assign regs_324_clock = clock; // @[:@136689.4]
  assign regs_324_reset = io_reset; // @[:@136690.4 RegFile.scala 76:16:@136697.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@136696.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@136700.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@136694.4]
  assign regs_325_clock = clock; // @[:@136703.4]
  assign regs_325_reset = io_reset; // @[:@136704.4 RegFile.scala 76:16:@136711.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@136710.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@136714.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@136708.4]
  assign regs_326_clock = clock; // @[:@136717.4]
  assign regs_326_reset = io_reset; // @[:@136718.4 RegFile.scala 76:16:@136725.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@136724.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@136728.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@136722.4]
  assign regs_327_clock = clock; // @[:@136731.4]
  assign regs_327_reset = io_reset; // @[:@136732.4 RegFile.scala 76:16:@136739.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@136738.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@136742.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@136736.4]
  assign regs_328_clock = clock; // @[:@136745.4]
  assign regs_328_reset = io_reset; // @[:@136746.4 RegFile.scala 76:16:@136753.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@136752.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@136756.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@136750.4]
  assign regs_329_clock = clock; // @[:@136759.4]
  assign regs_329_reset = io_reset; // @[:@136760.4 RegFile.scala 76:16:@136767.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@136766.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@136770.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@136764.4]
  assign regs_330_clock = clock; // @[:@136773.4]
  assign regs_330_reset = io_reset; // @[:@136774.4 RegFile.scala 76:16:@136781.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@136780.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@136784.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@136778.4]
  assign regs_331_clock = clock; // @[:@136787.4]
  assign regs_331_reset = io_reset; // @[:@136788.4 RegFile.scala 76:16:@136795.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@136794.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@136798.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@136792.4]
  assign regs_332_clock = clock; // @[:@136801.4]
  assign regs_332_reset = io_reset; // @[:@136802.4 RegFile.scala 76:16:@136809.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@136808.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@136812.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@136806.4]
  assign regs_333_clock = clock; // @[:@136815.4]
  assign regs_333_reset = io_reset; // @[:@136816.4 RegFile.scala 76:16:@136823.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@136822.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@136826.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@136820.4]
  assign regs_334_clock = clock; // @[:@136829.4]
  assign regs_334_reset = io_reset; // @[:@136830.4 RegFile.scala 76:16:@136837.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@136836.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@136840.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@136834.4]
  assign regs_335_clock = clock; // @[:@136843.4]
  assign regs_335_reset = io_reset; // @[:@136844.4 RegFile.scala 76:16:@136851.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@136850.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@136854.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@136848.4]
  assign regs_336_clock = clock; // @[:@136857.4]
  assign regs_336_reset = io_reset; // @[:@136858.4 RegFile.scala 76:16:@136865.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@136864.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@136868.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@136862.4]
  assign regs_337_clock = clock; // @[:@136871.4]
  assign regs_337_reset = io_reset; // @[:@136872.4 RegFile.scala 76:16:@136879.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@136878.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@136882.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@136876.4]
  assign regs_338_clock = clock; // @[:@136885.4]
  assign regs_338_reset = io_reset; // @[:@136886.4 RegFile.scala 76:16:@136893.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@136892.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@136896.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@136890.4]
  assign regs_339_clock = clock; // @[:@136899.4]
  assign regs_339_reset = io_reset; // @[:@136900.4 RegFile.scala 76:16:@136907.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@136906.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@136910.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@136904.4]
  assign regs_340_clock = clock; // @[:@136913.4]
  assign regs_340_reset = io_reset; // @[:@136914.4 RegFile.scala 76:16:@136921.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@136920.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@136924.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@136918.4]
  assign regs_341_clock = clock; // @[:@136927.4]
  assign regs_341_reset = io_reset; // @[:@136928.4 RegFile.scala 76:16:@136935.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@136934.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@136938.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@136932.4]
  assign regs_342_clock = clock; // @[:@136941.4]
  assign regs_342_reset = io_reset; // @[:@136942.4 RegFile.scala 76:16:@136949.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@136948.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@136952.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@136946.4]
  assign regs_343_clock = clock; // @[:@136955.4]
  assign regs_343_reset = io_reset; // @[:@136956.4 RegFile.scala 76:16:@136963.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@136962.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@136966.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@136960.4]
  assign regs_344_clock = clock; // @[:@136969.4]
  assign regs_344_reset = io_reset; // @[:@136970.4 RegFile.scala 76:16:@136977.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@136976.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@136980.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@136974.4]
  assign regs_345_clock = clock; // @[:@136983.4]
  assign regs_345_reset = io_reset; // @[:@136984.4 RegFile.scala 76:16:@136991.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@136990.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@136994.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@136988.4]
  assign regs_346_clock = clock; // @[:@136997.4]
  assign regs_346_reset = io_reset; // @[:@136998.4 RegFile.scala 76:16:@137005.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@137004.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@137008.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@137002.4]
  assign regs_347_clock = clock; // @[:@137011.4]
  assign regs_347_reset = io_reset; // @[:@137012.4 RegFile.scala 76:16:@137019.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@137018.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@137022.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@137016.4]
  assign regs_348_clock = clock; // @[:@137025.4]
  assign regs_348_reset = io_reset; // @[:@137026.4 RegFile.scala 76:16:@137033.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@137032.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@137036.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@137030.4]
  assign regs_349_clock = clock; // @[:@137039.4]
  assign regs_349_reset = io_reset; // @[:@137040.4 RegFile.scala 76:16:@137047.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@137046.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@137050.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@137044.4]
  assign regs_350_clock = clock; // @[:@137053.4]
  assign regs_350_reset = io_reset; // @[:@137054.4 RegFile.scala 76:16:@137061.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@137060.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@137064.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@137058.4]
  assign regs_351_clock = clock; // @[:@137067.4]
  assign regs_351_reset = io_reset; // @[:@137068.4 RegFile.scala 76:16:@137075.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@137074.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@137078.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@137072.4]
  assign regs_352_clock = clock; // @[:@137081.4]
  assign regs_352_reset = io_reset; // @[:@137082.4 RegFile.scala 76:16:@137089.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@137088.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@137092.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@137086.4]
  assign regs_353_clock = clock; // @[:@137095.4]
  assign regs_353_reset = io_reset; // @[:@137096.4 RegFile.scala 76:16:@137103.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@137102.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@137106.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@137100.4]
  assign regs_354_clock = clock; // @[:@137109.4]
  assign regs_354_reset = io_reset; // @[:@137110.4 RegFile.scala 76:16:@137117.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@137116.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@137120.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@137114.4]
  assign regs_355_clock = clock; // @[:@137123.4]
  assign regs_355_reset = io_reset; // @[:@137124.4 RegFile.scala 76:16:@137131.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@137130.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@137134.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@137128.4]
  assign regs_356_clock = clock; // @[:@137137.4]
  assign regs_356_reset = io_reset; // @[:@137138.4 RegFile.scala 76:16:@137145.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@137144.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@137148.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@137142.4]
  assign regs_357_clock = clock; // @[:@137151.4]
  assign regs_357_reset = io_reset; // @[:@137152.4 RegFile.scala 76:16:@137159.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@137158.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@137162.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@137156.4]
  assign regs_358_clock = clock; // @[:@137165.4]
  assign regs_358_reset = io_reset; // @[:@137166.4 RegFile.scala 76:16:@137173.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@137172.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@137176.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@137170.4]
  assign regs_359_clock = clock; // @[:@137179.4]
  assign regs_359_reset = io_reset; // @[:@137180.4 RegFile.scala 76:16:@137187.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@137186.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@137190.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@137184.4]
  assign regs_360_clock = clock; // @[:@137193.4]
  assign regs_360_reset = io_reset; // @[:@137194.4 RegFile.scala 76:16:@137201.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@137200.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@137204.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@137198.4]
  assign regs_361_clock = clock; // @[:@137207.4]
  assign regs_361_reset = io_reset; // @[:@137208.4 RegFile.scala 76:16:@137215.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@137214.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@137218.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@137212.4]
  assign regs_362_clock = clock; // @[:@137221.4]
  assign regs_362_reset = io_reset; // @[:@137222.4 RegFile.scala 76:16:@137229.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@137228.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@137232.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@137226.4]
  assign regs_363_clock = clock; // @[:@137235.4]
  assign regs_363_reset = io_reset; // @[:@137236.4 RegFile.scala 76:16:@137243.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@137242.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@137246.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@137240.4]
  assign regs_364_clock = clock; // @[:@137249.4]
  assign regs_364_reset = io_reset; // @[:@137250.4 RegFile.scala 76:16:@137257.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@137256.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@137260.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@137254.4]
  assign regs_365_clock = clock; // @[:@137263.4]
  assign regs_365_reset = io_reset; // @[:@137264.4 RegFile.scala 76:16:@137271.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@137270.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@137274.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@137268.4]
  assign regs_366_clock = clock; // @[:@137277.4]
  assign regs_366_reset = io_reset; // @[:@137278.4 RegFile.scala 76:16:@137285.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@137284.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@137288.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@137282.4]
  assign regs_367_clock = clock; // @[:@137291.4]
  assign regs_367_reset = io_reset; // @[:@137292.4 RegFile.scala 76:16:@137299.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@137298.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@137302.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@137296.4]
  assign regs_368_clock = clock; // @[:@137305.4]
  assign regs_368_reset = io_reset; // @[:@137306.4 RegFile.scala 76:16:@137313.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@137312.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@137316.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@137310.4]
  assign regs_369_clock = clock; // @[:@137319.4]
  assign regs_369_reset = io_reset; // @[:@137320.4 RegFile.scala 76:16:@137327.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@137326.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@137330.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@137324.4]
  assign regs_370_clock = clock; // @[:@137333.4]
  assign regs_370_reset = io_reset; // @[:@137334.4 RegFile.scala 76:16:@137341.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@137340.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@137344.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@137338.4]
  assign regs_371_clock = clock; // @[:@137347.4]
  assign regs_371_reset = io_reset; // @[:@137348.4 RegFile.scala 76:16:@137355.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@137354.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@137358.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@137352.4]
  assign regs_372_clock = clock; // @[:@137361.4]
  assign regs_372_reset = io_reset; // @[:@137362.4 RegFile.scala 76:16:@137369.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@137368.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@137372.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@137366.4]
  assign regs_373_clock = clock; // @[:@137375.4]
  assign regs_373_reset = io_reset; // @[:@137376.4 RegFile.scala 76:16:@137383.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@137382.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@137386.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@137380.4]
  assign regs_374_clock = clock; // @[:@137389.4]
  assign regs_374_reset = io_reset; // @[:@137390.4 RegFile.scala 76:16:@137397.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@137396.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@137400.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@137394.4]
  assign regs_375_clock = clock; // @[:@137403.4]
  assign regs_375_reset = io_reset; // @[:@137404.4 RegFile.scala 76:16:@137411.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@137410.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@137414.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@137408.4]
  assign regs_376_clock = clock; // @[:@137417.4]
  assign regs_376_reset = io_reset; // @[:@137418.4 RegFile.scala 76:16:@137425.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@137424.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@137428.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@137422.4]
  assign regs_377_clock = clock; // @[:@137431.4]
  assign regs_377_reset = io_reset; // @[:@137432.4 RegFile.scala 76:16:@137439.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@137438.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@137442.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@137436.4]
  assign regs_378_clock = clock; // @[:@137445.4]
  assign regs_378_reset = io_reset; // @[:@137446.4 RegFile.scala 76:16:@137453.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@137452.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@137456.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@137450.4]
  assign regs_379_clock = clock; // @[:@137459.4]
  assign regs_379_reset = io_reset; // @[:@137460.4 RegFile.scala 76:16:@137467.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@137466.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@137470.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@137464.4]
  assign regs_380_clock = clock; // @[:@137473.4]
  assign regs_380_reset = io_reset; // @[:@137474.4 RegFile.scala 76:16:@137481.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@137480.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@137484.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@137478.4]
  assign regs_381_clock = clock; // @[:@137487.4]
  assign regs_381_reset = io_reset; // @[:@137488.4 RegFile.scala 76:16:@137495.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@137494.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@137498.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@137492.4]
  assign regs_382_clock = clock; // @[:@137501.4]
  assign regs_382_reset = io_reset; // @[:@137502.4 RegFile.scala 76:16:@137509.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@137508.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@137512.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@137506.4]
  assign regs_383_clock = clock; // @[:@137515.4]
  assign regs_383_reset = io_reset; // @[:@137516.4 RegFile.scala 76:16:@137523.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@137522.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@137526.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@137520.4]
  assign regs_384_clock = clock; // @[:@137529.4]
  assign regs_384_reset = io_reset; // @[:@137530.4 RegFile.scala 76:16:@137537.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@137536.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@137540.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@137534.4]
  assign regs_385_clock = clock; // @[:@137543.4]
  assign regs_385_reset = io_reset; // @[:@137544.4 RegFile.scala 76:16:@137551.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@137550.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@137554.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@137548.4]
  assign regs_386_clock = clock; // @[:@137557.4]
  assign regs_386_reset = io_reset; // @[:@137558.4 RegFile.scala 76:16:@137565.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@137564.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@137568.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@137562.4]
  assign regs_387_clock = clock; // @[:@137571.4]
  assign regs_387_reset = io_reset; // @[:@137572.4 RegFile.scala 76:16:@137579.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@137578.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@137582.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@137576.4]
  assign regs_388_clock = clock; // @[:@137585.4]
  assign regs_388_reset = io_reset; // @[:@137586.4 RegFile.scala 76:16:@137593.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@137592.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@137596.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@137590.4]
  assign regs_389_clock = clock; // @[:@137599.4]
  assign regs_389_reset = io_reset; // @[:@137600.4 RegFile.scala 76:16:@137607.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@137606.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@137610.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@137604.4]
  assign regs_390_clock = clock; // @[:@137613.4]
  assign regs_390_reset = io_reset; // @[:@137614.4 RegFile.scala 76:16:@137621.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@137620.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@137624.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@137618.4]
  assign regs_391_clock = clock; // @[:@137627.4]
  assign regs_391_reset = io_reset; // @[:@137628.4 RegFile.scala 76:16:@137635.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@137634.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@137638.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@137632.4]
  assign regs_392_clock = clock; // @[:@137641.4]
  assign regs_392_reset = io_reset; // @[:@137642.4 RegFile.scala 76:16:@137649.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@137648.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@137652.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@137646.4]
  assign regs_393_clock = clock; // @[:@137655.4]
  assign regs_393_reset = io_reset; // @[:@137656.4 RegFile.scala 76:16:@137663.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@137662.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@137666.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@137660.4]
  assign regs_394_clock = clock; // @[:@137669.4]
  assign regs_394_reset = io_reset; // @[:@137670.4 RegFile.scala 76:16:@137677.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@137676.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@137680.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@137674.4]
  assign regs_395_clock = clock; // @[:@137683.4]
  assign regs_395_reset = io_reset; // @[:@137684.4 RegFile.scala 76:16:@137691.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@137690.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@137694.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@137688.4]
  assign regs_396_clock = clock; // @[:@137697.4]
  assign regs_396_reset = io_reset; // @[:@137698.4 RegFile.scala 76:16:@137705.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@137704.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@137708.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@137702.4]
  assign regs_397_clock = clock; // @[:@137711.4]
  assign regs_397_reset = io_reset; // @[:@137712.4 RegFile.scala 76:16:@137719.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@137718.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@137722.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@137716.4]
  assign regs_398_clock = clock; // @[:@137725.4]
  assign regs_398_reset = io_reset; // @[:@137726.4 RegFile.scala 76:16:@137733.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@137732.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@137736.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@137730.4]
  assign regs_399_clock = clock; // @[:@137739.4]
  assign regs_399_reset = io_reset; // @[:@137740.4 RegFile.scala 76:16:@137747.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@137746.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@137750.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@137744.4]
  assign regs_400_clock = clock; // @[:@137753.4]
  assign regs_400_reset = io_reset; // @[:@137754.4 RegFile.scala 76:16:@137761.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@137760.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@137764.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@137758.4]
  assign regs_401_clock = clock; // @[:@137767.4]
  assign regs_401_reset = io_reset; // @[:@137768.4 RegFile.scala 76:16:@137775.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@137774.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@137778.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@137772.4]
  assign regs_402_clock = clock; // @[:@137781.4]
  assign regs_402_reset = io_reset; // @[:@137782.4 RegFile.scala 76:16:@137789.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@137788.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@137792.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@137786.4]
  assign regs_403_clock = clock; // @[:@137795.4]
  assign regs_403_reset = io_reset; // @[:@137796.4 RegFile.scala 76:16:@137803.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@137802.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@137806.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@137800.4]
  assign regs_404_clock = clock; // @[:@137809.4]
  assign regs_404_reset = io_reset; // @[:@137810.4 RegFile.scala 76:16:@137817.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@137816.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@137820.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@137814.4]
  assign regs_405_clock = clock; // @[:@137823.4]
  assign regs_405_reset = io_reset; // @[:@137824.4 RegFile.scala 76:16:@137831.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@137830.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@137834.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@137828.4]
  assign regs_406_clock = clock; // @[:@137837.4]
  assign regs_406_reset = io_reset; // @[:@137838.4 RegFile.scala 76:16:@137845.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@137844.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@137848.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@137842.4]
  assign regs_407_clock = clock; // @[:@137851.4]
  assign regs_407_reset = io_reset; // @[:@137852.4 RegFile.scala 76:16:@137859.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@137858.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@137862.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@137856.4]
  assign regs_408_clock = clock; // @[:@137865.4]
  assign regs_408_reset = io_reset; // @[:@137866.4 RegFile.scala 76:16:@137873.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@137872.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@137876.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@137870.4]
  assign regs_409_clock = clock; // @[:@137879.4]
  assign regs_409_reset = io_reset; // @[:@137880.4 RegFile.scala 76:16:@137887.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@137886.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@137890.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@137884.4]
  assign regs_410_clock = clock; // @[:@137893.4]
  assign regs_410_reset = io_reset; // @[:@137894.4 RegFile.scala 76:16:@137901.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@137900.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@137904.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@137898.4]
  assign regs_411_clock = clock; // @[:@137907.4]
  assign regs_411_reset = io_reset; // @[:@137908.4 RegFile.scala 76:16:@137915.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@137914.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@137918.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@137912.4]
  assign regs_412_clock = clock; // @[:@137921.4]
  assign regs_412_reset = io_reset; // @[:@137922.4 RegFile.scala 76:16:@137929.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@137928.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@137932.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@137926.4]
  assign regs_413_clock = clock; // @[:@137935.4]
  assign regs_413_reset = io_reset; // @[:@137936.4 RegFile.scala 76:16:@137943.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@137942.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@137946.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@137940.4]
  assign regs_414_clock = clock; // @[:@137949.4]
  assign regs_414_reset = io_reset; // @[:@137950.4 RegFile.scala 76:16:@137957.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@137956.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@137960.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@137954.4]
  assign regs_415_clock = clock; // @[:@137963.4]
  assign regs_415_reset = io_reset; // @[:@137964.4 RegFile.scala 76:16:@137971.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@137970.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@137974.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@137968.4]
  assign regs_416_clock = clock; // @[:@137977.4]
  assign regs_416_reset = io_reset; // @[:@137978.4 RegFile.scala 76:16:@137985.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@137984.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@137988.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@137982.4]
  assign regs_417_clock = clock; // @[:@137991.4]
  assign regs_417_reset = io_reset; // @[:@137992.4 RegFile.scala 76:16:@137999.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@137998.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@138002.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@137996.4]
  assign regs_418_clock = clock; // @[:@138005.4]
  assign regs_418_reset = io_reset; // @[:@138006.4 RegFile.scala 76:16:@138013.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@138012.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@138016.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@138010.4]
  assign regs_419_clock = clock; // @[:@138019.4]
  assign regs_419_reset = io_reset; // @[:@138020.4 RegFile.scala 76:16:@138027.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@138026.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@138030.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@138024.4]
  assign regs_420_clock = clock; // @[:@138033.4]
  assign regs_420_reset = io_reset; // @[:@138034.4 RegFile.scala 76:16:@138041.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@138040.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@138044.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@138038.4]
  assign regs_421_clock = clock; // @[:@138047.4]
  assign regs_421_reset = io_reset; // @[:@138048.4 RegFile.scala 76:16:@138055.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@138054.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@138058.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@138052.4]
  assign regs_422_clock = clock; // @[:@138061.4]
  assign regs_422_reset = io_reset; // @[:@138062.4 RegFile.scala 76:16:@138069.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@138068.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@138072.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@138066.4]
  assign regs_423_clock = clock; // @[:@138075.4]
  assign regs_423_reset = io_reset; // @[:@138076.4 RegFile.scala 76:16:@138083.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@138082.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@138086.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@138080.4]
  assign regs_424_clock = clock; // @[:@138089.4]
  assign regs_424_reset = io_reset; // @[:@138090.4 RegFile.scala 76:16:@138097.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@138096.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@138100.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@138094.4]
  assign regs_425_clock = clock; // @[:@138103.4]
  assign regs_425_reset = io_reset; // @[:@138104.4 RegFile.scala 76:16:@138111.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@138110.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@138114.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@138108.4]
  assign regs_426_clock = clock; // @[:@138117.4]
  assign regs_426_reset = io_reset; // @[:@138118.4 RegFile.scala 76:16:@138125.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@138124.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@138128.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@138122.4]
  assign regs_427_clock = clock; // @[:@138131.4]
  assign regs_427_reset = io_reset; // @[:@138132.4 RegFile.scala 76:16:@138139.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@138138.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@138142.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@138136.4]
  assign regs_428_clock = clock; // @[:@138145.4]
  assign regs_428_reset = io_reset; // @[:@138146.4 RegFile.scala 76:16:@138153.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@138152.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@138156.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@138150.4]
  assign regs_429_clock = clock; // @[:@138159.4]
  assign regs_429_reset = io_reset; // @[:@138160.4 RegFile.scala 76:16:@138167.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@138166.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@138170.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@138164.4]
  assign regs_430_clock = clock; // @[:@138173.4]
  assign regs_430_reset = io_reset; // @[:@138174.4 RegFile.scala 76:16:@138181.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@138180.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@138184.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@138178.4]
  assign regs_431_clock = clock; // @[:@138187.4]
  assign regs_431_reset = io_reset; // @[:@138188.4 RegFile.scala 76:16:@138195.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@138194.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@138198.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@138192.4]
  assign regs_432_clock = clock; // @[:@138201.4]
  assign regs_432_reset = io_reset; // @[:@138202.4 RegFile.scala 76:16:@138209.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@138208.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@138212.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@138206.4]
  assign regs_433_clock = clock; // @[:@138215.4]
  assign regs_433_reset = io_reset; // @[:@138216.4 RegFile.scala 76:16:@138223.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@138222.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@138226.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@138220.4]
  assign regs_434_clock = clock; // @[:@138229.4]
  assign regs_434_reset = io_reset; // @[:@138230.4 RegFile.scala 76:16:@138237.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@138236.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@138240.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@138234.4]
  assign regs_435_clock = clock; // @[:@138243.4]
  assign regs_435_reset = io_reset; // @[:@138244.4 RegFile.scala 76:16:@138251.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@138250.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@138254.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@138248.4]
  assign regs_436_clock = clock; // @[:@138257.4]
  assign regs_436_reset = io_reset; // @[:@138258.4 RegFile.scala 76:16:@138265.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@138264.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@138268.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@138262.4]
  assign regs_437_clock = clock; // @[:@138271.4]
  assign regs_437_reset = io_reset; // @[:@138272.4 RegFile.scala 76:16:@138279.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@138278.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@138282.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@138276.4]
  assign regs_438_clock = clock; // @[:@138285.4]
  assign regs_438_reset = io_reset; // @[:@138286.4 RegFile.scala 76:16:@138293.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@138292.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@138296.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@138290.4]
  assign regs_439_clock = clock; // @[:@138299.4]
  assign regs_439_reset = io_reset; // @[:@138300.4 RegFile.scala 76:16:@138307.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@138306.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@138310.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@138304.4]
  assign regs_440_clock = clock; // @[:@138313.4]
  assign regs_440_reset = io_reset; // @[:@138314.4 RegFile.scala 76:16:@138321.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@138320.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@138324.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@138318.4]
  assign regs_441_clock = clock; // @[:@138327.4]
  assign regs_441_reset = io_reset; // @[:@138328.4 RegFile.scala 76:16:@138335.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@138334.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@138338.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@138332.4]
  assign regs_442_clock = clock; // @[:@138341.4]
  assign regs_442_reset = io_reset; // @[:@138342.4 RegFile.scala 76:16:@138349.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@138348.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@138352.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@138346.4]
  assign regs_443_clock = clock; // @[:@138355.4]
  assign regs_443_reset = io_reset; // @[:@138356.4 RegFile.scala 76:16:@138363.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@138362.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@138366.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@138360.4]
  assign regs_444_clock = clock; // @[:@138369.4]
  assign regs_444_reset = io_reset; // @[:@138370.4 RegFile.scala 76:16:@138377.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@138376.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@138380.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@138374.4]
  assign regs_445_clock = clock; // @[:@138383.4]
  assign regs_445_reset = io_reset; // @[:@138384.4 RegFile.scala 76:16:@138391.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@138390.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@138394.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@138388.4]
  assign regs_446_clock = clock; // @[:@138397.4]
  assign regs_446_reset = io_reset; // @[:@138398.4 RegFile.scala 76:16:@138405.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@138404.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@138408.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@138402.4]
  assign regs_447_clock = clock; // @[:@138411.4]
  assign regs_447_reset = io_reset; // @[:@138412.4 RegFile.scala 76:16:@138419.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@138418.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@138422.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@138416.4]
  assign regs_448_clock = clock; // @[:@138425.4]
  assign regs_448_reset = io_reset; // @[:@138426.4 RegFile.scala 76:16:@138433.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@138432.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@138436.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@138430.4]
  assign regs_449_clock = clock; // @[:@138439.4]
  assign regs_449_reset = io_reset; // @[:@138440.4 RegFile.scala 76:16:@138447.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@138446.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@138450.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@138444.4]
  assign regs_450_clock = clock; // @[:@138453.4]
  assign regs_450_reset = io_reset; // @[:@138454.4 RegFile.scala 76:16:@138461.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@138460.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@138464.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@138458.4]
  assign regs_451_clock = clock; // @[:@138467.4]
  assign regs_451_reset = io_reset; // @[:@138468.4 RegFile.scala 76:16:@138475.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@138474.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@138478.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@138472.4]
  assign regs_452_clock = clock; // @[:@138481.4]
  assign regs_452_reset = io_reset; // @[:@138482.4 RegFile.scala 76:16:@138489.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@138488.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@138492.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@138486.4]
  assign regs_453_clock = clock; // @[:@138495.4]
  assign regs_453_reset = io_reset; // @[:@138496.4 RegFile.scala 76:16:@138503.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@138502.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@138506.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@138500.4]
  assign regs_454_clock = clock; // @[:@138509.4]
  assign regs_454_reset = io_reset; // @[:@138510.4 RegFile.scala 76:16:@138517.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@138516.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@138520.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@138514.4]
  assign regs_455_clock = clock; // @[:@138523.4]
  assign regs_455_reset = io_reset; // @[:@138524.4 RegFile.scala 76:16:@138531.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@138530.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@138534.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@138528.4]
  assign regs_456_clock = clock; // @[:@138537.4]
  assign regs_456_reset = io_reset; // @[:@138538.4 RegFile.scala 76:16:@138545.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@138544.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@138548.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@138542.4]
  assign regs_457_clock = clock; // @[:@138551.4]
  assign regs_457_reset = io_reset; // @[:@138552.4 RegFile.scala 76:16:@138559.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@138558.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@138562.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@138556.4]
  assign regs_458_clock = clock; // @[:@138565.4]
  assign regs_458_reset = io_reset; // @[:@138566.4 RegFile.scala 76:16:@138573.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@138572.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@138576.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@138570.4]
  assign regs_459_clock = clock; // @[:@138579.4]
  assign regs_459_reset = io_reset; // @[:@138580.4 RegFile.scala 76:16:@138587.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@138586.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@138590.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@138584.4]
  assign regs_460_clock = clock; // @[:@138593.4]
  assign regs_460_reset = io_reset; // @[:@138594.4 RegFile.scala 76:16:@138601.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@138600.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@138604.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@138598.4]
  assign regs_461_clock = clock; // @[:@138607.4]
  assign regs_461_reset = io_reset; // @[:@138608.4 RegFile.scala 76:16:@138615.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@138614.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@138618.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@138612.4]
  assign regs_462_clock = clock; // @[:@138621.4]
  assign regs_462_reset = io_reset; // @[:@138622.4 RegFile.scala 76:16:@138629.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@138628.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@138632.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@138626.4]
  assign regs_463_clock = clock; // @[:@138635.4]
  assign regs_463_reset = io_reset; // @[:@138636.4 RegFile.scala 76:16:@138643.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@138642.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@138646.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@138640.4]
  assign regs_464_clock = clock; // @[:@138649.4]
  assign regs_464_reset = io_reset; // @[:@138650.4 RegFile.scala 76:16:@138657.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@138656.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@138660.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@138654.4]
  assign regs_465_clock = clock; // @[:@138663.4]
  assign regs_465_reset = io_reset; // @[:@138664.4 RegFile.scala 76:16:@138671.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@138670.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@138674.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@138668.4]
  assign regs_466_clock = clock; // @[:@138677.4]
  assign regs_466_reset = io_reset; // @[:@138678.4 RegFile.scala 76:16:@138685.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@138684.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@138688.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@138682.4]
  assign regs_467_clock = clock; // @[:@138691.4]
  assign regs_467_reset = io_reset; // @[:@138692.4 RegFile.scala 76:16:@138699.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@138698.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@138702.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@138696.4]
  assign regs_468_clock = clock; // @[:@138705.4]
  assign regs_468_reset = io_reset; // @[:@138706.4 RegFile.scala 76:16:@138713.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@138712.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@138716.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@138710.4]
  assign regs_469_clock = clock; // @[:@138719.4]
  assign regs_469_reset = io_reset; // @[:@138720.4 RegFile.scala 76:16:@138727.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@138726.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@138730.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@138724.4]
  assign regs_470_clock = clock; // @[:@138733.4]
  assign regs_470_reset = io_reset; // @[:@138734.4 RegFile.scala 76:16:@138741.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@138740.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@138744.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@138738.4]
  assign regs_471_clock = clock; // @[:@138747.4]
  assign regs_471_reset = io_reset; // @[:@138748.4 RegFile.scala 76:16:@138755.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@138754.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@138758.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@138752.4]
  assign regs_472_clock = clock; // @[:@138761.4]
  assign regs_472_reset = io_reset; // @[:@138762.4 RegFile.scala 76:16:@138769.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@138768.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@138772.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@138766.4]
  assign regs_473_clock = clock; // @[:@138775.4]
  assign regs_473_reset = io_reset; // @[:@138776.4 RegFile.scala 76:16:@138783.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@138782.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@138786.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@138780.4]
  assign regs_474_clock = clock; // @[:@138789.4]
  assign regs_474_reset = io_reset; // @[:@138790.4 RegFile.scala 76:16:@138797.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@138796.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@138800.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@138794.4]
  assign regs_475_clock = clock; // @[:@138803.4]
  assign regs_475_reset = io_reset; // @[:@138804.4 RegFile.scala 76:16:@138811.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@138810.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@138814.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@138808.4]
  assign regs_476_clock = clock; // @[:@138817.4]
  assign regs_476_reset = io_reset; // @[:@138818.4 RegFile.scala 76:16:@138825.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@138824.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@138828.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@138822.4]
  assign regs_477_clock = clock; // @[:@138831.4]
  assign regs_477_reset = io_reset; // @[:@138832.4 RegFile.scala 76:16:@138839.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@138838.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@138842.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@138836.4]
  assign regs_478_clock = clock; // @[:@138845.4]
  assign regs_478_reset = io_reset; // @[:@138846.4 RegFile.scala 76:16:@138853.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@138852.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@138856.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@138850.4]
  assign regs_479_clock = clock; // @[:@138859.4]
  assign regs_479_reset = io_reset; // @[:@138860.4 RegFile.scala 76:16:@138867.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@138866.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@138870.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@138864.4]
  assign regs_480_clock = clock; // @[:@138873.4]
  assign regs_480_reset = io_reset; // @[:@138874.4 RegFile.scala 76:16:@138881.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@138880.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@138884.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@138878.4]
  assign regs_481_clock = clock; // @[:@138887.4]
  assign regs_481_reset = io_reset; // @[:@138888.4 RegFile.scala 76:16:@138895.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@138894.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@138898.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@138892.4]
  assign regs_482_clock = clock; // @[:@138901.4]
  assign regs_482_reset = io_reset; // @[:@138902.4 RegFile.scala 76:16:@138909.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@138908.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@138912.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@138906.4]
  assign regs_483_clock = clock; // @[:@138915.4]
  assign regs_483_reset = io_reset; // @[:@138916.4 RegFile.scala 76:16:@138923.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@138922.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@138926.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@138920.4]
  assign regs_484_clock = clock; // @[:@138929.4]
  assign regs_484_reset = io_reset; // @[:@138930.4 RegFile.scala 76:16:@138937.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@138936.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@138940.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@138934.4]
  assign regs_485_clock = clock; // @[:@138943.4]
  assign regs_485_reset = io_reset; // @[:@138944.4 RegFile.scala 76:16:@138951.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@138950.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@138954.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@138948.4]
  assign regs_486_clock = clock; // @[:@138957.4]
  assign regs_486_reset = io_reset; // @[:@138958.4 RegFile.scala 76:16:@138965.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@138964.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@138968.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@138962.4]
  assign regs_487_clock = clock; // @[:@138971.4]
  assign regs_487_reset = io_reset; // @[:@138972.4 RegFile.scala 76:16:@138979.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@138978.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@138982.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@138976.4]
  assign regs_488_clock = clock; // @[:@138985.4]
  assign regs_488_reset = io_reset; // @[:@138986.4 RegFile.scala 76:16:@138993.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@138992.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@138996.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@138990.4]
  assign regs_489_clock = clock; // @[:@138999.4]
  assign regs_489_reset = io_reset; // @[:@139000.4 RegFile.scala 76:16:@139007.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@139006.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@139010.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@139004.4]
  assign regs_490_clock = clock; // @[:@139013.4]
  assign regs_490_reset = io_reset; // @[:@139014.4 RegFile.scala 76:16:@139021.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@139020.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@139024.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@139018.4]
  assign regs_491_clock = clock; // @[:@139027.4]
  assign regs_491_reset = io_reset; // @[:@139028.4 RegFile.scala 76:16:@139035.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@139034.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@139038.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@139032.4]
  assign regs_492_clock = clock; // @[:@139041.4]
  assign regs_492_reset = io_reset; // @[:@139042.4 RegFile.scala 76:16:@139049.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@139048.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@139052.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@139046.4]
  assign regs_493_clock = clock; // @[:@139055.4]
  assign regs_493_reset = io_reset; // @[:@139056.4 RegFile.scala 76:16:@139063.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@139062.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@139066.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@139060.4]
  assign regs_494_clock = clock; // @[:@139069.4]
  assign regs_494_reset = io_reset; // @[:@139070.4 RegFile.scala 76:16:@139077.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@139076.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@139080.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@139074.4]
  assign regs_495_clock = clock; // @[:@139083.4]
  assign regs_495_reset = io_reset; // @[:@139084.4 RegFile.scala 76:16:@139091.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@139090.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@139094.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@139088.4]
  assign regs_496_clock = clock; // @[:@139097.4]
  assign regs_496_reset = io_reset; // @[:@139098.4 RegFile.scala 76:16:@139105.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@139104.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@139108.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@139102.4]
  assign regs_497_clock = clock; // @[:@139111.4]
  assign regs_497_reset = io_reset; // @[:@139112.4 RegFile.scala 76:16:@139119.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@139118.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@139122.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@139116.4]
  assign regs_498_clock = clock; // @[:@139125.4]
  assign regs_498_reset = io_reset; // @[:@139126.4 RegFile.scala 76:16:@139133.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@139132.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@139136.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@139130.4]
  assign regs_499_clock = clock; // @[:@139139.4]
  assign regs_499_reset = io_reset; // @[:@139140.4 RegFile.scala 76:16:@139147.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@139146.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@139150.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@139144.4]
  assign regs_500_clock = clock; // @[:@139153.4]
  assign regs_500_reset = io_reset; // @[:@139154.4 RegFile.scala 76:16:@139161.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@139160.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@139164.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@139158.4]
  assign regs_501_clock = clock; // @[:@139167.4]
  assign regs_501_reset = io_reset; // @[:@139168.4 RegFile.scala 76:16:@139175.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@139174.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@139178.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@139172.4]
  assign regs_502_clock = clock; // @[:@139181.4]
  assign regs_502_reset = io_reset; // @[:@139182.4 RegFile.scala 76:16:@139189.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@139188.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@139192.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@139186.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@139701.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@139702.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@139703.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@139704.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@139705.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@139706.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@139707.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@139708.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@139709.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@139710.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@139711.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@139712.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@139713.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@139714.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@139715.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@139716.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@139717.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@139718.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@139719.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@139720.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@139721.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@139722.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@139723.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@139724.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@139725.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@139726.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@139727.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@139728.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@139729.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@139730.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@139731.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@139732.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@139733.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@139734.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@139735.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@139736.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@139737.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@139738.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@139739.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@139740.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@139741.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@139742.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@139743.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@139744.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@139745.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@139746.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@139747.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@139748.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@139749.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@139750.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@139751.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@139752.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@139753.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@139754.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@139755.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@139756.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@139757.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@139758.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@139759.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@139760.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@139761.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@139762.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@139763.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@139764.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@139765.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@139766.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@139767.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@139768.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@139769.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@139770.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@139771.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@139772.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@139773.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@139774.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@139775.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@139776.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@139777.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@139778.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@139779.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@139780.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@139781.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@139782.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@139783.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@139784.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@139785.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@139786.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@139787.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@139788.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@139789.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@139790.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@139791.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@139792.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@139793.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@139794.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@139795.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@139796.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@139797.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@139798.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@139799.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@139800.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@139801.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@139802.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@139803.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@139804.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@139805.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@139806.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@139807.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@139808.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@139809.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@139810.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@139811.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@139812.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@139813.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@139814.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@139815.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@139816.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@139817.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@139818.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@139819.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@139820.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@139821.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@139822.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@139823.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@139824.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@139825.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@139826.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@139827.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@139828.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@139829.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@139830.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@139831.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@139832.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@139833.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@139834.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@139835.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@139836.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@139837.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@139838.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@139839.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@139840.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@139841.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@139842.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@139843.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@139844.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@139845.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@139846.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@139847.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@139848.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@139849.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@139850.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@139851.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@139852.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@139853.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@139854.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@139855.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@139856.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@139857.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@139858.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@139859.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@139860.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@139861.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@139862.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@139863.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@139864.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@139865.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@139866.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@139867.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@139868.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@139869.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@139870.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@139871.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@139872.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@139873.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@139874.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@139875.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@139876.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@139877.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@139878.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@139879.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@139880.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@139881.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@139882.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@139883.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@139884.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@139885.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@139886.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@139887.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@139888.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@139889.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@139890.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@139891.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@139892.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@139893.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@139894.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@139895.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@139896.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@139897.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@139898.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@139899.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@139900.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@139901.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@139902.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@139903.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@139904.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@139905.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@139906.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@139907.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@139908.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@139909.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@139910.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@139911.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@139912.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@139913.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@139914.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@139915.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@139916.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@139917.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@139918.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@139919.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@139920.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@139921.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@139922.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@139923.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@139924.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@139925.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@139926.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@139927.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@139928.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@139929.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@139930.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@139931.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@139932.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@139933.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@139934.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@139935.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@139936.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@139937.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@139938.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@139939.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@139940.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@139941.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@139942.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@139943.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@139944.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@139945.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@139946.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@139947.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@139948.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@139949.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@139950.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@139951.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@139952.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@139953.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@139954.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@139955.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@139956.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@139957.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@139958.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@139959.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@139960.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@139961.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@139962.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@139963.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@139964.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@139965.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@139966.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@139967.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@139968.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@139969.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@139970.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@139971.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@139972.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@139973.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@139974.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@139975.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@139976.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@139977.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@139978.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@139979.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@139980.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@139981.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@139982.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@139983.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@139984.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@139985.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@139986.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@139987.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@139988.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@139989.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@139990.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@139991.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@139992.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@139993.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@139994.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@139995.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@139996.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@139997.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@139998.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@139999.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@140000.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@140001.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@140002.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@140003.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@140004.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@140005.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@140006.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@140007.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@140008.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@140009.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@140010.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@140011.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@140012.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@140013.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@140014.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@140015.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@140016.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@140017.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@140018.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@140019.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@140020.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@140021.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@140022.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@140023.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@140024.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@140025.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@140026.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@140027.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@140028.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@140029.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@140030.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@140031.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@140032.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@140033.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@140034.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@140035.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@140036.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@140037.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@140038.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@140039.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@140040.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@140041.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@140042.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@140043.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@140044.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@140045.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@140046.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@140047.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@140048.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@140049.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@140050.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@140051.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@140052.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@140053.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@140054.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@140055.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@140056.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@140057.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@140058.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@140059.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@140060.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@140061.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@140062.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@140063.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@140064.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@140065.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@140066.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@140067.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@140068.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@140069.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@140070.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@140071.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@140072.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@140073.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@140074.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@140075.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@140076.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@140077.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@140078.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@140079.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@140080.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@140081.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@140082.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@140083.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@140084.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@140085.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@140086.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@140087.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@140088.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@140089.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@140090.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@140091.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@140092.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@140093.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@140094.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@140095.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@140096.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@140097.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@140098.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@140099.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@140100.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@140101.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@140102.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@140103.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@140104.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@140105.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@140106.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@140107.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@140108.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@140109.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@140110.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@140111.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@140112.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@140113.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@140114.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@140115.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@140116.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@140117.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@140118.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@140119.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@140120.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@140121.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@140122.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@140123.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@140124.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@140125.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@140126.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@140127.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@140128.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@140129.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@140130.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@140131.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@140132.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@140133.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@140134.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@140135.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@140136.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@140137.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@140138.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@140139.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@140140.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@140141.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@140142.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@140143.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@140144.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@140145.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@140146.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@140147.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@140148.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@140149.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@140150.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@140151.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@140152.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@140153.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@140154.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@140155.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@140156.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@140157.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@140158.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@140159.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@140160.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@140161.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@140162.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@140163.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@140164.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@140165.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@140166.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@140167.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@140168.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@140169.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@140170.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@140171.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@140172.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@140173.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@140174.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@140175.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@140176.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@140177.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@140178.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@140179.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@140180.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@140181.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@140182.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@140183.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@140184.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@140185.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@140186.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@140187.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@140188.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@140189.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@140190.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@140191.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@140192.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@140193.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@140194.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@140195.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@140196.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@140197.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@140198.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@140199.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@140200.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@140201.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@140202.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@140203.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@140204.4]
endmodule
module RetimeWrapper_930( // @[:@140228.2]
  input         clock, // @[:@140229.4]
  input         reset, // @[:@140230.4]
  input  [39:0] io_in, // @[:@140231.4]
  output [39:0] io_out // @[:@140231.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@140233.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@140233.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@140233.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@140233.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@140233.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@140233.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@140233.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@140246.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@140245.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@140244.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@140243.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@140242.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@140240.4]
endmodule
module FringeFF_503( // @[:@140248.2]
  input         clock, // @[:@140249.4]
  input         reset, // @[:@140250.4]
  input  [39:0] io_in, // @[:@140251.4]
  output [39:0] io_out, // @[:@140251.4]
  input         io_enable // @[:@140251.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@140254.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@140254.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@140254.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@140254.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@140259.4 package.scala 96:25:@140260.4]
  RetimeWrapper_930 RetimeWrapper ( // @[package.scala 93:22:@140254.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@140259.4 package.scala 96:25:@140260.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@140271.4]
  assign RetimeWrapper_clock = clock; // @[:@140255.4]
  assign RetimeWrapper_reset = reset; // @[:@140256.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@140257.4]
endmodule
module FringeCounter( // @[:@140273.2]
  input   clock, // @[:@140274.4]
  input   reset, // @[:@140275.4]
  input   io_enable, // @[:@140276.4]
  output  io_done // @[:@140276.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@140278.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@140278.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@140278.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@140278.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@140278.4]
  wire [40:0] count; // @[Cat.scala 30:58:@140285.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@140286.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@140287.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@140288.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@140290.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@140278.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@140285.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@140286.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@140287.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@140288.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@140290.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@140301.4]
  assign reg$_clock = clock; // @[:@140279.4]
  assign reg$_reset = reset; // @[:@140280.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@140292.6 FringeCounter.scala 37:15:@140295.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@140283.4]
endmodule
module FringeFF_504( // @[:@140335.2]
  input   clock, // @[:@140336.4]
  input   reset, // @[:@140337.4]
  input   io_in, // @[:@140338.4]
  input   io_reset, // @[:@140338.4]
  output  io_out, // @[:@140338.4]
  input   io_enable // @[:@140338.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@140341.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@140341.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@140341.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@140341.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@140341.4]
  wire  _T_18; // @[package.scala 96:25:@140346.4 package.scala 96:25:@140347.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@140352.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@140341.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@140346.4 package.scala 96:25:@140347.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@140352.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@140358.4]
  assign RetimeWrapper_clock = clock; // @[:@140342.4]
  assign RetimeWrapper_reset = reset; // @[:@140343.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@140345.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@140344.4]
endmodule
module Depulser( // @[:@140360.2]
  input   clock, // @[:@140361.4]
  input   reset, // @[:@140362.4]
  input   io_in, // @[:@140363.4]
  input   io_rst, // @[:@140363.4]
  output  io_out // @[:@140363.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@140365.4]
  wire  r_reset; // @[Depulser.scala 14:17:@140365.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@140365.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@140365.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@140365.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@140365.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@140365.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@140374.4]
  assign r_clock = clock; // @[:@140366.4]
  assign r_reset = reset; // @[:@140367.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@140369.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@140373.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@140372.4]
endmodule
module Fringe( // @[:@140376.2]
  input         clock, // @[:@140377.4]
  input         reset, // @[:@140378.4]
  input  [31:0] io_raddr, // @[:@140379.4]
  input         io_wen, // @[:@140379.4]
  input  [31:0] io_waddr, // @[:@140379.4]
  input  [63:0] io_wdata, // @[:@140379.4]
  output [63:0] io_rdata, // @[:@140379.4]
  output        io_enable, // @[:@140379.4]
  input         io_done, // @[:@140379.4]
  output        io_reset, // @[:@140379.4]
  output [63:0] io_argIns_0, // @[:@140379.4]
  output [63:0] io_argIns_1, // @[:@140379.4]
  input         io_argOuts_0_valid, // @[:@140379.4]
  input  [63:0] io_argOuts_0_bits, // @[:@140379.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@140379.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@140379.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@140379.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@140379.4]
  output        io_memStreams_stores_0_data_ready, // @[:@140379.4]
  input         io_memStreams_stores_0_data_valid, // @[:@140379.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@140379.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@140379.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@140379.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@140379.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@140379.4]
  input         io_dram_0_cmd_ready, // @[:@140379.4]
  output        io_dram_0_cmd_valid, // @[:@140379.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@140379.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@140379.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@140379.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@140379.4]
  input         io_dram_0_wdata_ready, // @[:@140379.4]
  output        io_dram_0_wdata_valid, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@140379.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@140379.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@140379.4]
  output        io_dram_0_rresp_ready, // @[:@140379.4]
  output        io_dram_0_wresp_ready, // @[:@140379.4]
  input         io_dram_0_wresp_valid, // @[:@140379.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@140379.4]
  input         io_dram_1_cmd_ready, // @[:@140379.4]
  output        io_dram_1_cmd_valid, // @[:@140379.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@140379.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@140379.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@140379.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@140379.4]
  input         io_dram_1_wdata_ready, // @[:@140379.4]
  output        io_dram_1_wdata_valid, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@140379.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@140379.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@140379.4]
  output        io_dram_1_rresp_ready, // @[:@140379.4]
  output        io_dram_1_wresp_ready, // @[:@140379.4]
  input         io_dram_1_wresp_valid, // @[:@140379.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@140379.4]
  input         io_dram_2_cmd_ready, // @[:@140379.4]
  output        io_dram_2_cmd_valid, // @[:@140379.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@140379.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@140379.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@140379.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@140379.4]
  input         io_dram_2_wdata_ready, // @[:@140379.4]
  output        io_dram_2_wdata_valid, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@140379.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@140379.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@140379.4]
  output        io_dram_2_rresp_ready, // @[:@140379.4]
  output        io_dram_2_wresp_ready, // @[:@140379.4]
  input         io_dram_2_wresp_valid, // @[:@140379.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@140379.4]
  input         io_dram_3_cmd_ready, // @[:@140379.4]
  output        io_dram_3_cmd_valid, // @[:@140379.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@140379.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@140379.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@140379.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@140379.4]
  input         io_dram_3_wdata_ready, // @[:@140379.4]
  output        io_dram_3_wdata_valid, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@140379.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@140379.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@140379.4]
  output        io_dram_3_rresp_ready, // @[:@140379.4]
  output        io_dram_3_wresp_ready, // @[:@140379.4]
  input         io_dram_3_wresp_valid, // @[:@140379.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@140379.4]
  input         io_heap_0_req_valid, // @[:@140379.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@140379.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@140379.4]
  output        io_heap_0_resp_valid, // @[:@140379.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@140379.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@140379.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@140385.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@140385.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@140385.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@140385.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@141378.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@141378.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@141378.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@142338.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@142338.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@142338.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@143298.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@143298.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@143298.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@143298.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@144258.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@144258.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@144258.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@144258.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@144258.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@144258.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@144267.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@144267.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@144267.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@144267.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@144267.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@144267.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@144267.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@144267.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@144267.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@146317.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@146317.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@146317.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@146317.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@146336.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@146336.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@146336.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@146336.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@146336.4]
  wire [63:0] _T_1020; // @[:@146294.4 :@146295.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@146296.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@146298.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@146300.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@146302.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@146304.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@146306.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@146308.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@146344.4]
  reg  _T_1047; // @[package.scala 152:20:@146347.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@146349.4]
  wire  _T_1049; // @[package.scala 153:8:@146350.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@146354.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@146355.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@146358.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@146359.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@146361.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@146362.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@146364.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@146367.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@146346.4 Fringe.scala 163:24:@146365.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@146346.4 Fringe.scala 162:28:@146363.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@146368.4]
  wire  alloc; // @[Fringe.scala 202:38:@147998.4]
  wire  dealloc; // @[Fringe.scala 203:40:@147999.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@148000.4]
  reg  _T_1572; // @[package.scala 152:20:@148001.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@148003.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@140385.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@141378.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@142338.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@143298.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@144258.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@144267.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@146317.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@146336.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@146294.4 :@146295.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@146296.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@146298.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@146300.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@146302.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@146304.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@146306.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@146308.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@146344.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@146349.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@146350.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@146354.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@146355.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@146358.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@146359.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@146361.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@146362.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@146364.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@146367.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@146346.4 Fringe.scala 163:24:@146365.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@146346.4 Fringe.scala 162:28:@146363.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@146368.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@147998.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@147999.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@148000.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@148003.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@146292.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@146312.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@146313.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@146334.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@146335.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@141304.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@141300.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@141295.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@141294.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@147496.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@147495.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@147494.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@147492.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@147491.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@147489.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@147473.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@147474.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@147475.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@147476.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@147477.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@147478.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@147479.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@147480.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@147481.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@147482.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@147483.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@147484.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@147485.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@147486.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@147487.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@147488.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@147409.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@147410.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@147411.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@147412.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@147413.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@147414.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@147415.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@147416.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@147417.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@147418.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@147419.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@147420.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@147421.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@147422.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@147423.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@147424.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@147425.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@147426.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@147427.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@147428.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@147429.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@147430.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@147431.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@147432.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@147433.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@147434.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@147435.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@147436.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@147437.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@147438.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@147439.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@147440.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@147441.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@147442.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@147443.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@147444.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@147445.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@147446.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@147447.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@147448.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@147449.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@147450.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@147451.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@147452.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@147453.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@147454.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@147455.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@147456.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@147457.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@147458.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@147459.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@147460.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@147461.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@147462.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@147463.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@147464.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@147465.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@147466.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@147467.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@147468.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@147469.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@147470.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@147471.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@147472.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@147408.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@147407.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@147388.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@147608.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@147607.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@147606.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@147604.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@147603.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@147601.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@147585.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@147586.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@147587.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@147588.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@147589.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@147590.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@147591.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@147592.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@147593.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@147594.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@147595.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@147596.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@147597.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@147598.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@147599.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@147600.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@147521.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@147522.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@147523.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@147524.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@147525.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@147526.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@147527.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@147528.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@147529.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@147530.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@147531.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@147532.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@147533.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@147534.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@147535.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@147536.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@147537.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@147538.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@147539.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@147540.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@147541.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@147542.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@147543.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@147544.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@147545.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@147546.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@147547.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@147548.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@147549.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@147550.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@147551.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@147552.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@147553.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@147554.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@147555.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@147556.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@147557.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@147558.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@147559.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@147560.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@147561.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@147562.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@147563.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@147564.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@147565.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@147566.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@147567.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@147568.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@147569.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@147570.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@147571.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@147572.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@147573.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@147574.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@147575.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@147576.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@147577.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@147578.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@147579.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@147580.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@147581.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@147582.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@147583.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@147584.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@147520.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@147519.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@147500.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@147720.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@147719.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@147718.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@147716.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@147715.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@147713.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@147697.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@147698.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@147699.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@147700.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@147701.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@147702.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@147703.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@147704.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@147705.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@147706.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@147707.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@147708.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@147709.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@147710.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@147711.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@147712.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@147633.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@147634.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@147635.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@147636.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@147637.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@147638.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@147639.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@147640.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@147641.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@147642.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@147643.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@147644.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@147645.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@147646.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@147647.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@147648.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@147649.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@147650.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@147651.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@147652.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@147653.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@147654.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@147655.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@147656.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@147657.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@147658.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@147659.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@147660.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@147661.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@147662.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@147663.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@147664.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@147665.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@147666.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@147667.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@147668.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@147669.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@147670.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@147671.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@147672.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@147673.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@147674.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@147675.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@147676.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@147677.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@147678.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@147679.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@147680.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@147681.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@147682.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@147683.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@147684.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@147685.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@147686.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@147687.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@147688.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@147689.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@147690.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@147691.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@147692.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@147693.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@147694.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@147695.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@147696.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@147632.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@147631.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@147612.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@147832.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@147831.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@147830.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@147828.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@147827.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@147825.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@147809.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@147810.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@147811.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@147812.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@147813.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@147814.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@147815.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@147816.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@147817.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@147818.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@147819.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@147820.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@147821.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@147822.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@147823.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@147824.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@147745.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@147746.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@147747.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@147748.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@147749.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@147750.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@147751.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@147752.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@147753.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@147754.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@147755.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@147756.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@147757.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@147758.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@147759.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@147760.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@147761.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@147762.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@147763.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@147764.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@147765.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@147766.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@147767.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@147768.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@147769.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@147770.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@147771.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@147772.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@147773.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@147774.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@147775.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@147776.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@147777.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@147778.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@147779.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@147780.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@147781.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@147782.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@147783.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@147784.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@147785.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@147786.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@147787.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@147788.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@147789.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@147790.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@147791.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@147792.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@147793.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@147794.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@147795.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@147796.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@147797.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@147798.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@147799.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@147800.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@147801.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@147802.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@147803.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@147804.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@147805.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@147806.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@147807.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@147808.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@147744.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@147743.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@147724.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@144263.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@144262.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@144261.4]
  assign dramArbs_0_clock = clock; // @[:@140386.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@140387.4 Fringe.scala 187:30:@147378.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147382.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@141303.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@141302.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@141301.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@141299.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@141298.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@141297.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@141296.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@147497.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@147490.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@147387.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@147386.4]
  assign dramArbs_1_clock = clock; // @[:@141379.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@141380.4 Fringe.scala 187:30:@147379.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147383.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@147609.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@147602.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@147499.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@147498.4]
  assign dramArbs_2_clock = clock; // @[:@142339.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@142340.4 Fringe.scala 187:30:@147380.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147384.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@147721.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@147714.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@147611.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@147610.4]
  assign dramArbs_3_clock = clock; // @[:@143299.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@143300.4 Fringe.scala 187:30:@147381.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@147385.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@147833.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@147826.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@147723.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@147722.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@144266.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@144265.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@144264.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@148005.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@148006.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@148007.4]
  assign regs_clock = clock; // @[:@144268.4]
  assign regs_reset = reset; // @[:@144269.4 Fringe.scala 139:14:@146316.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@146288.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@146290.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@146289.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@146291.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@146314.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@146366.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@146370.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@146373.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@146372.4]
  assign timeoutCtr_clock = clock; // @[:@146318.4]
  assign timeoutCtr_reset = reset; // @[:@146319.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@146333.4]
  assign depulser_clock = clock; // @[:@146337.4]
  assign depulser_reset = reset; // @[:@146338.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@146343.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@146345.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@148022.2]
  input         clock, // @[:@148023.4]
  input         reset, // @[:@148024.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@148025.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@148025.4]
  input         io_S_AXI_AWVALID, // @[:@148025.4]
  output        io_S_AXI_AWREADY, // @[:@148025.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@148025.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@148025.4]
  input         io_S_AXI_ARVALID, // @[:@148025.4]
  output        io_S_AXI_ARREADY, // @[:@148025.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@148025.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@148025.4]
  input         io_S_AXI_WVALID, // @[:@148025.4]
  output        io_S_AXI_WREADY, // @[:@148025.4]
  output [31:0] io_S_AXI_RDATA, // @[:@148025.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@148025.4]
  output        io_S_AXI_RVALID, // @[:@148025.4]
  input         io_S_AXI_RREADY, // @[:@148025.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@148025.4]
  output        io_S_AXI_BVALID, // @[:@148025.4]
  input         io_S_AXI_BREADY, // @[:@148025.4]
  output [31:0] io_raddr, // @[:@148025.4]
  output        io_wen, // @[:@148025.4]
  output [31:0] io_waddr, // @[:@148025.4]
  output [31:0] io_wdata, // @[:@148025.4]
  input  [31:0] io_rdata // @[:@148025.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@148027.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148051.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148047.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148043.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@148042.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@148041.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148040.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@148038.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148037.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@148059.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@148062.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@148060.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@148061.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@148063.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@148058.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@148055.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@148054.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@148053.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148052.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@148050.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@148049.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148048.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@148046.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@148045.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@148044.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148039.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@148036.4]
endmodule
module MAGToAXI4Bridge( // @[:@148065.2]
  output         io_in_cmd_ready, // @[:@148068.4]
  input          io_in_cmd_valid, // @[:@148068.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@148068.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@148068.4]
  input          io_in_cmd_bits_isWr, // @[:@148068.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@148068.4]
  output         io_in_wdata_ready, // @[:@148068.4]
  input          io_in_wdata_valid, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@148068.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@148068.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@148068.4]
  input          io_in_wdata_bits_wlast, // @[:@148068.4]
  input          io_in_rresp_ready, // @[:@148068.4]
  input          io_in_wresp_ready, // @[:@148068.4]
  output         io_in_wresp_valid, // @[:@148068.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@148068.4]
  output [31:0]  io_M_AXI_AWID, // @[:@148068.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@148068.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@148068.4]
  output         io_M_AXI_AWVALID, // @[:@148068.4]
  input          io_M_AXI_AWREADY, // @[:@148068.4]
  output [31:0]  io_M_AXI_ARID, // @[:@148068.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@148068.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@148068.4]
  output         io_M_AXI_ARVALID, // @[:@148068.4]
  input          io_M_AXI_ARREADY, // @[:@148068.4]
  output [511:0] io_M_AXI_WDATA, // @[:@148068.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@148068.4]
  output         io_M_AXI_WLAST, // @[:@148068.4]
  output         io_M_AXI_WVALID, // @[:@148068.4]
  input          io_M_AXI_WREADY, // @[:@148068.4]
  output         io_M_AXI_RREADY, // @[:@148068.4]
  input  [31:0]  io_M_AXI_BID, // @[:@148068.4]
  input          io_M_AXI_BVALID, // @[:@148068.4]
  output         io_M_AXI_BREADY // @[:@148068.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@148225.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@148226.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@148227.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@148235.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@148262.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@148267.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@148278.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@148287.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@148296.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@148305.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@148314.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@148323.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@148331.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@148225.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@148226.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@148227.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@148235.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@148262.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@148267.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@148278.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@148287.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@148296.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@148305.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@148314.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@148323.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@148331.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@148239.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@148336.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@148389.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@148391.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@148240.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@148241.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@148245.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@148253.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@148223.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@148224.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@148228.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@148237.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@148269.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@148333.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@148334.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@148335.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@148386.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@148387.4]
endmodule
module FringeZynq( // @[:@149377.2]
  input          clock, // @[:@149378.4]
  input          reset, // @[:@149379.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@149380.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@149380.4]
  input          io_S_AXI_AWVALID, // @[:@149380.4]
  output         io_S_AXI_AWREADY, // @[:@149380.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@149380.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@149380.4]
  input          io_S_AXI_ARVALID, // @[:@149380.4]
  output         io_S_AXI_ARREADY, // @[:@149380.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@149380.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@149380.4]
  input          io_S_AXI_WVALID, // @[:@149380.4]
  output         io_S_AXI_WREADY, // @[:@149380.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@149380.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@149380.4]
  output         io_S_AXI_RVALID, // @[:@149380.4]
  input          io_S_AXI_RREADY, // @[:@149380.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@149380.4]
  output         io_S_AXI_BVALID, // @[:@149380.4]
  input          io_S_AXI_BREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@149380.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@149380.4]
  output         io_M_AXI_0_AWVALID, // @[:@149380.4]
  input          io_M_AXI_0_AWREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@149380.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@149380.4]
  output         io_M_AXI_0_ARVALID, // @[:@149380.4]
  input          io_M_AXI_0_ARREADY, // @[:@149380.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@149380.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@149380.4]
  output         io_M_AXI_0_WLAST, // @[:@149380.4]
  output         io_M_AXI_0_WVALID, // @[:@149380.4]
  input          io_M_AXI_0_WREADY, // @[:@149380.4]
  output         io_M_AXI_0_RREADY, // @[:@149380.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@149380.4]
  input          io_M_AXI_0_BVALID, // @[:@149380.4]
  output         io_M_AXI_0_BREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@149380.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@149380.4]
  output         io_M_AXI_1_AWVALID, // @[:@149380.4]
  input          io_M_AXI_1_AWREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@149380.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@149380.4]
  output         io_M_AXI_1_ARVALID, // @[:@149380.4]
  input          io_M_AXI_1_ARREADY, // @[:@149380.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@149380.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@149380.4]
  output         io_M_AXI_1_WLAST, // @[:@149380.4]
  output         io_M_AXI_1_WVALID, // @[:@149380.4]
  input          io_M_AXI_1_WREADY, // @[:@149380.4]
  output         io_M_AXI_1_RREADY, // @[:@149380.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@149380.4]
  input          io_M_AXI_1_BVALID, // @[:@149380.4]
  output         io_M_AXI_1_BREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@149380.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@149380.4]
  output         io_M_AXI_2_AWVALID, // @[:@149380.4]
  input          io_M_AXI_2_AWREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@149380.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@149380.4]
  output         io_M_AXI_2_ARVALID, // @[:@149380.4]
  input          io_M_AXI_2_ARREADY, // @[:@149380.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@149380.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@149380.4]
  output         io_M_AXI_2_WLAST, // @[:@149380.4]
  output         io_M_AXI_2_WVALID, // @[:@149380.4]
  input          io_M_AXI_2_WREADY, // @[:@149380.4]
  output         io_M_AXI_2_RREADY, // @[:@149380.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@149380.4]
  input          io_M_AXI_2_BVALID, // @[:@149380.4]
  output         io_M_AXI_2_BREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@149380.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@149380.4]
  output         io_M_AXI_3_AWVALID, // @[:@149380.4]
  input          io_M_AXI_3_AWREADY, // @[:@149380.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@149380.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@149380.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@149380.4]
  output         io_M_AXI_3_ARVALID, // @[:@149380.4]
  input          io_M_AXI_3_ARREADY, // @[:@149380.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@149380.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@149380.4]
  output         io_M_AXI_3_WLAST, // @[:@149380.4]
  output         io_M_AXI_3_WVALID, // @[:@149380.4]
  input          io_M_AXI_3_WREADY, // @[:@149380.4]
  output         io_M_AXI_3_RREADY, // @[:@149380.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@149380.4]
  input          io_M_AXI_3_BVALID, // @[:@149380.4]
  output         io_M_AXI_3_BREADY, // @[:@149380.4]
  output         io_enable, // @[:@149380.4]
  input          io_done, // @[:@149380.4]
  output         io_reset, // @[:@149380.4]
  output [63:0]  io_argIns_0, // @[:@149380.4]
  output [63:0]  io_argIns_1, // @[:@149380.4]
  input          io_argOuts_0_valid, // @[:@149380.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@149380.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@149380.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@149380.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@149380.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@149380.4]
  output         io_memStreams_stores_0_data_ready, // @[:@149380.4]
  input          io_memStreams_stores_0_data_valid, // @[:@149380.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@149380.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@149380.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@149380.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@149380.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@149380.4]
  input          io_heap_0_req_valid, // @[:@149380.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@149380.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@149380.4]
  output         io_heap_0_resp_valid, // @[:@149380.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@149380.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@149380.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@149851.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@149851.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@149851.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@150757.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@150757.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@150757.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@150757.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@150757.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@150757.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@150757.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@150757.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@150907.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@150907.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@150907.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@150907.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@150907.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@150907.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@150907.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151063.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151063.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151063.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151063.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151063.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151063.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151063.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151219.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151219.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151219.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151219.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151219.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151219.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151219.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@151375.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@151375.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@151375.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@151375.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@151375.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@151375.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@151375.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@151375.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@149851.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@150757.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@150907.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@151063.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@151219.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@151375.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@150775.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@150771.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@150767.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@150766.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@150765.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@150764.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@150762.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@150761.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151062.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151060.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151059.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151052.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151050.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151048.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151047.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151040.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151038.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151037.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151036.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151035.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151027.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151022.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151218.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151216.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151215.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151208.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151206.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151204.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151203.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151196.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151194.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151193.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151192.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151191.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151183.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151178.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151374.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151372.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151371.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151364.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151362.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151360.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151359.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151352.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151350.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151349.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151348.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151347.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151339.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151334.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@151530.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@151528.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@151527.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@151520.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@151518.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@151516.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@151515.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@151508.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@151506.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@151505.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@151504.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@151503.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@151495.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@151490.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@150785.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@150789.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@150790.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@150791.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@150878.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@150874.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@150869.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@150868.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@150903.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@150902.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@150901.4]
  assign fringeCommon_clock = clock; // @[:@149852.4]
  assign fringeCommon_reset = reset; // @[:@149853.4 FringeZynq.scala 117:22:@150788.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@150779.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@150780.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@150781.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@150782.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@150786.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@150793.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@150792.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@150877.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@150876.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@150875.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@150873.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@150872.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@150871.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@150870.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151021.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151014.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@150911.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@150910.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151177.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151170.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151067.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151066.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151333.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151326.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151223.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151222.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@151489.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@151482.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@151379.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@151378.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@150906.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@150905.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@150904.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@150758.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@150759.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@150778.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@150777.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@150776.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@150774.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@150773.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@150772.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@150770.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@150769.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@150768.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@150763.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@150760.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@150783.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@151020.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151019.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@151018.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151016.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151015.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@151013.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@150997.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@150998.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@150999.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151000.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151001.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151002.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151003.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151004.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151005.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151006.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151007.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151008.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151009.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151010.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151011.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151012.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@150933.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@150934.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@150935.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@150936.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@150937.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@150938.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@150939.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@150940.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@150941.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@150942.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@150943.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@150944.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@150945.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@150946.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@150947.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@150948.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@150949.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@150950.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@150951.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@150952.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@150953.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@150954.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@150955.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@150956.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@150957.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@150958.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@150959.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@150960.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@150961.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@150962.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@150963.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@150964.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@150965.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@150966.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@150967.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@150968.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@150969.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@150970.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@150971.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@150972.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@150973.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@150974.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@150975.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@150976.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@150977.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@150978.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@150979.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@150980.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@150981.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@150982.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@150983.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@150984.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@150985.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@150986.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@150987.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@150988.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@150989.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@150990.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@150991.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@150992.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@150993.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@150994.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@150995.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@150996.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@150932.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@150931.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@150912.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@151051.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@151039.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@151034.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@151026.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@151023.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@151176.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151175.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@151174.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151172.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151171.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@151169.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@151153.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@151154.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@151155.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151156.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151157.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151158.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151159.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151160.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151161.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151162.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151163.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151164.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151165.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151166.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151167.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151168.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151089.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151090.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151091.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151092.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151093.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151094.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151095.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151096.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151097.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151098.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151099.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151100.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151101.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151102.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151103.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151104.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151105.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151106.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151107.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151108.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151109.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151110.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151111.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151112.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151113.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151114.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151115.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151116.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151117.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@151118.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@151119.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@151120.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@151121.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@151122.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@151123.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@151124.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@151125.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@151126.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@151127.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@151128.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@151129.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@151130.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@151131.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@151132.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@151133.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@151134.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@151135.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@151136.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@151137.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@151138.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@151139.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@151140.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@151141.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@151142.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@151143.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@151144.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@151145.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@151146.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@151147.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@151148.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@151149.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@151150.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@151151.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@151152.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151088.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@151087.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@151068.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@151207.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@151195.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@151190.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@151182.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@151179.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@151332.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151331.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@151330.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151328.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151327.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@151325.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@151309.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@151310.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@151311.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151312.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151313.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151314.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151315.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151316.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151317.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151318.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151319.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151320.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151321.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151322.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151323.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151324.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151245.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151246.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151247.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151248.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151249.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151250.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151251.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151252.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151253.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151254.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151255.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151256.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151257.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151258.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151259.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151260.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151261.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151262.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151263.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151264.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151265.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151266.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151267.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151268.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151269.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151270.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151271.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151272.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151273.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@151274.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@151275.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@151276.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@151277.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@151278.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@151279.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@151280.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@151281.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@151282.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@151283.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@151284.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@151285.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@151286.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@151287.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@151288.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@151289.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@151290.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@151291.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@151292.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@151293.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@151294.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@151295.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@151296.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@151297.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@151298.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@151299.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@151300.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@151301.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@151302.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@151303.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@151304.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@151305.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@151306.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@151307.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@151308.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151244.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@151243.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@151224.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@151363.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@151351.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@151346.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@151338.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@151335.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@151488.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@151487.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@151486.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@151484.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@151483.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@151481.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@151465.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@151466.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@151467.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@151468.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@151469.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@151470.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@151471.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@151472.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@151473.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@151474.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@151475.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@151476.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@151477.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@151478.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@151479.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@151480.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@151401.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@151402.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@151403.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@151404.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@151405.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@151406.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@151407.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@151408.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@151409.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@151410.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@151411.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@151412.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@151413.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@151414.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@151415.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@151416.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@151417.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@151418.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@151419.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@151420.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@151421.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@151422.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@151423.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@151424.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@151425.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@151426.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@151427.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@151428.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@151429.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@151430.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@151431.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@151432.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@151433.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@151434.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@151435.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@151436.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@151437.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@151438.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@151439.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@151440.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@151441.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@151442.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@151443.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@151444.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@151445.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@151446.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@151447.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@151448.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@151449.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@151450.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@151451.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@151452.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@151453.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@151454.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@151455.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@151456.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@151457.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@151458.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@151459.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@151460.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@151461.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@151462.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@151463.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@151464.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@151400.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@151399.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@151380.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@151519.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@151507.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@151502.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@151494.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@151491.4]
endmodule
module SpatialIP( // @[:@151532.2]
  input          clock, // @[:@151533.4]
  input          reset, // @[:@151534.4]
  input          io_raddr, // @[:@151535.4]
  input          io_wen, // @[:@151535.4]
  input          io_waddr, // @[:@151535.4]
  input          io_wdata, // @[:@151535.4]
  output         io_rdata, // @[:@151535.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@151535.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@151535.4]
  input          io_S_AXI_AWVALID, // @[:@151535.4]
  output         io_S_AXI_AWREADY, // @[:@151535.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@151535.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@151535.4]
  input          io_S_AXI_ARVALID, // @[:@151535.4]
  output         io_S_AXI_ARREADY, // @[:@151535.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@151535.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@151535.4]
  input          io_S_AXI_WVALID, // @[:@151535.4]
  output         io_S_AXI_WREADY, // @[:@151535.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@151535.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@151535.4]
  output         io_S_AXI_RVALID, // @[:@151535.4]
  input          io_S_AXI_RREADY, // @[:@151535.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@151535.4]
  output         io_S_AXI_BVALID, // @[:@151535.4]
  input          io_S_AXI_BREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@151535.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@151535.4]
  output         io_M_AXI_0_AWLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@151535.4]
  output         io_M_AXI_0_AWVALID, // @[:@151535.4]
  input          io_M_AXI_0_AWREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@151535.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@151535.4]
  output         io_M_AXI_0_ARLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@151535.4]
  output         io_M_AXI_0_ARVALID, // @[:@151535.4]
  input          io_M_AXI_0_ARREADY, // @[:@151535.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@151535.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@151535.4]
  output         io_M_AXI_0_WLAST, // @[:@151535.4]
  output         io_M_AXI_0_WVALID, // @[:@151535.4]
  input          io_M_AXI_0_WREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@151535.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@151535.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@151535.4]
  input          io_M_AXI_0_RLAST, // @[:@151535.4]
  input          io_M_AXI_0_RVALID, // @[:@151535.4]
  output         io_M_AXI_0_RREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@151535.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@151535.4]
  input          io_M_AXI_0_BVALID, // @[:@151535.4]
  output         io_M_AXI_0_BREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@151535.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@151535.4]
  output         io_M_AXI_1_AWLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@151535.4]
  output         io_M_AXI_1_AWVALID, // @[:@151535.4]
  input          io_M_AXI_1_AWREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@151535.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@151535.4]
  output         io_M_AXI_1_ARLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@151535.4]
  output         io_M_AXI_1_ARVALID, // @[:@151535.4]
  input          io_M_AXI_1_ARREADY, // @[:@151535.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@151535.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@151535.4]
  output         io_M_AXI_1_WLAST, // @[:@151535.4]
  output         io_M_AXI_1_WVALID, // @[:@151535.4]
  input          io_M_AXI_1_WREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@151535.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@151535.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@151535.4]
  input          io_M_AXI_1_RLAST, // @[:@151535.4]
  input          io_M_AXI_1_RVALID, // @[:@151535.4]
  output         io_M_AXI_1_RREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@151535.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@151535.4]
  input          io_M_AXI_1_BVALID, // @[:@151535.4]
  output         io_M_AXI_1_BREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@151535.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@151535.4]
  output         io_M_AXI_2_AWLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@151535.4]
  output         io_M_AXI_2_AWVALID, // @[:@151535.4]
  input          io_M_AXI_2_AWREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@151535.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@151535.4]
  output         io_M_AXI_2_ARLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@151535.4]
  output         io_M_AXI_2_ARVALID, // @[:@151535.4]
  input          io_M_AXI_2_ARREADY, // @[:@151535.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@151535.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@151535.4]
  output         io_M_AXI_2_WLAST, // @[:@151535.4]
  output         io_M_AXI_2_WVALID, // @[:@151535.4]
  input          io_M_AXI_2_WREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@151535.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@151535.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@151535.4]
  input          io_M_AXI_2_RLAST, // @[:@151535.4]
  input          io_M_AXI_2_RVALID, // @[:@151535.4]
  output         io_M_AXI_2_RREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@151535.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@151535.4]
  input          io_M_AXI_2_BVALID, // @[:@151535.4]
  output         io_M_AXI_2_BREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@151535.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@151535.4]
  output         io_M_AXI_3_AWLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@151535.4]
  output         io_M_AXI_3_AWVALID, // @[:@151535.4]
  input          io_M_AXI_3_AWREADY, // @[:@151535.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@151535.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@151535.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@151535.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@151535.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@151535.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@151535.4]
  output         io_M_AXI_3_ARLOCK, // @[:@151535.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@151535.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@151535.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@151535.4]
  output         io_M_AXI_3_ARVALID, // @[:@151535.4]
  input          io_M_AXI_3_ARREADY, // @[:@151535.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@151535.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@151535.4]
  output         io_M_AXI_3_WLAST, // @[:@151535.4]
  output         io_M_AXI_3_WVALID, // @[:@151535.4]
  input          io_M_AXI_3_WREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@151535.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@151535.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@151535.4]
  input          io_M_AXI_3_RLAST, // @[:@151535.4]
  input          io_M_AXI_3_RVALID, // @[:@151535.4]
  output         io_M_AXI_3_RREADY, // @[:@151535.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@151535.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@151535.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@151535.4]
  input          io_M_AXI_3_BVALID, // @[:@151535.4]
  output         io_M_AXI_3_BREADY, // @[:@151535.4]
  input          io_TOP_AXI_AWID, // @[:@151535.4]
  input          io_TOP_AXI_AWUSER, // @[:@151535.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@151535.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@151535.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@151535.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@151535.4]
  input          io_TOP_AXI_AWLOCK, // @[:@151535.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@151535.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@151535.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@151535.4]
  input          io_TOP_AXI_AWVALID, // @[:@151535.4]
  input          io_TOP_AXI_AWREADY, // @[:@151535.4]
  input          io_TOP_AXI_ARID, // @[:@151535.4]
  input          io_TOP_AXI_ARUSER, // @[:@151535.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@151535.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@151535.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@151535.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@151535.4]
  input          io_TOP_AXI_ARLOCK, // @[:@151535.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@151535.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@151535.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@151535.4]
  input          io_TOP_AXI_ARVALID, // @[:@151535.4]
  input          io_TOP_AXI_ARREADY, // @[:@151535.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@151535.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@151535.4]
  input          io_TOP_AXI_WLAST, // @[:@151535.4]
  input          io_TOP_AXI_WVALID, // @[:@151535.4]
  input          io_TOP_AXI_WREADY, // @[:@151535.4]
  input          io_TOP_AXI_RID, // @[:@151535.4]
  input          io_TOP_AXI_RUSER, // @[:@151535.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@151535.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@151535.4]
  input          io_TOP_AXI_RLAST, // @[:@151535.4]
  input          io_TOP_AXI_RVALID, // @[:@151535.4]
  input          io_TOP_AXI_RREADY, // @[:@151535.4]
  input          io_TOP_AXI_BID, // @[:@151535.4]
  input          io_TOP_AXI_BUSER, // @[:@151535.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@151535.4]
  input          io_TOP_AXI_BVALID, // @[:@151535.4]
  input          io_TOP_AXI_BREADY, // @[:@151535.4]
  input          io_DWIDTH_AXI_AWID, // @[:@151535.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@151535.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@151535.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@151535.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@151535.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@151535.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@151535.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@151535.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@151535.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@151535.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@151535.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@151535.4]
  input          io_DWIDTH_AXI_ARID, // @[:@151535.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@151535.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@151535.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@151535.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@151535.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@151535.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@151535.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@151535.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@151535.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@151535.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@151535.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@151535.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@151535.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@151535.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@151535.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@151535.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@151535.4]
  input          io_DWIDTH_AXI_RID, // @[:@151535.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@151535.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@151535.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@151535.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@151535.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@151535.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@151535.4]
  input          io_DWIDTH_AXI_BID, // @[:@151535.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@151535.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@151535.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@151535.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@151535.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@151535.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@151535.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@151535.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@151535.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@151535.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@151535.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@151535.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@151535.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@151535.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@151535.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@151535.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@151535.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@151535.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@151535.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@151535.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@151535.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@151535.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@151535.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@151535.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@151535.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@151535.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@151535.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@151535.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@151535.4]
  input          io_PROTOCOL_AXI_RID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@151535.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@151535.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@151535.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@151535.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@151535.4]
  input          io_PROTOCOL_AXI_BID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@151535.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@151535.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@151535.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@151535.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@151535.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@151535.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@151535.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@151535.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@151535.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@151535.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@151535.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@151535.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@151535.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@151535.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@151535.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@151535.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@151535.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@151535.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@151535.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@151535.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@151535.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@151535.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@151535.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@151535.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@151537.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@151537.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@151537.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@151537.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@151537.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@151537.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@151537.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@151537.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@151537.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@151537.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@151679.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@151679.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@151679.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@151679.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@151679.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@151679.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@151679.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@151537.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@151679.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@151697.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@151693.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@151689.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@151688.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@151687.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@151686.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@151684.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@151683.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@151741.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@151740.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@151739.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@151738.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@151737.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@151736.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@151735.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@151734.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@151733.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@151732.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@151731.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@151729.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@151728.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@151727.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@151726.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@151725.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@151724.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@151723.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@151722.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@151721.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@151720.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@151719.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@151717.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@151716.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@151715.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@151714.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@151706.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@151701.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@151782.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@151781.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@151780.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@151779.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@151778.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@151777.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@151776.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@151775.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@151774.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@151773.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@151772.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@151770.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@151769.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@151768.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@151767.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@151766.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@151765.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@151764.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@151763.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@151762.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@151761.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@151760.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@151758.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@151757.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@151756.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@151755.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@151747.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@151742.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@151823.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@151822.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@151821.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@151820.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@151819.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@151818.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@151817.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@151816.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@151815.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@151814.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@151813.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@151811.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@151810.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@151809.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@151808.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@151807.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@151806.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@151805.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@151804.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@151803.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@151802.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@151801.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@151799.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@151798.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@151797.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@151796.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@151788.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@151783.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@151864.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@151863.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@151862.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@151861.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@151860.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@151859.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@151858.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@151857.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@151856.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@151855.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@151854.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@151852.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@151851.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@151850.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@151849.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@151848.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@151847.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@151846.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@151845.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@151844.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@151843.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@151842.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@151840.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@151839.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@151838.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@151837.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@151829.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@151824.4]
  assign accel_clock = clock; // @[:@151538.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@151539.4 Zynq.scala 54:17:@152153.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@152148.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@152141.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@152136.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@152120.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@152121.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@152122.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@152123.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@152124.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@152125.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@152126.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@152127.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@152128.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@152129.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@152130.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@152131.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@152132.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@152133.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@152134.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@152135.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@152119.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@152115.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@152110.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@152109.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@152108.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@152089.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@152073.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@152074.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@152075.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@152076.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@152077.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@152078.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@152079.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@152080.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@152081.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@152082.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@152083.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@152084.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@152085.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@152086.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@152087.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@152088.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@152072.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@152037.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@152036.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@152144.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@152143.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@152142.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@152030.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@152031.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@152034.4]
  assign FringeZynq_clock = clock; // @[:@151680.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@151681.4 Zynq.scala 53:18:@152152.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@151700.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@151699.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@151698.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@151696.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@151695.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@151694.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@151692.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@151691.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@151690.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@151685.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@151682.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@151730.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@151718.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@151713.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@151705.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@151702.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@151771.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@151759.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@151754.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@151746.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@151743.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@151812.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@151800.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@151795.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@151787.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@151784.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@151853.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@151841.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@151836.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@151828.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@151825.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@152149.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@152033.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@152032.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@152118.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@152117.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@152116.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@152114.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@152113.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@152112.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@152111.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@152147.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@152146.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@152145.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




