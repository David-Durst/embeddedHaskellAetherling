// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  output [31:0] O_0,
  output [31:0] O_1
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x253_TREADY(dontcare), // @[:@1298.4]
    .io_in_x253_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x253_TID(8'h0),
    .io_in_x253_TDEST(8'h0),
    .io_in_x254_TVALID(valid_down), // @[:@1298.4]
    .io_in_x254_TDATA({O_0,O_1}), // @[:@1298.4]
    .io_in_x254_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x261_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule


// End boilerplate
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh22); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh22); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x255_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x522_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x447_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x256_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x257_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x261_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x279_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x496_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x267_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x279_inr_Foreach_kernelx279_inr_Foreach_concrete1( // @[:@5106.2]
  input         clock, // @[:@5107.4]
  input         reset, // @[:@5108.4]
  output        io_in_x257_fifoinpacked_0_wPort_0_en_0, // @[:@5109.4]
  input         io_in_x257_fifoinpacked_0_full, // @[:@5109.4]
  output        io_in_x257_fifoinpacked_0_active_0_in, // @[:@5109.4]
  input         io_in_x257_fifoinpacked_0_active_0_out, // @[:@5109.4]
  input         io_sigsIn_backpressure, // @[:@5109.4]
  input         io_sigsIn_datapathEn, // @[:@5109.4]
  input         io_sigsIn_break, // @[:@5109.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5109.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5109.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5109.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5109.4]
  input         io_rr // @[:@5109.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@5143.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@5143.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@5155.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@5155.4]
  wire  x496_sub_1_clock; // @[Math.scala 191:24:@5182.4]
  wire  x496_sub_1_reset; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x496_sub_1_io_a; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x496_sub_1_io_b; // @[Math.scala 191:24:@5182.4]
  wire  x496_sub_1_io_flow; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x496_sub_1_io_result; // @[Math.scala 191:24:@5182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5192.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5192.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5192.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5192.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5192.4]
  wire  x267_sum_1_clock; // @[Math.scala 150:24:@5201.4]
  wire  x267_sum_1_reset; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x267_sum_1_io_a; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x267_sum_1_io_b; // @[Math.scala 150:24:@5201.4]
  wire  x267_sum_1_io_flow; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x267_sum_1_io_result; // @[Math.scala 150:24:@5201.4]
  wire  x268_sum_1_clock; // @[Math.scala 150:24:@5213.4]
  wire  x268_sum_1_reset; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x268_sum_1_io_a; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x268_sum_1_io_b; // @[Math.scala 150:24:@5213.4]
  wire  x268_sum_1_io_flow; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x268_sum_1_io_result; // @[Math.scala 150:24:@5213.4]
  wire  x498_sum_1_clock; // @[Math.scala 150:24:@5228.4]
  wire  x498_sum_1_reset; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x498_sum_1_io_a; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x498_sum_1_io_b; // @[Math.scala 150:24:@5228.4]
  wire  x498_sum_1_io_flow; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x498_sum_1_io_result; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x271_1_io_b; // @[Math.scala 720:24:@5249.4]
  wire [31:0] x271_1_io_result; // @[Math.scala 720:24:@5249.4]
  wire  x272_sum_1_clock; // @[Math.scala 150:24:@5260.4]
  wire  x272_sum_1_reset; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x272_sum_1_io_a; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x272_sum_1_io_b; // @[Math.scala 150:24:@5260.4]
  wire  x272_sum_1_io_flow; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x272_sum_1_io_result; // @[Math.scala 150:24:@5260.4]
  wire  x501_sum_1_clock; // @[Math.scala 150:24:@5275.4]
  wire  x501_sum_1_reset; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x501_sum_1_io_a; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x501_sum_1_io_b; // @[Math.scala 150:24:@5275.4]
  wire  x501_sum_1_io_flow; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x501_sum_1_io_result; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x275_1_io_b; // @[Math.scala 720:24:@5296.4]
  wire [31:0] x275_1_io_result; // @[Math.scala 720:24:@5296.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5331.4]
  wire  _T_327; // @[sm_x279_inr_Foreach.scala 62:18:@5168.4]
  wire  _T_328; // @[sm_x279_inr_Foreach.scala 62:55:@5169.4]
  wire [31:0] b262_number; // @[Math.scala 723:22:@5148.4 Math.scala 724:14:@5149.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@5173.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@5173.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@5178.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@5178.4]
  wire [31:0] x268_sum_number; // @[Math.scala 154:22:@5219.4 Math.scala 155:14:@5220.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@5224.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@5224.4]
  wire [31:0] x498_sum_number; // @[Math.scala 154:22:@5234.4 Math.scala 155:14:@5235.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@5241.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@5243.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@5244.4]
  wire [31:0] x272_sum_number; // @[Math.scala 154:22:@5266.4 Math.scala 155:14:@5267.4]
  wire [33:0] _GEN_3; // @[Math.scala 461:32:@5271.4]
  wire [33:0] _T_381; // @[Math.scala 461:32:@5271.4]
  wire [31:0] x501_sum_number; // @[Math.scala 154:22:@5281.4 Math.scala 155:14:@5282.4]
  wire [31:0] _T_392; // @[Math.scala 406:49:@5288.4]
  wire [31:0] _T_394; // @[Math.scala 406:56:@5290.4]
  wire [31:0] _T_395; // @[Math.scala 406:56:@5291.4]
  wire  _T_415; // @[sm_x279_inr_Foreach.scala 103:131:@5328.4]
  wire  _T_419; // @[package.scala 96:25:@5336.4 package.scala 96:25:@5337.4]
  wire  _T_421; // @[implicits.scala 55:10:@5338.4]
  wire  _T_422; // @[sm_x279_inr_Foreach.scala 103:148:@5339.4]
  wire  _T_424; // @[sm_x279_inr_Foreach.scala 103:236:@5341.4]
  wire  _T_425; // @[sm_x279_inr_Foreach.scala 103:255:@5342.4]
  wire  x525_b264_D4; // @[package.scala 96:25:@5316.4 package.scala 96:25:@5317.4]
  wire  _T_428; // @[sm_x279_inr_Foreach.scala 103:291:@5344.4]
  wire  x526_b265_D4; // @[package.scala 96:25:@5325.4 package.scala 96:25:@5326.4]
  _ _ ( // @[Math.scala 720:24:@5143.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@5155.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x496_sub x496_sub_1 ( // @[Math.scala 191:24:@5182.4]
    .clock(x496_sub_1_clock),
    .reset(x496_sub_1_reset),
    .io_a(x496_sub_1_io_a),
    .io_b(x496_sub_1_io_b),
    .io_flow(x496_sub_1_io_flow),
    .io_result(x496_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5192.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x267_sum x267_sum_1 ( // @[Math.scala 150:24:@5201.4]
    .clock(x267_sum_1_clock),
    .reset(x267_sum_1_reset),
    .io_a(x267_sum_1_io_a),
    .io_b(x267_sum_1_io_b),
    .io_flow(x267_sum_1_io_flow),
    .io_result(x267_sum_1_io_result)
  );
  x267_sum x268_sum_1 ( // @[Math.scala 150:24:@5213.4]
    .clock(x268_sum_1_clock),
    .reset(x268_sum_1_reset),
    .io_a(x268_sum_1_io_a),
    .io_b(x268_sum_1_io_b),
    .io_flow(x268_sum_1_io_flow),
    .io_result(x268_sum_1_io_result)
  );
  x267_sum x498_sum_1 ( // @[Math.scala 150:24:@5228.4]
    .clock(x498_sum_1_clock),
    .reset(x498_sum_1_reset),
    .io_a(x498_sum_1_io_a),
    .io_b(x498_sum_1_io_b),
    .io_flow(x498_sum_1_io_flow),
    .io_result(x498_sum_1_io_result)
  );
  _ x271_1 ( // @[Math.scala 720:24:@5249.4]
    .io_b(x271_1_io_b),
    .io_result(x271_1_io_result)
  );
  x267_sum x272_sum_1 ( // @[Math.scala 150:24:@5260.4]
    .clock(x272_sum_1_clock),
    .reset(x272_sum_1_reset),
    .io_a(x272_sum_1_io_a),
    .io_b(x272_sum_1_io_b),
    .io_flow(x272_sum_1_io_flow),
    .io_result(x272_sum_1_io_result)
  );
  x267_sum x501_sum_1 ( // @[Math.scala 150:24:@5275.4]
    .clock(x501_sum_1_clock),
    .reset(x501_sum_1_reset),
    .io_a(x501_sum_1_io_a),
    .io_b(x501_sum_1_io_b),
    .io_flow(x501_sum_1_io_flow),
    .io_result(x501_sum_1_io_result)
  );
  _ x275_1 ( // @[Math.scala 720:24:@5296.4]
    .io_b(x275_1_io_b),
    .io_result(x275_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@5311.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@5320.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@5331.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x257_fifoinpacked_0_full; // @[sm_x279_inr_Foreach.scala 62:18:@5168.4]
  assign _T_328 = ~ io_in_x257_fifoinpacked_0_active_0_out; // @[sm_x279_inr_Foreach.scala 62:55:@5169.4]
  assign b262_number = __io_result; // @[Math.scala 723:22:@5148.4 Math.scala 724:14:@5149.4]
  assign _GEN_0 = {{11'd0}, b262_number}; // @[Math.scala 461:32:@5173.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@5173.4]
  assign _GEN_1 = {{7'd0}, b262_number}; // @[Math.scala 461:32:@5178.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@5178.4]
  assign x268_sum_number = x268_sum_1_io_result; // @[Math.scala 154:22:@5219.4 Math.scala 155:14:@5220.4]
  assign _GEN_2 = {{2'd0}, x268_sum_number}; // @[Math.scala 461:32:@5224.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@5224.4]
  assign x498_sum_number = x498_sum_1_io_result; // @[Math.scala 154:22:@5234.4 Math.scala 155:14:@5235.4]
  assign _T_364 = $signed(x498_sum_number); // @[Math.scala 406:49:@5241.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@5243.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@5244.4]
  assign x272_sum_number = x272_sum_1_io_result; // @[Math.scala 154:22:@5266.4 Math.scala 155:14:@5267.4]
  assign _GEN_3 = {{2'd0}, x272_sum_number}; // @[Math.scala 461:32:@5271.4]
  assign _T_381 = _GEN_3 << 2; // @[Math.scala 461:32:@5271.4]
  assign x501_sum_number = x501_sum_1_io_result; // @[Math.scala 154:22:@5281.4 Math.scala 155:14:@5282.4]
  assign _T_392 = $signed(x501_sum_number); // @[Math.scala 406:49:@5288.4]
  assign _T_394 = $signed(_T_392) & $signed(32'shff); // @[Math.scala 406:56:@5290.4]
  assign _T_395 = $signed(_T_394); // @[Math.scala 406:56:@5291.4]
  assign _T_415 = ~ io_sigsIn_break; // @[sm_x279_inr_Foreach.scala 103:131:@5328.4]
  assign _T_419 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5336.4 package.scala 96:25:@5337.4]
  assign _T_421 = io_rr ? _T_419 : 1'h0; // @[implicits.scala 55:10:@5338.4]
  assign _T_422 = _T_415 & _T_421; // @[sm_x279_inr_Foreach.scala 103:148:@5339.4]
  assign _T_424 = _T_422 & _T_415; // @[sm_x279_inr_Foreach.scala 103:236:@5341.4]
  assign _T_425 = _T_424 & io_sigsIn_backpressure; // @[sm_x279_inr_Foreach.scala 103:255:@5342.4]
  assign x525_b264_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5316.4 package.scala 96:25:@5317.4]
  assign _T_428 = _T_425 & x525_b264_D4; // @[sm_x279_inr_Foreach.scala 103:291:@5344.4]
  assign x526_b265_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5325.4 package.scala 96:25:@5326.4]
  assign io_in_x257_fifoinpacked_0_wPort_0_en_0 = _T_428 & x526_b265_D4; // @[MemInterfaceType.scala 93:57:@5348.4]
  assign io_in_x257_fifoinpacked_0_active_0_in = x525_b264_D4 & x526_b265_D4; // @[MemInterfaceType.scala 147:18:@5351.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@5146.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@5158.4]
  assign x496_sub_1_clock = clock; // @[:@5183.4]
  assign x496_sub_1_reset = reset; // @[:@5184.4]
  assign x496_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@5185.4]
  assign x496_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@5186.4]
  assign x496_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5187.4]
  assign RetimeWrapper_clock = clock; // @[:@5193.4]
  assign RetimeWrapper_reset = reset; // @[:@5194.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5196.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5195.4]
  assign x267_sum_1_clock = clock; // @[:@5202.4]
  assign x267_sum_1_reset = reset; // @[:@5203.4]
  assign x267_sum_1_io_a = x496_sub_1_io_result; // @[Math.scala 151:17:@5204.4]
  assign x267_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5205.4]
  assign x267_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5206.4]
  assign x268_sum_1_clock = clock; // @[:@5214.4]
  assign x268_sum_1_reset = reset; // @[:@5215.4]
  assign x268_sum_1_io_a = x267_sum_1_io_result; // @[Math.scala 151:17:@5216.4]
  assign x268_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@5217.4]
  assign x268_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5218.4]
  assign x498_sum_1_clock = clock; // @[:@5229.4]
  assign x498_sum_1_reset = reset; // @[:@5230.4]
  assign x498_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@5231.4]
  assign x498_sum_1_io_b = x268_sum_1_io_result; // @[Math.scala 152:17:@5232.4]
  assign x498_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5233.4]
  assign x271_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@5252.4]
  assign x272_sum_1_clock = clock; // @[:@5261.4]
  assign x272_sum_1_reset = reset; // @[:@5262.4]
  assign x272_sum_1_io_a = x267_sum_1_io_result; // @[Math.scala 151:17:@5263.4]
  assign x272_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@5264.4]
  assign x272_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5265.4]
  assign x501_sum_1_clock = clock; // @[:@5276.4]
  assign x501_sum_1_reset = reset; // @[:@5277.4]
  assign x501_sum_1_io_a = _T_381[31:0]; // @[Math.scala 151:17:@5278.4]
  assign x501_sum_1_io_b = x272_sum_1_io_result; // @[Math.scala 152:17:@5279.4]
  assign x501_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5280.4]
  assign x275_1_io_b = $unsigned(_T_395); // @[Math.scala 721:17:@5299.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5312.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5313.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5315.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5314.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5321.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5322.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5324.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@5323.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5332.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5333.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5335.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5334.4]
endmodule
module RetimeWrapper_44( // @[:@6469.2]
  input   clock, // @[:@6470.4]
  input   reset, // @[:@6471.4]
  input   io_flow, // @[:@6472.4]
  input   io_in, // @[:@6472.4]
  output  io_out // @[:@6472.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(34)) sr ( // @[RetimeShiftRegister.scala 15:20:@6474.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6487.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6486.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6485.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6484.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6483.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6481.4]
endmodule
module RetimeWrapper_48( // @[:@6597.2]
  input   clock, // @[:@6598.4]
  input   reset, // @[:@6599.4]
  input   io_flow, // @[:@6600.4]
  input   io_in, // @[:@6600.4]
  output  io_out // @[:@6600.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(33)) sr ( // @[RetimeShiftRegister.scala 15:20:@6602.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6615.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6614.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6613.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6612.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6611.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6609.4]
endmodule
module x445_inr_Foreach_SAMPLER_BOX_sm( // @[:@6617.2]
  input   clock, // @[:@6618.4]
  input   reset, // @[:@6619.4]
  input   io_enable, // @[:@6620.4]
  output  io_done, // @[:@6620.4]
  output  io_doneLatch, // @[:@6620.4]
  input   io_ctrDone, // @[:@6620.4]
  output  io_datapathEn, // @[:@6620.4]
  output  io_ctrInc, // @[:@6620.4]
  output  io_ctrRst, // @[:@6620.4]
  input   io_parentAck, // @[:@6620.4]
  input   io_backpressure, // @[:@6620.4]
  input   io_break // @[:@6620.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6622.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6622.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6625.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6717.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6630.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6631.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6632.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6633.4]
  wire  _T_100; // @[package.scala 100:49:@6650.4]
  reg  _T_103; // @[package.scala 48:56:@6651.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6664.4 package.scala 96:25:@6665.4]
  wire  _T_110; // @[package.scala 100:49:@6666.4]
  reg  _T_113; // @[package.scala 48:56:@6667.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6669.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6674.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6675.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6678.4]
  wire  _T_124; // @[package.scala 96:25:@6686.4 package.scala 96:25:@6687.4]
  wire  _T_126; // @[package.scala 100:49:@6688.4]
  reg  _T_129; // @[package.scala 48:56:@6689.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6711.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6713.4]
  reg  _T_153; // @[package.scala 48:56:@6714.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6722.4 package.scala 96:25:@6723.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6724.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6725.4]
  SRFF active ( // @[Controllers.scala 261:22:@6622.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6625.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@6659.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@6681.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6693.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6701.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_4 ( // @[package.scala 93:22:@6717.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6630.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6631.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6632.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6633.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6650.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6664.4 package.scala 96:25:@6665.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6666.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6669.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6674.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6675.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6678.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6686.4 package.scala 96:25:@6687.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6688.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6713.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6722.4 package.scala 96:25:@6723.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6724.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6725.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6692.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6727.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6677.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6680.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6672.4]
  assign active_clock = clock; // @[:@6623.4]
  assign active_reset = reset; // @[:@6624.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6635.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6639.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6640.4]
  assign done_clock = clock; // @[:@6626.4]
  assign done_reset = reset; // @[:@6627.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6655.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6648.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6649.4]
  assign RetimeWrapper_clock = clock; // @[:@6660.4]
  assign RetimeWrapper_reset = reset; // @[:@6661.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6663.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6662.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6682.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6683.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6685.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6684.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6694.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6695.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6697.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6696.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6702.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6703.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6705.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6704.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6718.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6719.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6721.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6720.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_52( // @[:@6918.2]
  input         clock, // @[:@6919.4]
  input         reset, // @[:@6920.4]
  input         io_flow, // @[:@6921.4]
  input  [63:0] io_in, // @[:@6921.4]
  output [63:0] io_out // @[:@6921.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6923.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6936.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6935.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@6934.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6933.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6932.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6930.4]
endmodule
module SRAM_1( // @[:@6954.2]
  input         clock, // @[:@6955.4]
  input         reset, // @[:@6956.4]
  input  [8:0]  io_raddr, // @[:@6957.4]
  input         io_wen, // @[:@6957.4]
  input  [8:0]  io_waddr, // @[:@6957.4]
  input  [31:0] io_wdata, // @[:@6957.4]
  output [31:0] io_rdata, // @[:@6957.4]
  input         io_backpressure // @[:@6957.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6959.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6959.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6959.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6959.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6977.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6978.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6979.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6981.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(480), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6959.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6977.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6978.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6986.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6973.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6974.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6971.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6976.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6975.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6972.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6970.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6969.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_53( // @[:@7000.2]
  input        clock, // @[:@7001.4]
  input        reset, // @[:@7002.4]
  input        io_flow, // @[:@7003.4]
  input  [8:0] io_in, // @[:@7003.4]
  output [8:0] io_out // @[:@7003.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7005.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7018.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7017.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7016.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7015.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7014.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7012.4]
endmodule
module Mem1D_5( // @[:@7020.2]
  input         clock, // @[:@7021.4]
  input         reset, // @[:@7022.4]
  input  [8:0]  io_r_ofs_0, // @[:@7023.4]
  input         io_r_backpressure, // @[:@7023.4]
  input  [8:0]  io_w_ofs_0, // @[:@7023.4]
  input  [31:0] io_w_data_0, // @[:@7023.4]
  input         io_w_en_0, // @[:@7023.4]
  output [31:0] io_output // @[:@7023.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7030.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7030.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7030.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7030.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7030.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@7025.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@7027.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_53 RetimeWrapper ( // @[package.scala 93:22:@7030.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h1e0; // @[MemPrimitives.scala 702:32:@7025.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@7043.4]
  assign SRAM_clock = clock; // @[:@7028.4]
  assign SRAM_reset = reset; // @[:@7029.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@7037.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@7040.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@7038.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@7041.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@7042.4]
  assign RetimeWrapper_clock = clock; // @[:@7031.4]
  assign RetimeWrapper_reset = reset; // @[:@7032.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7034.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7033.4]
endmodule
module StickySelects_1( // @[:@8650.2]
  input   clock, // @[:@8651.4]
  input   reset, // @[:@8652.4]
  input   io_ins_0, // @[:@8653.4]
  input   io_ins_1, // @[:@8653.4]
  input   io_ins_2, // @[:@8653.4]
  input   io_ins_3, // @[:@8653.4]
  input   io_ins_4, // @[:@8653.4]
  input   io_ins_5, // @[:@8653.4]
  output  io_outs_0, // @[:@8653.4]
  output  io_outs_1, // @[:@8653.4]
  output  io_outs_2, // @[:@8653.4]
  output  io_outs_3, // @[:@8653.4]
  output  io_outs_4, // @[:@8653.4]
  output  io_outs_5 // @[:@8653.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@8655.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@8656.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@8657.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@8658.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@8659.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@8660.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@8661.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@8662.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@8663.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@8664.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@8665.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@8666.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@8668.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@8669.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@8670.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@8671.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@8672.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@8673.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@8675.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@8676.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@8677.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@8678.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@8679.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@8680.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@8683.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@8684.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@8685.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@8686.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@8687.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@8691.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@8692.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@8693.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@8694.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@8699.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@8700.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@8701.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@8661.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@8662.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@8663.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@8664.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@8665.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@8666.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@8668.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@8669.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@8670.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@8671.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@8672.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@8673.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@8675.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@8676.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@8677.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@8678.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@8679.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@8680.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@8683.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@8684.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@8685.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@8686.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@8687.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@8691.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@8692.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@8693.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@8694.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@8699.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@8700.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@8701.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@8703.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@8704.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@8705.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@8706.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@8707.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@8708.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x290_lb_0( // @[:@12682.2]
  input         clock, // @[:@12683.4]
  input         reset, // @[:@12684.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@12685.4]
  input         io_rPort_11_en_0, // @[:@12685.4]
  input         io_rPort_11_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_11_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@12685.4]
  input         io_rPort_10_en_0, // @[:@12685.4]
  input         io_rPort_10_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_10_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@12685.4]
  input         io_rPort_9_en_0, // @[:@12685.4]
  input         io_rPort_9_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_9_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@12685.4]
  input         io_rPort_8_en_0, // @[:@12685.4]
  input         io_rPort_8_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_8_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@12685.4]
  input         io_rPort_7_en_0, // @[:@12685.4]
  input         io_rPort_7_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_7_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@12685.4]
  input         io_rPort_6_en_0, // @[:@12685.4]
  input         io_rPort_6_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_6_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@12685.4]
  input         io_rPort_5_en_0, // @[:@12685.4]
  input         io_rPort_5_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_5_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@12685.4]
  input         io_rPort_4_en_0, // @[:@12685.4]
  input         io_rPort_4_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_4_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@12685.4]
  input         io_rPort_3_en_0, // @[:@12685.4]
  input         io_rPort_3_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_3_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@12685.4]
  input         io_rPort_2_en_0, // @[:@12685.4]
  input         io_rPort_2_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_2_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@12685.4]
  input         io_rPort_1_en_0, // @[:@12685.4]
  input         io_rPort_1_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_1_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@12685.4]
  input         io_rPort_0_en_0, // @[:@12685.4]
  input         io_rPort_0_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_0_output_0, // @[:@12685.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@12685.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@12685.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@12685.4]
  input  [31:0] io_wPort_1_data_0, // @[:@12685.4]
  input         io_wPort_1_en_0, // @[:@12685.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@12685.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12685.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@12685.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12685.4]
  input         io_wPort_0_en_0 // @[:@12685.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15353.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@13032.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@13033.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@13034.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@13035.4]
  wire [41:0] _T_450; // @[Cat.scala 30:58:@13037.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@13044.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@13045.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@13046.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@13047.4]
  wire [41:0] _T_461; // @[Cat.scala 30:58:@13049.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@13057.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@13058.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@13059.4]
  wire [41:0] _T_472; // @[Cat.scala 30:58:@13061.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@13069.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@13070.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@13071.4]
  wire [41:0] _T_483; // @[Cat.scala 30:58:@13073.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@13080.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@13082.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@13083.4]
  wire [41:0] _T_494; // @[Cat.scala 30:58:@13085.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@13092.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@13094.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@13095.4]
  wire [41:0] _T_505; // @[Cat.scala 30:58:@13097.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@13106.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@13107.4]
  wire [41:0] _T_516; // @[Cat.scala 30:58:@13109.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@13118.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@13119.4]
  wire [41:0] _T_527; // @[Cat.scala 30:58:@13121.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@13128.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@13130.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@13131.4]
  wire [41:0] _T_538; // @[Cat.scala 30:58:@13133.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@13140.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@13142.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@13143.4]
  wire [41:0] _T_549; // @[Cat.scala 30:58:@13145.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@13154.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@13155.4]
  wire [41:0] _T_560; // @[Cat.scala 30:58:@13157.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@13166.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@13167.4]
  wire [41:0] _T_571; // @[Cat.scala 30:58:@13169.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@13176.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@13178.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@13179.4]
  wire [41:0] _T_582; // @[Cat.scala 30:58:@13181.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@13188.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@13190.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@13191.4]
  wire [41:0] _T_593; // @[Cat.scala 30:58:@13193.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@13202.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@13203.4]
  wire [41:0] _T_604; // @[Cat.scala 30:58:@13205.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@13214.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@13215.4]
  wire [41:0] _T_615; // @[Cat.scala 30:58:@13217.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@13224.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@13225.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@13226.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@13228.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@13229.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@13230.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@13232.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13233.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13234.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@13236.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13237.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13238.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@13240.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13241.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13242.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@13244.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13245.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13246.4]
  wire  _T_655; // @[MemPrimitives.scala 126:35:@13257.4]
  wire  _T_656; // @[MemPrimitives.scala 126:35:@13258.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@13259.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@13260.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@13261.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@13262.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@13264.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@13266.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@13268.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@13270.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@13272.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@13274.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@13275.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@13276.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@13277.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@13278.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@13279.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13286.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@13287.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@13290.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@13291.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@13294.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@13295.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@13296.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@13298.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@13299.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@13300.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@13302.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@13303.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@13304.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@13306.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@13307.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@13308.4]
  wire  _T_717; // @[MemPrimitives.scala 126:35:@13319.4]
  wire  _T_718; // @[MemPrimitives.scala 126:35:@13320.4]
  wire  _T_719; // @[MemPrimitives.scala 126:35:@13321.4]
  wire  _T_720; // @[MemPrimitives.scala 126:35:@13322.4]
  wire  _T_721; // @[MemPrimitives.scala 126:35:@13323.4]
  wire  _T_722; // @[MemPrimitives.scala 126:35:@13324.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@13326.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@13328.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@13330.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@13332.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@13334.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@13336.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@13337.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@13338.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@13339.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@13340.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@13341.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@13349.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@13350.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@13353.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@13354.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@13357.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@13358.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@13361.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@13362.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@13365.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@13366.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@13369.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@13370.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13381.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13382.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13383.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13384.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13385.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13386.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@13388.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@13390.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@13392.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@13394.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@13396.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@13398.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@13399.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@13400.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@13401.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@13402.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@13403.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@13411.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@13412.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@13415.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@13416.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@13419.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@13420.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@13423.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@13424.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@13427.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@13428.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@13431.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@13432.4]
  wire  _T_841; // @[MemPrimitives.scala 126:35:@13443.4]
  wire  _T_842; // @[MemPrimitives.scala 126:35:@13444.4]
  wire  _T_843; // @[MemPrimitives.scala 126:35:@13445.4]
  wire  _T_844; // @[MemPrimitives.scala 126:35:@13446.4]
  wire  _T_845; // @[MemPrimitives.scala 126:35:@13447.4]
  wire  _T_846; // @[MemPrimitives.scala 126:35:@13448.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@13450.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@13452.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@13454.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@13456.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@13458.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@13460.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@13461.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@13462.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@13463.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@13464.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@13465.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@13472.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@13476.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@13480.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@13482.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@13484.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@13486.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@13488.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@13490.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@13492.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@13494.4]
  wire  _T_903; // @[MemPrimitives.scala 126:35:@13505.4]
  wire  _T_904; // @[MemPrimitives.scala 126:35:@13506.4]
  wire  _T_905; // @[MemPrimitives.scala 126:35:@13507.4]
  wire  _T_906; // @[MemPrimitives.scala 126:35:@13508.4]
  wire  _T_907; // @[MemPrimitives.scala 126:35:@13509.4]
  wire  _T_908; // @[MemPrimitives.scala 126:35:@13510.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@13512.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@13514.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@13516.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@13518.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@13520.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@13522.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@13523.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@13524.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@13525.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@13526.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@13527.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@13534.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@13536.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@13538.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@13540.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@13542.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@13544.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@13546.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@13548.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@13550.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@13552.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@13554.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@13556.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13567.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13568.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13569.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13570.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13571.4]
  wire  _T_970; // @[MemPrimitives.scala 126:35:@13572.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@13574.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@13576.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@13578.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@13580.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@13582.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@13584.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@13585.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@13586.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@13587.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@13588.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@13589.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@13598.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@13602.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@13606.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@13610.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@13614.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@13618.4]
  wire  _T_1027; // @[MemPrimitives.scala 126:35:@13629.4]
  wire  _T_1028; // @[MemPrimitives.scala 126:35:@13630.4]
  wire  _T_1029; // @[MemPrimitives.scala 126:35:@13631.4]
  wire  _T_1030; // @[MemPrimitives.scala 126:35:@13632.4]
  wire  _T_1031; // @[MemPrimitives.scala 126:35:@13633.4]
  wire  _T_1032; // @[MemPrimitives.scala 126:35:@13634.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@13636.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@13638.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@13640.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@13642.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@13644.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@13646.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@13647.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@13648.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@13649.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@13650.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@13651.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@13668.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@13672.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@13676.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@13680.4]
  wire  _T_1089; // @[MemPrimitives.scala 126:35:@13691.4]
  wire  _T_1090; // @[MemPrimitives.scala 126:35:@13692.4]
  wire  _T_1091; // @[MemPrimitives.scala 126:35:@13693.4]
  wire  _T_1092; // @[MemPrimitives.scala 126:35:@13694.4]
  wire  _T_1093; // @[MemPrimitives.scala 126:35:@13695.4]
  wire  _T_1094; // @[MemPrimitives.scala 126:35:@13696.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@13698.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@13700.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@13702.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@13704.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@13706.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@13708.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@13709.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@13710.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@13711.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@13712.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@13713.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@13720.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13722.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@13724.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13726.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@13728.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13730.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@13732.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13734.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@13736.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13738.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@13740.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@13742.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13753.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13754.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13755.4]
  wire  _T_1154; // @[MemPrimitives.scala 126:35:@13756.4]
  wire  _T_1155; // @[MemPrimitives.scala 126:35:@13757.4]
  wire  _T_1156; // @[MemPrimitives.scala 126:35:@13758.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@13760.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@13762.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@13764.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@13766.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@13768.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@13770.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@13771.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@13772.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@13773.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@13774.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@13775.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@13782.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@13784.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@13786.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13788.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@13790.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13792.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@13794.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13796.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@13798.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13800.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@13802.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13804.4]
  wire  _T_1213; // @[MemPrimitives.scala 126:35:@13815.4]
  wire  _T_1214; // @[MemPrimitives.scala 126:35:@13816.4]
  wire  _T_1215; // @[MemPrimitives.scala 126:35:@13817.4]
  wire  _T_1216; // @[MemPrimitives.scala 126:35:@13818.4]
  wire  _T_1217; // @[MemPrimitives.scala 126:35:@13819.4]
  wire  _T_1218; // @[MemPrimitives.scala 126:35:@13820.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@13822.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@13824.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@13826.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@13828.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@13830.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@13832.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@13833.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@13834.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@13835.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@13836.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@13837.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@13846.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@13850.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@13854.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@13858.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@13862.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@13866.4]
  wire  _T_1275; // @[MemPrimitives.scala 126:35:@13877.4]
  wire  _T_1276; // @[MemPrimitives.scala 126:35:@13878.4]
  wire  _T_1277; // @[MemPrimitives.scala 126:35:@13879.4]
  wire  _T_1278; // @[MemPrimitives.scala 126:35:@13880.4]
  wire  _T_1279; // @[MemPrimitives.scala 126:35:@13881.4]
  wire  _T_1280; // @[MemPrimitives.scala 126:35:@13882.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@13884.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@13886.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@13888.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@13890.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@13892.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@13894.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@13895.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@13896.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@13897.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@13898.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@13899.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@13908.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@13912.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@13916.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@13920.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@13924.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@13928.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13939.4]
  wire  _T_1338; // @[MemPrimitives.scala 126:35:@13940.4]
  wire  _T_1339; // @[MemPrimitives.scala 126:35:@13941.4]
  wire  _T_1340; // @[MemPrimitives.scala 126:35:@13942.4]
  wire  _T_1341; // @[MemPrimitives.scala 126:35:@13943.4]
  wire  _T_1342; // @[MemPrimitives.scala 126:35:@13944.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@13946.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@13948.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@13950.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@13952.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@13954.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@13956.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@13957.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@13958.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@13959.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@13960.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@13961.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@13968.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@13970.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@13972.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@13974.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@13976.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@13978.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@13980.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@13982.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@13984.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@13986.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@13988.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@13990.4]
  wire  _T_1399; // @[MemPrimitives.scala 126:35:@14001.4]
  wire  _T_1400; // @[MemPrimitives.scala 126:35:@14002.4]
  wire  _T_1401; // @[MemPrimitives.scala 126:35:@14003.4]
  wire  _T_1402; // @[MemPrimitives.scala 126:35:@14004.4]
  wire  _T_1403; // @[MemPrimitives.scala 126:35:@14005.4]
  wire  _T_1404; // @[MemPrimitives.scala 126:35:@14006.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@14008.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@14010.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@14012.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@14014.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@14016.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@14018.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@14019.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@14020.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@14021.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@14022.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@14023.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@14030.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@14032.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@14034.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@14036.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@14038.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@14040.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@14042.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@14044.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@14046.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@14048.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@14050.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@14052.4]
  wire  _T_1461; // @[MemPrimitives.scala 126:35:@14063.4]
  wire  _T_1462; // @[MemPrimitives.scala 126:35:@14064.4]
  wire  _T_1463; // @[MemPrimitives.scala 126:35:@14065.4]
  wire  _T_1464; // @[MemPrimitives.scala 126:35:@14066.4]
  wire  _T_1465; // @[MemPrimitives.scala 126:35:@14067.4]
  wire  _T_1466; // @[MemPrimitives.scala 126:35:@14068.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@14070.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@14072.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@14074.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@14076.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@14078.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@14080.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@14081.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@14082.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@14083.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@14084.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@14085.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@14094.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@14098.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@14102.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@14106.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@14110.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@14114.4]
  wire  _T_1523; // @[MemPrimitives.scala 126:35:@14125.4]
  wire  _T_1524; // @[MemPrimitives.scala 126:35:@14126.4]
  wire  _T_1525; // @[MemPrimitives.scala 126:35:@14127.4]
  wire  _T_1526; // @[MemPrimitives.scala 126:35:@14128.4]
  wire  _T_1527; // @[MemPrimitives.scala 126:35:@14129.4]
  wire  _T_1528; // @[MemPrimitives.scala 126:35:@14130.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@14132.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@14134.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@14136.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@14138.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@14140.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@14142.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@14143.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@14144.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@14145.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@14146.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@14147.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@14156.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@14160.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@14164.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@14168.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@14172.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@14176.4]
  wire  _T_1585; // @[MemPrimitives.scala 126:35:@14187.4]
  wire  _T_1586; // @[MemPrimitives.scala 126:35:@14188.4]
  wire  _T_1587; // @[MemPrimitives.scala 126:35:@14189.4]
  wire  _T_1588; // @[MemPrimitives.scala 126:35:@14190.4]
  wire  _T_1589; // @[MemPrimitives.scala 126:35:@14191.4]
  wire  _T_1590; // @[MemPrimitives.scala 126:35:@14192.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@14194.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@14196.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@14198.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@14200.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@14202.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@14204.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@14205.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@14206.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@14207.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@14208.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1671; // @[package.scala 96:25:@14294.4 package.scala 96:25:@14295.4]
  wire [31:0] _T_1675; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1668; // @[package.scala 96:25:@14286.4 package.scala 96:25:@14287.4]
  wire [31:0] _T_1676; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1665; // @[package.scala 96:25:@14278.4 package.scala 96:25:@14279.4]
  wire [31:0] _T_1677; // @[Mux.scala 31:69:@14306.4]
  wire  _T_1662; // @[package.scala 96:25:@14270.4 package.scala 96:25:@14271.4]
  wire [31:0] _T_1678; // @[Mux.scala 31:69:@14307.4]
  wire  _T_1659; // @[package.scala 96:25:@14262.4 package.scala 96:25:@14263.4]
  wire [31:0] _T_1679; // @[Mux.scala 31:69:@14308.4]
  wire  _T_1656; // @[package.scala 96:25:@14254.4 package.scala 96:25:@14255.4]
  wire [31:0] _T_1680; // @[Mux.scala 31:69:@14309.4]
  wire  _T_1653; // @[package.scala 96:25:@14246.4 package.scala 96:25:@14247.4]
  wire  _T_1742; // @[package.scala 96:25:@14390.4 package.scala 96:25:@14391.4]
  wire [31:0] _T_1746; // @[Mux.scala 31:69:@14400.4]
  wire  _T_1739; // @[package.scala 96:25:@14382.4 package.scala 96:25:@14383.4]
  wire [31:0] _T_1747; // @[Mux.scala 31:69:@14401.4]
  wire  _T_1736; // @[package.scala 96:25:@14374.4 package.scala 96:25:@14375.4]
  wire [31:0] _T_1748; // @[Mux.scala 31:69:@14402.4]
  wire  _T_1733; // @[package.scala 96:25:@14366.4 package.scala 96:25:@14367.4]
  wire [31:0] _T_1749; // @[Mux.scala 31:69:@14403.4]
  wire  _T_1730; // @[package.scala 96:25:@14358.4 package.scala 96:25:@14359.4]
  wire [31:0] _T_1750; // @[Mux.scala 31:69:@14404.4]
  wire  _T_1727; // @[package.scala 96:25:@14350.4 package.scala 96:25:@14351.4]
  wire [31:0] _T_1751; // @[Mux.scala 31:69:@14405.4]
  wire  _T_1724; // @[package.scala 96:25:@14342.4 package.scala 96:25:@14343.4]
  wire  _T_1813; // @[package.scala 96:25:@14486.4 package.scala 96:25:@14487.4]
  wire [31:0] _T_1817; // @[Mux.scala 31:69:@14496.4]
  wire  _T_1810; // @[package.scala 96:25:@14478.4 package.scala 96:25:@14479.4]
  wire [31:0] _T_1818; // @[Mux.scala 31:69:@14497.4]
  wire  _T_1807; // @[package.scala 96:25:@14470.4 package.scala 96:25:@14471.4]
  wire [31:0] _T_1819; // @[Mux.scala 31:69:@14498.4]
  wire  _T_1804; // @[package.scala 96:25:@14462.4 package.scala 96:25:@14463.4]
  wire [31:0] _T_1820; // @[Mux.scala 31:69:@14499.4]
  wire  _T_1801; // @[package.scala 96:25:@14454.4 package.scala 96:25:@14455.4]
  wire [31:0] _T_1821; // @[Mux.scala 31:69:@14500.4]
  wire  _T_1798; // @[package.scala 96:25:@14446.4 package.scala 96:25:@14447.4]
  wire [31:0] _T_1822; // @[Mux.scala 31:69:@14501.4]
  wire  _T_1795; // @[package.scala 96:25:@14438.4 package.scala 96:25:@14439.4]
  wire  _T_1884; // @[package.scala 96:25:@14582.4 package.scala 96:25:@14583.4]
  wire [31:0] _T_1888; // @[Mux.scala 31:69:@14592.4]
  wire  _T_1881; // @[package.scala 96:25:@14574.4 package.scala 96:25:@14575.4]
  wire [31:0] _T_1889; // @[Mux.scala 31:69:@14593.4]
  wire  _T_1878; // @[package.scala 96:25:@14566.4 package.scala 96:25:@14567.4]
  wire [31:0] _T_1890; // @[Mux.scala 31:69:@14594.4]
  wire  _T_1875; // @[package.scala 96:25:@14558.4 package.scala 96:25:@14559.4]
  wire [31:0] _T_1891; // @[Mux.scala 31:69:@14595.4]
  wire  _T_1872; // @[package.scala 96:25:@14550.4 package.scala 96:25:@14551.4]
  wire [31:0] _T_1892; // @[Mux.scala 31:69:@14596.4]
  wire  _T_1869; // @[package.scala 96:25:@14542.4 package.scala 96:25:@14543.4]
  wire [31:0] _T_1893; // @[Mux.scala 31:69:@14597.4]
  wire  _T_1866; // @[package.scala 96:25:@14534.4 package.scala 96:25:@14535.4]
  wire  _T_1955; // @[package.scala 96:25:@14678.4 package.scala 96:25:@14679.4]
  wire [31:0] _T_1959; // @[Mux.scala 31:69:@14688.4]
  wire  _T_1952; // @[package.scala 96:25:@14670.4 package.scala 96:25:@14671.4]
  wire [31:0] _T_1960; // @[Mux.scala 31:69:@14689.4]
  wire  _T_1949; // @[package.scala 96:25:@14662.4 package.scala 96:25:@14663.4]
  wire [31:0] _T_1961; // @[Mux.scala 31:69:@14690.4]
  wire  _T_1946; // @[package.scala 96:25:@14654.4 package.scala 96:25:@14655.4]
  wire [31:0] _T_1962; // @[Mux.scala 31:69:@14691.4]
  wire  _T_1943; // @[package.scala 96:25:@14646.4 package.scala 96:25:@14647.4]
  wire [31:0] _T_1963; // @[Mux.scala 31:69:@14692.4]
  wire  _T_1940; // @[package.scala 96:25:@14638.4 package.scala 96:25:@14639.4]
  wire [31:0] _T_1964; // @[Mux.scala 31:69:@14693.4]
  wire  _T_1937; // @[package.scala 96:25:@14630.4 package.scala 96:25:@14631.4]
  wire  _T_2026; // @[package.scala 96:25:@14774.4 package.scala 96:25:@14775.4]
  wire [31:0] _T_2030; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2023; // @[package.scala 96:25:@14766.4 package.scala 96:25:@14767.4]
  wire [31:0] _T_2031; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2020; // @[package.scala 96:25:@14758.4 package.scala 96:25:@14759.4]
  wire [31:0] _T_2032; // @[Mux.scala 31:69:@14786.4]
  wire  _T_2017; // @[package.scala 96:25:@14750.4 package.scala 96:25:@14751.4]
  wire [31:0] _T_2033; // @[Mux.scala 31:69:@14787.4]
  wire  _T_2014; // @[package.scala 96:25:@14742.4 package.scala 96:25:@14743.4]
  wire [31:0] _T_2034; // @[Mux.scala 31:69:@14788.4]
  wire  _T_2011; // @[package.scala 96:25:@14734.4 package.scala 96:25:@14735.4]
  wire [31:0] _T_2035; // @[Mux.scala 31:69:@14789.4]
  wire  _T_2008; // @[package.scala 96:25:@14726.4 package.scala 96:25:@14727.4]
  wire  _T_2097; // @[package.scala 96:25:@14870.4 package.scala 96:25:@14871.4]
  wire [31:0] _T_2101; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2094; // @[package.scala 96:25:@14862.4 package.scala 96:25:@14863.4]
  wire [31:0] _T_2102; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2091; // @[package.scala 96:25:@14854.4 package.scala 96:25:@14855.4]
  wire [31:0] _T_2103; // @[Mux.scala 31:69:@14882.4]
  wire  _T_2088; // @[package.scala 96:25:@14846.4 package.scala 96:25:@14847.4]
  wire [31:0] _T_2104; // @[Mux.scala 31:69:@14883.4]
  wire  _T_2085; // @[package.scala 96:25:@14838.4 package.scala 96:25:@14839.4]
  wire [31:0] _T_2105; // @[Mux.scala 31:69:@14884.4]
  wire  _T_2082; // @[package.scala 96:25:@14830.4 package.scala 96:25:@14831.4]
  wire [31:0] _T_2106; // @[Mux.scala 31:69:@14885.4]
  wire  _T_2079; // @[package.scala 96:25:@14822.4 package.scala 96:25:@14823.4]
  wire  _T_2168; // @[package.scala 96:25:@14966.4 package.scala 96:25:@14967.4]
  wire [31:0] _T_2172; // @[Mux.scala 31:69:@14976.4]
  wire  _T_2165; // @[package.scala 96:25:@14958.4 package.scala 96:25:@14959.4]
  wire [31:0] _T_2173; // @[Mux.scala 31:69:@14977.4]
  wire  _T_2162; // @[package.scala 96:25:@14950.4 package.scala 96:25:@14951.4]
  wire [31:0] _T_2174; // @[Mux.scala 31:69:@14978.4]
  wire  _T_2159; // @[package.scala 96:25:@14942.4 package.scala 96:25:@14943.4]
  wire [31:0] _T_2175; // @[Mux.scala 31:69:@14979.4]
  wire  _T_2156; // @[package.scala 96:25:@14934.4 package.scala 96:25:@14935.4]
  wire [31:0] _T_2176; // @[Mux.scala 31:69:@14980.4]
  wire  _T_2153; // @[package.scala 96:25:@14926.4 package.scala 96:25:@14927.4]
  wire [31:0] _T_2177; // @[Mux.scala 31:69:@14981.4]
  wire  _T_2150; // @[package.scala 96:25:@14918.4 package.scala 96:25:@14919.4]
  wire  _T_2239; // @[package.scala 96:25:@15062.4 package.scala 96:25:@15063.4]
  wire [31:0] _T_2243; // @[Mux.scala 31:69:@15072.4]
  wire  _T_2236; // @[package.scala 96:25:@15054.4 package.scala 96:25:@15055.4]
  wire [31:0] _T_2244; // @[Mux.scala 31:69:@15073.4]
  wire  _T_2233; // @[package.scala 96:25:@15046.4 package.scala 96:25:@15047.4]
  wire [31:0] _T_2245; // @[Mux.scala 31:69:@15074.4]
  wire  _T_2230; // @[package.scala 96:25:@15038.4 package.scala 96:25:@15039.4]
  wire [31:0] _T_2246; // @[Mux.scala 31:69:@15075.4]
  wire  _T_2227; // @[package.scala 96:25:@15030.4 package.scala 96:25:@15031.4]
  wire [31:0] _T_2247; // @[Mux.scala 31:69:@15076.4]
  wire  _T_2224; // @[package.scala 96:25:@15022.4 package.scala 96:25:@15023.4]
  wire [31:0] _T_2248; // @[Mux.scala 31:69:@15077.4]
  wire  _T_2221; // @[package.scala 96:25:@15014.4 package.scala 96:25:@15015.4]
  wire  _T_2310; // @[package.scala 96:25:@15158.4 package.scala 96:25:@15159.4]
  wire [31:0] _T_2314; // @[Mux.scala 31:69:@15168.4]
  wire  _T_2307; // @[package.scala 96:25:@15150.4 package.scala 96:25:@15151.4]
  wire [31:0] _T_2315; // @[Mux.scala 31:69:@15169.4]
  wire  _T_2304; // @[package.scala 96:25:@15142.4 package.scala 96:25:@15143.4]
  wire [31:0] _T_2316; // @[Mux.scala 31:69:@15170.4]
  wire  _T_2301; // @[package.scala 96:25:@15134.4 package.scala 96:25:@15135.4]
  wire [31:0] _T_2317; // @[Mux.scala 31:69:@15171.4]
  wire  _T_2298; // @[package.scala 96:25:@15126.4 package.scala 96:25:@15127.4]
  wire [31:0] _T_2318; // @[Mux.scala 31:69:@15172.4]
  wire  _T_2295; // @[package.scala 96:25:@15118.4 package.scala 96:25:@15119.4]
  wire [31:0] _T_2319; // @[Mux.scala 31:69:@15173.4]
  wire  _T_2292; // @[package.scala 96:25:@15110.4 package.scala 96:25:@15111.4]
  wire  _T_2381; // @[package.scala 96:25:@15254.4 package.scala 96:25:@15255.4]
  wire [31:0] _T_2385; // @[Mux.scala 31:69:@15264.4]
  wire  _T_2378; // @[package.scala 96:25:@15246.4 package.scala 96:25:@15247.4]
  wire [31:0] _T_2386; // @[Mux.scala 31:69:@15265.4]
  wire  _T_2375; // @[package.scala 96:25:@15238.4 package.scala 96:25:@15239.4]
  wire [31:0] _T_2387; // @[Mux.scala 31:69:@15266.4]
  wire  _T_2372; // @[package.scala 96:25:@15230.4 package.scala 96:25:@15231.4]
  wire [31:0] _T_2388; // @[Mux.scala 31:69:@15267.4]
  wire  _T_2369; // @[package.scala 96:25:@15222.4 package.scala 96:25:@15223.4]
  wire [31:0] _T_2389; // @[Mux.scala 31:69:@15268.4]
  wire  _T_2366; // @[package.scala 96:25:@15214.4 package.scala 96:25:@15215.4]
  wire [31:0] _T_2390; // @[Mux.scala 31:69:@15269.4]
  wire  _T_2363; // @[package.scala 96:25:@15206.4 package.scala 96:25:@15207.4]
  wire  _T_2452; // @[package.scala 96:25:@15350.4 package.scala 96:25:@15351.4]
  wire [31:0] _T_2456; // @[Mux.scala 31:69:@15360.4]
  wire  _T_2449; // @[package.scala 96:25:@15342.4 package.scala 96:25:@15343.4]
  wire [31:0] _T_2457; // @[Mux.scala 31:69:@15361.4]
  wire  _T_2446; // @[package.scala 96:25:@15334.4 package.scala 96:25:@15335.4]
  wire [31:0] _T_2458; // @[Mux.scala 31:69:@15362.4]
  wire  _T_2443; // @[package.scala 96:25:@15326.4 package.scala 96:25:@15327.4]
  wire [31:0] _T_2459; // @[Mux.scala 31:69:@15363.4]
  wire  _T_2440; // @[package.scala 96:25:@15318.4 package.scala 96:25:@15319.4]
  wire [31:0] _T_2460; // @[Mux.scala 31:69:@15364.4]
  wire  _T_2437; // @[package.scala 96:25:@15310.4 package.scala 96:25:@15311.4]
  wire [31:0] _T_2461; // @[Mux.scala 31:69:@15365.4]
  wire  _T_2434; // @[package.scala 96:25:@15302.4 package.scala 96:25:@15303.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12776.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12792.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12808.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12824.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12840.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12856.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12872.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12888.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12904.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12920.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12936.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12952.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@12968.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@12984.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@13000.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@13016.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@13248.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@13310.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13372.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13434.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13496.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13558.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13620.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13682.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13744.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13806.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13868.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13930.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@13992.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@14054.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@14116.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@14178.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14241.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14249.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14257.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14265.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14273.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14281.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14289.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14297.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14337.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14345.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14353.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14361.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14369.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14377.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14385.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14393.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14433.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14441.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14449.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14457.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14465.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14473.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14481.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14489.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14529.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14537.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14545.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14553.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14561.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14569.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14577.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14585.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14625.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14633.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14641.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14649.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14657.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14665.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14673.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14681.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14721.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14729.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14737.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14745.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14753.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14761.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14769.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14777.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14817.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14825.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14833.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14841.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14849.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14857.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14865.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14873.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14913.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14921.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14929.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14937.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14945.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14953.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14961.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14969.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@15009.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@15017.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@15025.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@15033.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@15041.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@15049.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@15057.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@15065.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@15105.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@15113.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@15121.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@15129.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@15137.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@15145.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@15153.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15161.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15201.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15209.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15217.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15225.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15233.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15241.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15249.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15257.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15297.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15305.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15313.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15321.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15329.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15337.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15345.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15353.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13032.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@13033.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@13034.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@13035.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13037.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13044.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@13045.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@13046.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@13047.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13049.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@13057.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@13058.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@13059.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13061.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@13069.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@13070.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@13071.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13073.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13080.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@13082.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@13083.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13085.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13092.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@13094.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@13095.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13097.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@13106.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@13107.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13109.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@13118.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@13119.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13121.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13128.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@13130.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@13131.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13133.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13140.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@13142.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@13143.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13145.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@13154.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@13155.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13157.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@13166.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@13167.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13169.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13176.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@13178.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@13179.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13181.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13188.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@13190.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@13191.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13193.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@13202.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@13203.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13205.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@13214.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@13215.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13217.4]
  assign _T_620 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13224.4]
  assign _T_622 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13225.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@13226.4]
  assign _T_626 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13228.4]
  assign _T_628 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13229.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@13230.4]
  assign _T_632 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13232.4]
  assign _T_634 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13233.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@13234.4]
  assign _T_638 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13236.4]
  assign _T_640 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13237.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@13238.4]
  assign _T_644 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13240.4]
  assign _T_646 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13241.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@13242.4]
  assign _T_650 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13244.4]
  assign _T_652 = io_rPort_9_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13245.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@13246.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@13257.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@13258.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@13259.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@13260.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@13261.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@13262.4]
  assign _T_662 = {_T_655,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13264.4]
  assign _T_664 = {_T_656,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13266.4]
  assign _T_666 = {_T_657,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13268.4]
  assign _T_668 = {_T_658,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13270.4]
  assign _T_670 = {_T_659,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13272.4]
  assign _T_672 = {_T_660,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13274.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@13275.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@13276.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@13277.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@13278.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@13279.4]
  assign _T_682 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13286.4]
  assign _T_684 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13287.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_688 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13290.4]
  assign _T_690 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13291.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_694 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13294.4]
  assign _T_696 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13295.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@13296.4]
  assign _T_700 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13298.4]
  assign _T_702 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13299.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@13300.4]
  assign _T_706 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13302.4]
  assign _T_708 = io_rPort_10_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13303.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@13304.4]
  assign _T_712 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13306.4]
  assign _T_714 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13307.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@13308.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@13319.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@13320.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@13321.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@13322.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@13323.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@13324.4]
  assign _T_724 = {_T_717,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13326.4]
  assign _T_726 = {_T_718,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13328.4]
  assign _T_728 = {_T_719,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13330.4]
  assign _T_730 = {_T_720,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_732 = {_T_721,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13334.4]
  assign _T_734 = {_T_722,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13336.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@13337.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@13338.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@13339.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@13340.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@13341.4]
  assign _T_746 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13349.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@13350.4]
  assign _T_752 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13353.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@13354.4]
  assign _T_758 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13357.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@13358.4]
  assign _T_764 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13361.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@13362.4]
  assign _T_770 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13365.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@13366.4]
  assign _T_776 = io_rPort_9_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13369.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@13370.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13381.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13382.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13383.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13384.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13385.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13386.4]
  assign _T_786 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13388.4]
  assign _T_788 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13390.4]
  assign _T_790 = {_T_781,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13392.4]
  assign _T_792 = {_T_782,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13394.4]
  assign _T_794 = {_T_783,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13396.4]
  assign _T_796 = {_T_784,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13398.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@13399.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@13400.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@13401.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@13402.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@13403.4]
  assign _T_808 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13411.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@13412.4]
  assign _T_814 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13415.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@13416.4]
  assign _T_820 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13419.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@13420.4]
  assign _T_826 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13423.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@13424.4]
  assign _T_832 = io_rPort_10_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13427.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@13428.4]
  assign _T_838 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13431.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@13432.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13443.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13444.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13445.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13446.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13447.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13448.4]
  assign _T_848 = {_T_841,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13450.4]
  assign _T_850 = {_T_842,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13452.4]
  assign _T_852 = {_T_843,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13454.4]
  assign _T_854 = {_T_844,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13456.4]
  assign _T_856 = {_T_845,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13458.4]
  assign _T_858 = {_T_846,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13460.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@13461.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@13462.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@13463.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@13464.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@13465.4]
  assign _T_868 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13472.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_874 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13476.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_880 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13480.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@13482.4]
  assign _T_886 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13484.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@13486.4]
  assign _T_892 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13488.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@13490.4]
  assign _T_898 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13492.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@13494.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13505.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13506.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13507.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13508.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13509.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13510.4]
  assign _T_910 = {_T_903,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13512.4]
  assign _T_912 = {_T_904,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13514.4]
  assign _T_914 = {_T_905,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13516.4]
  assign _T_916 = {_T_906,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13518.4]
  assign _T_918 = {_T_907,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13520.4]
  assign _T_920 = {_T_908,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13522.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@13523.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@13524.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@13525.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@13526.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@13527.4]
  assign _T_930 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13534.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@13536.4]
  assign _T_936 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13538.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@13540.4]
  assign _T_942 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13542.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@13544.4]
  assign _T_948 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13546.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@13548.4]
  assign _T_954 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13550.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@13552.4]
  assign _T_960 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13554.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@13556.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13567.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13568.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13569.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13570.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13571.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13572.4]
  assign _T_972 = {_T_965,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13574.4]
  assign _T_974 = {_T_966,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13576.4]
  assign _T_976 = {_T_967,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13578.4]
  assign _T_978 = {_T_968,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13580.4]
  assign _T_980 = {_T_969,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13582.4]
  assign _T_982 = {_T_970,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13584.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@13585.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@13586.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@13587.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@13588.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@13589.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@13598.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@13602.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@13606.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@13610.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@13614.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@13618.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13629.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13630.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13631.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13632.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13633.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13634.4]
  assign _T_1034 = {_T_1027,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13636.4]
  assign _T_1036 = {_T_1028,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13638.4]
  assign _T_1038 = {_T_1029,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13640.4]
  assign _T_1040 = {_T_1030,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13642.4]
  assign _T_1042 = {_T_1031,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13644.4]
  assign _T_1044 = {_T_1032,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13646.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@13647.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@13648.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@13649.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@13650.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@13651.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@13668.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@13672.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@13676.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@13680.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13691.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13692.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13693.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13694.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13695.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13696.4]
  assign _T_1096 = {_T_1089,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13698.4]
  assign _T_1098 = {_T_1090,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13700.4]
  assign _T_1100 = {_T_1091,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13702.4]
  assign _T_1102 = {_T_1092,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13704.4]
  assign _T_1104 = {_T_1093,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13706.4]
  assign _T_1106 = {_T_1094,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13708.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@13709.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@13710.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@13711.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@13712.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@13713.4]
  assign _T_1116 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13720.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@13722.4]
  assign _T_1122 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13724.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@13726.4]
  assign _T_1128 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13728.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@13730.4]
  assign _T_1134 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13732.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@13734.4]
  assign _T_1140 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13736.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@13738.4]
  assign _T_1146 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13740.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@13742.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13753.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13754.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13755.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13756.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13757.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13758.4]
  assign _T_1158 = {_T_1151,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13760.4]
  assign _T_1160 = {_T_1152,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13762.4]
  assign _T_1162 = {_T_1153,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13764.4]
  assign _T_1164 = {_T_1154,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13766.4]
  assign _T_1166 = {_T_1155,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13768.4]
  assign _T_1168 = {_T_1156,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13770.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@13771.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@13772.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@13773.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@13774.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@13775.4]
  assign _T_1178 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13782.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@13784.4]
  assign _T_1184 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13786.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@13788.4]
  assign _T_1190 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13790.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@13792.4]
  assign _T_1196 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13794.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@13796.4]
  assign _T_1202 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13798.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@13800.4]
  assign _T_1208 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13802.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@13804.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13815.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13816.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13817.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13818.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13819.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13820.4]
  assign _T_1220 = {_T_1213,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13822.4]
  assign _T_1222 = {_T_1214,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13824.4]
  assign _T_1224 = {_T_1215,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13826.4]
  assign _T_1226 = {_T_1216,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13828.4]
  assign _T_1228 = {_T_1217,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13830.4]
  assign _T_1230 = {_T_1218,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13832.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@13833.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@13834.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@13835.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@13836.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@13837.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@13846.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@13850.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@13854.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@13858.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@13862.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@13866.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13877.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13878.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13879.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13880.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13881.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13882.4]
  assign _T_1282 = {_T_1275,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13884.4]
  assign _T_1284 = {_T_1276,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13886.4]
  assign _T_1286 = {_T_1277,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13888.4]
  assign _T_1288 = {_T_1278,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13890.4]
  assign _T_1290 = {_T_1279,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13892.4]
  assign _T_1292 = {_T_1280,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13894.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@13895.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@13896.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@13897.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@13898.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@13899.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@13908.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@13912.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@13916.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@13920.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@13924.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@13928.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13939.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13940.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13941.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13942.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13943.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13944.4]
  assign _T_1344 = {_T_1337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13946.4]
  assign _T_1346 = {_T_1338,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13948.4]
  assign _T_1348 = {_T_1339,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13950.4]
  assign _T_1350 = {_T_1340,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13952.4]
  assign _T_1352 = {_T_1341,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13954.4]
  assign _T_1354 = {_T_1342,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13956.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@13957.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@13958.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@13959.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@13960.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@13961.4]
  assign _T_1364 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13968.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@13970.4]
  assign _T_1370 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13972.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@13974.4]
  assign _T_1376 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13976.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@13978.4]
  assign _T_1382 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13980.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@13982.4]
  assign _T_1388 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13984.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@13986.4]
  assign _T_1394 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13988.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@13990.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@14001.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@14002.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@14003.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@14004.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@14005.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@14006.4]
  assign _T_1406 = {_T_1399,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14008.4]
  assign _T_1408 = {_T_1400,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14010.4]
  assign _T_1410 = {_T_1401,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14012.4]
  assign _T_1412 = {_T_1402,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14014.4]
  assign _T_1414 = {_T_1403,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14016.4]
  assign _T_1416 = {_T_1404,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14018.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@14019.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@14020.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@14021.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@14022.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@14023.4]
  assign _T_1426 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14030.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@14032.4]
  assign _T_1432 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14034.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@14036.4]
  assign _T_1438 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14038.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@14040.4]
  assign _T_1444 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14042.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@14044.4]
  assign _T_1450 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14046.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@14048.4]
  assign _T_1456 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14050.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@14052.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@14063.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@14064.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@14065.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@14066.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@14067.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@14068.4]
  assign _T_1468 = {_T_1461,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14070.4]
  assign _T_1470 = {_T_1462,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14072.4]
  assign _T_1472 = {_T_1463,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14074.4]
  assign _T_1474 = {_T_1464,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14076.4]
  assign _T_1476 = {_T_1465,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14078.4]
  assign _T_1478 = {_T_1466,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14080.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@14081.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@14082.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@14083.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@14084.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@14085.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@14094.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@14098.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@14102.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@14106.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@14110.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@14114.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@14125.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@14126.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@14127.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@14128.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@14129.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@14130.4]
  assign _T_1530 = {_T_1523,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14132.4]
  assign _T_1532 = {_T_1524,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14134.4]
  assign _T_1534 = {_T_1525,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14136.4]
  assign _T_1536 = {_T_1526,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14138.4]
  assign _T_1538 = {_T_1527,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14140.4]
  assign _T_1540 = {_T_1528,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14142.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@14143.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@14144.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@14145.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@14146.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@14147.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@14156.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@14160.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@14164.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@14168.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@14172.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@14176.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@14187.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@14188.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@14189.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@14190.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@14191.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@14192.4]
  assign _T_1592 = {_T_1585,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14194.4]
  assign _T_1594 = {_T_1586,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14196.4]
  assign _T_1596 = {_T_1587,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14198.4]
  assign _T_1598 = {_T_1588,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14200.4]
  assign _T_1600 = {_T_1589,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14202.4]
  assign _T_1602 = {_T_1590,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14204.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@14205.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@14206.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@14207.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@14208.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@14209.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14294.4 package.scala 96:25:@14295.4]
  assign _T_1675 = _T_1671 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14304.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14286.4 package.scala 96:25:@14287.4]
  assign _T_1676 = _T_1668 ? Mem1D_11_io_output : _T_1675; // @[Mux.scala 31:69:@14305.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14278.4 package.scala 96:25:@14279.4]
  assign _T_1677 = _T_1665 ? Mem1D_9_io_output : _T_1676; // @[Mux.scala 31:69:@14306.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14270.4 package.scala 96:25:@14271.4]
  assign _T_1678 = _T_1662 ? Mem1D_7_io_output : _T_1677; // @[Mux.scala 31:69:@14307.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14262.4 package.scala 96:25:@14263.4]
  assign _T_1679 = _T_1659 ? Mem1D_5_io_output : _T_1678; // @[Mux.scala 31:69:@14308.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14254.4 package.scala 96:25:@14255.4]
  assign _T_1680 = _T_1656 ? Mem1D_3_io_output : _T_1679; // @[Mux.scala 31:69:@14309.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@14246.4 package.scala 96:25:@14247.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14390.4 package.scala 96:25:@14391.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14400.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14382.4 package.scala 96:25:@14383.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@14401.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14374.4 package.scala 96:25:@14375.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@14402.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@14366.4 package.scala 96:25:@14367.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@14403.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14358.4 package.scala 96:25:@14359.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@14404.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14350.4 package.scala 96:25:@14351.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@14405.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14342.4 package.scala 96:25:@14343.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14486.4 package.scala 96:25:@14487.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14496.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14478.4 package.scala 96:25:@14479.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@14497.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14470.4 package.scala 96:25:@14471.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@14498.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14462.4 package.scala 96:25:@14463.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@14499.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14454.4 package.scala 96:25:@14455.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@14500.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14446.4 package.scala 96:25:@14447.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@14501.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14438.4 package.scala 96:25:@14439.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14582.4 package.scala 96:25:@14583.4]
  assign _T_1888 = _T_1884 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14592.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14574.4 package.scala 96:25:@14575.4]
  assign _T_1889 = _T_1881 ? Mem1D_10_io_output : _T_1888; // @[Mux.scala 31:69:@14593.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14566.4 package.scala 96:25:@14567.4]
  assign _T_1890 = _T_1878 ? Mem1D_8_io_output : _T_1889; // @[Mux.scala 31:69:@14594.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14558.4 package.scala 96:25:@14559.4]
  assign _T_1891 = _T_1875 ? Mem1D_6_io_output : _T_1890; // @[Mux.scala 31:69:@14595.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14550.4 package.scala 96:25:@14551.4]
  assign _T_1892 = _T_1872 ? Mem1D_4_io_output : _T_1891; // @[Mux.scala 31:69:@14596.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14542.4 package.scala 96:25:@14543.4]
  assign _T_1893 = _T_1869 ? Mem1D_2_io_output : _T_1892; // @[Mux.scala 31:69:@14597.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14534.4 package.scala 96:25:@14535.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14678.4 package.scala 96:25:@14679.4]
  assign _T_1959 = _T_1955 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14688.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14670.4 package.scala 96:25:@14671.4]
  assign _T_1960 = _T_1952 ? Mem1D_11_io_output : _T_1959; // @[Mux.scala 31:69:@14689.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14662.4 package.scala 96:25:@14663.4]
  assign _T_1961 = _T_1949 ? Mem1D_9_io_output : _T_1960; // @[Mux.scala 31:69:@14690.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@14654.4 package.scala 96:25:@14655.4]
  assign _T_1962 = _T_1946 ? Mem1D_7_io_output : _T_1961; // @[Mux.scala 31:69:@14691.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14646.4 package.scala 96:25:@14647.4]
  assign _T_1963 = _T_1943 ? Mem1D_5_io_output : _T_1962; // @[Mux.scala 31:69:@14692.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14638.4 package.scala 96:25:@14639.4]
  assign _T_1964 = _T_1940 ? Mem1D_3_io_output : _T_1963; // @[Mux.scala 31:69:@14693.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14630.4 package.scala 96:25:@14631.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14774.4 package.scala 96:25:@14775.4]
  assign _T_2030 = _T_2026 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14784.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14766.4 package.scala 96:25:@14767.4]
  assign _T_2031 = _T_2023 ? Mem1D_11_io_output : _T_2030; // @[Mux.scala 31:69:@14785.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14758.4 package.scala 96:25:@14759.4]
  assign _T_2032 = _T_2020 ? Mem1D_9_io_output : _T_2031; // @[Mux.scala 31:69:@14786.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14750.4 package.scala 96:25:@14751.4]
  assign _T_2033 = _T_2017 ? Mem1D_7_io_output : _T_2032; // @[Mux.scala 31:69:@14787.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14742.4 package.scala 96:25:@14743.4]
  assign _T_2034 = _T_2014 ? Mem1D_5_io_output : _T_2033; // @[Mux.scala 31:69:@14788.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14734.4 package.scala 96:25:@14735.4]
  assign _T_2035 = _T_2011 ? Mem1D_3_io_output : _T_2034; // @[Mux.scala 31:69:@14789.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14726.4 package.scala 96:25:@14727.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14870.4 package.scala 96:25:@14871.4]
  assign _T_2101 = _T_2097 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14880.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14862.4 package.scala 96:25:@14863.4]
  assign _T_2102 = _T_2094 ? Mem1D_10_io_output : _T_2101; // @[Mux.scala 31:69:@14881.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14854.4 package.scala 96:25:@14855.4]
  assign _T_2103 = _T_2091 ? Mem1D_8_io_output : _T_2102; // @[Mux.scala 31:69:@14882.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14846.4 package.scala 96:25:@14847.4]
  assign _T_2104 = _T_2088 ? Mem1D_6_io_output : _T_2103; // @[Mux.scala 31:69:@14883.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14838.4 package.scala 96:25:@14839.4]
  assign _T_2105 = _T_2085 ? Mem1D_4_io_output : _T_2104; // @[Mux.scala 31:69:@14884.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14830.4 package.scala 96:25:@14831.4]
  assign _T_2106 = _T_2082 ? Mem1D_2_io_output : _T_2105; // @[Mux.scala 31:69:@14885.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14822.4 package.scala 96:25:@14823.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14966.4 package.scala 96:25:@14967.4]
  assign _T_2172 = _T_2168 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14976.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14958.4 package.scala 96:25:@14959.4]
  assign _T_2173 = _T_2165 ? Mem1D_10_io_output : _T_2172; // @[Mux.scala 31:69:@14977.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14950.4 package.scala 96:25:@14951.4]
  assign _T_2174 = _T_2162 ? Mem1D_8_io_output : _T_2173; // @[Mux.scala 31:69:@14978.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14942.4 package.scala 96:25:@14943.4]
  assign _T_2175 = _T_2159 ? Mem1D_6_io_output : _T_2174; // @[Mux.scala 31:69:@14979.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14934.4 package.scala 96:25:@14935.4]
  assign _T_2176 = _T_2156 ? Mem1D_4_io_output : _T_2175; // @[Mux.scala 31:69:@14980.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14926.4 package.scala 96:25:@14927.4]
  assign _T_2177 = _T_2153 ? Mem1D_2_io_output : _T_2176; // @[Mux.scala 31:69:@14981.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14918.4 package.scala 96:25:@14919.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@15062.4 package.scala 96:25:@15063.4]
  assign _T_2243 = _T_2239 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15072.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@15054.4 package.scala 96:25:@15055.4]
  assign _T_2244 = _T_2236 ? Mem1D_10_io_output : _T_2243; // @[Mux.scala 31:69:@15073.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@15046.4 package.scala 96:25:@15047.4]
  assign _T_2245 = _T_2233 ? Mem1D_8_io_output : _T_2244; // @[Mux.scala 31:69:@15074.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@15038.4 package.scala 96:25:@15039.4]
  assign _T_2246 = _T_2230 ? Mem1D_6_io_output : _T_2245; // @[Mux.scala 31:69:@15075.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@15030.4 package.scala 96:25:@15031.4]
  assign _T_2247 = _T_2227 ? Mem1D_4_io_output : _T_2246; // @[Mux.scala 31:69:@15076.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@15022.4 package.scala 96:25:@15023.4]
  assign _T_2248 = _T_2224 ? Mem1D_2_io_output : _T_2247; // @[Mux.scala 31:69:@15077.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@15014.4 package.scala 96:25:@15015.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15158.4 package.scala 96:25:@15159.4]
  assign _T_2314 = _T_2310 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15168.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@15150.4 package.scala 96:25:@15151.4]
  assign _T_2315 = _T_2307 ? Mem1D_10_io_output : _T_2314; // @[Mux.scala 31:69:@15169.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@15142.4 package.scala 96:25:@15143.4]
  assign _T_2316 = _T_2304 ? Mem1D_8_io_output : _T_2315; // @[Mux.scala 31:69:@15170.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@15134.4 package.scala 96:25:@15135.4]
  assign _T_2317 = _T_2301 ? Mem1D_6_io_output : _T_2316; // @[Mux.scala 31:69:@15171.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@15126.4 package.scala 96:25:@15127.4]
  assign _T_2318 = _T_2298 ? Mem1D_4_io_output : _T_2317; // @[Mux.scala 31:69:@15172.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@15118.4 package.scala 96:25:@15119.4]
  assign _T_2319 = _T_2295 ? Mem1D_2_io_output : _T_2318; // @[Mux.scala 31:69:@15173.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@15110.4 package.scala 96:25:@15111.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15254.4 package.scala 96:25:@15255.4]
  assign _T_2385 = _T_2381 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15264.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15246.4 package.scala 96:25:@15247.4]
  assign _T_2386 = _T_2378 ? Mem1D_11_io_output : _T_2385; // @[Mux.scala 31:69:@15265.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15238.4 package.scala 96:25:@15239.4]
  assign _T_2387 = _T_2375 ? Mem1D_9_io_output : _T_2386; // @[Mux.scala 31:69:@15266.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@15230.4 package.scala 96:25:@15231.4]
  assign _T_2388 = _T_2372 ? Mem1D_7_io_output : _T_2387; // @[Mux.scala 31:69:@15267.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15222.4 package.scala 96:25:@15223.4]
  assign _T_2389 = _T_2369 ? Mem1D_5_io_output : _T_2388; // @[Mux.scala 31:69:@15268.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15214.4 package.scala 96:25:@15215.4]
  assign _T_2390 = _T_2366 ? Mem1D_3_io_output : _T_2389; // @[Mux.scala 31:69:@15269.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15206.4 package.scala 96:25:@15207.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15350.4 package.scala 96:25:@15351.4]
  assign _T_2456 = _T_2452 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15360.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15342.4 package.scala 96:25:@15343.4]
  assign _T_2457 = _T_2449 ? Mem1D_11_io_output : _T_2456; // @[Mux.scala 31:69:@15361.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15334.4 package.scala 96:25:@15335.4]
  assign _T_2458 = _T_2446 ? Mem1D_9_io_output : _T_2457; // @[Mux.scala 31:69:@15362.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15326.4 package.scala 96:25:@15327.4]
  assign _T_2459 = _T_2443 ? Mem1D_7_io_output : _T_2458; // @[Mux.scala 31:69:@15363.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15318.4 package.scala 96:25:@15319.4]
  assign _T_2460 = _T_2440 ? Mem1D_5_io_output : _T_2459; // @[Mux.scala 31:69:@15364.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15310.4 package.scala 96:25:@15311.4]
  assign _T_2461 = _T_2437 ? Mem1D_3_io_output : _T_2460; // @[Mux.scala 31:69:@15365.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15302.4 package.scala 96:25:@15303.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_1_io_output : _T_2461; // @[MemPrimitives.scala 152:13:@15367.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_1_io_output : _T_2390; // @[MemPrimitives.scala 152:13:@15271.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_io_output : _T_2319; // @[MemPrimitives.scala 152:13:@15175.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_io_output : _T_2248; // @[MemPrimitives.scala 152:13:@15079.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_io_output : _T_2177; // @[MemPrimitives.scala 152:13:@14983.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_io_output : _T_2106; // @[MemPrimitives.scala 152:13:@14887.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_1_io_output : _T_2035; // @[MemPrimitives.scala 152:13:@14791.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_1_io_output : _T_1964; // @[MemPrimitives.scala 152:13:@14695.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_io_output : _T_1893; // @[MemPrimitives.scala 152:13:@14599.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 152:13:@14503.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 152:13:@14407.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_1_io_output : _T_1680; // @[MemPrimitives.scala 152:13:@14311.4]
  assign Mem1D_clock = clock; // @[:@12777.4]
  assign Mem1D_reset = reset; // @[:@12778.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 131:28:@13283.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 132:32:@13284.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@13041.4]
  assign Mem1D_io_w_data_0 = _T_450[40:9]; // @[MemPrimitives.scala 95:29:@13042.4]
  assign Mem1D_io_w_en_0 = _T_450[41]; // @[MemPrimitives.scala 96:27:@13043.4]
  assign Mem1D_1_clock = clock; // @[:@12793.4]
  assign Mem1D_1_reset = reset; // @[:@12794.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 131:28:@13345.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 132:32:@13346.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@13053.4]
  assign Mem1D_1_io_w_data_0 = _T_461[40:9]; // @[MemPrimitives.scala 95:29:@13054.4]
  assign Mem1D_1_io_w_en_0 = _T_461[41]; // @[MemPrimitives.scala 96:27:@13055.4]
  assign Mem1D_2_clock = clock; // @[:@12809.4]
  assign Mem1D_2_reset = reset; // @[:@12810.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 131:28:@13407.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 132:32:@13408.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@13065.4]
  assign Mem1D_2_io_w_data_0 = _T_472[40:9]; // @[MemPrimitives.scala 95:29:@13066.4]
  assign Mem1D_2_io_w_en_0 = _T_472[41]; // @[MemPrimitives.scala 96:27:@13067.4]
  assign Mem1D_3_clock = clock; // @[:@12825.4]
  assign Mem1D_3_reset = reset; // @[:@12826.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 131:28:@13469.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 132:32:@13470.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@13077.4]
  assign Mem1D_3_io_w_data_0 = _T_483[40:9]; // @[MemPrimitives.scala 95:29:@13078.4]
  assign Mem1D_3_io_w_en_0 = _T_483[41]; // @[MemPrimitives.scala 96:27:@13079.4]
  assign Mem1D_4_clock = clock; // @[:@12841.4]
  assign Mem1D_4_reset = reset; // @[:@12842.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 131:28:@13531.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 132:32:@13532.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@13089.4]
  assign Mem1D_4_io_w_data_0 = _T_494[40:9]; // @[MemPrimitives.scala 95:29:@13090.4]
  assign Mem1D_4_io_w_en_0 = _T_494[41]; // @[MemPrimitives.scala 96:27:@13091.4]
  assign Mem1D_5_clock = clock; // @[:@12857.4]
  assign Mem1D_5_reset = reset; // @[:@12858.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 131:28:@13593.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 132:32:@13594.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@13101.4]
  assign Mem1D_5_io_w_data_0 = _T_505[40:9]; // @[MemPrimitives.scala 95:29:@13102.4]
  assign Mem1D_5_io_w_en_0 = _T_505[41]; // @[MemPrimitives.scala 96:27:@13103.4]
  assign Mem1D_6_clock = clock; // @[:@12873.4]
  assign Mem1D_6_reset = reset; // @[:@12874.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 131:28:@13655.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 132:32:@13656.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@13113.4]
  assign Mem1D_6_io_w_data_0 = _T_516[40:9]; // @[MemPrimitives.scala 95:29:@13114.4]
  assign Mem1D_6_io_w_en_0 = _T_516[41]; // @[MemPrimitives.scala 96:27:@13115.4]
  assign Mem1D_7_clock = clock; // @[:@12889.4]
  assign Mem1D_7_reset = reset; // @[:@12890.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 131:28:@13717.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 132:32:@13718.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@13125.4]
  assign Mem1D_7_io_w_data_0 = _T_527[40:9]; // @[MemPrimitives.scala 95:29:@13126.4]
  assign Mem1D_7_io_w_en_0 = _T_527[41]; // @[MemPrimitives.scala 96:27:@13127.4]
  assign Mem1D_8_clock = clock; // @[:@12905.4]
  assign Mem1D_8_reset = reset; // @[:@12906.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 131:28:@13779.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 132:32:@13780.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@13137.4]
  assign Mem1D_8_io_w_data_0 = _T_538[40:9]; // @[MemPrimitives.scala 95:29:@13138.4]
  assign Mem1D_8_io_w_en_0 = _T_538[41]; // @[MemPrimitives.scala 96:27:@13139.4]
  assign Mem1D_9_clock = clock; // @[:@12921.4]
  assign Mem1D_9_reset = reset; // @[:@12922.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 131:28:@13841.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 132:32:@13842.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@13149.4]
  assign Mem1D_9_io_w_data_0 = _T_549[40:9]; // @[MemPrimitives.scala 95:29:@13150.4]
  assign Mem1D_9_io_w_en_0 = _T_549[41]; // @[MemPrimitives.scala 96:27:@13151.4]
  assign Mem1D_10_clock = clock; // @[:@12937.4]
  assign Mem1D_10_reset = reset; // @[:@12938.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 131:28:@13903.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 132:32:@13904.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@13161.4]
  assign Mem1D_10_io_w_data_0 = _T_560[40:9]; // @[MemPrimitives.scala 95:29:@13162.4]
  assign Mem1D_10_io_w_en_0 = _T_560[41]; // @[MemPrimitives.scala 96:27:@13163.4]
  assign Mem1D_11_clock = clock; // @[:@12953.4]
  assign Mem1D_11_reset = reset; // @[:@12954.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@13965.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@13966.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@13173.4]
  assign Mem1D_11_io_w_data_0 = _T_571[40:9]; // @[MemPrimitives.scala 95:29:@13174.4]
  assign Mem1D_11_io_w_en_0 = _T_571[41]; // @[MemPrimitives.scala 96:27:@13175.4]
  assign Mem1D_12_clock = clock; // @[:@12969.4]
  assign Mem1D_12_reset = reset; // @[:@12970.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 131:28:@14027.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 132:32:@14028.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@13185.4]
  assign Mem1D_12_io_w_data_0 = _T_582[40:9]; // @[MemPrimitives.scala 95:29:@13186.4]
  assign Mem1D_12_io_w_en_0 = _T_582[41]; // @[MemPrimitives.scala 96:27:@13187.4]
  assign Mem1D_13_clock = clock; // @[:@12985.4]
  assign Mem1D_13_reset = reset; // @[:@12986.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 131:28:@14089.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 132:32:@14090.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@13197.4]
  assign Mem1D_13_io_w_data_0 = _T_593[40:9]; // @[MemPrimitives.scala 95:29:@13198.4]
  assign Mem1D_13_io_w_en_0 = _T_593[41]; // @[MemPrimitives.scala 96:27:@13199.4]
  assign Mem1D_14_clock = clock; // @[:@13001.4]
  assign Mem1D_14_reset = reset; // @[:@13002.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 131:28:@14151.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 132:32:@14152.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@13209.4]
  assign Mem1D_14_io_w_data_0 = _T_604[40:9]; // @[MemPrimitives.scala 95:29:@13210.4]
  assign Mem1D_14_io_w_en_0 = _T_604[41]; // @[MemPrimitives.scala 96:27:@13211.4]
  assign Mem1D_15_clock = clock; // @[:@13017.4]
  assign Mem1D_15_reset = reset; // @[:@13018.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 131:28:@14213.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 132:32:@14214.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@13221.4]
  assign Mem1D_15_io_w_data_0 = _T_615[40:9]; // @[MemPrimitives.scala 95:29:@13222.4]
  assign Mem1D_15_io_w_en_0 = _T_615[41]; // @[MemPrimitives.scala 96:27:@13223.4]
  assign StickySelects_clock = clock; // @[:@13249.4]
  assign StickySelects_reset = reset; // @[:@13250.4]
  assign StickySelects_io_ins_0 = io_rPort_2_en_0 & _T_623; // @[MemPrimitives.scala 125:64:@13251.4]
  assign StickySelects_io_ins_1 = io_rPort_3_en_0 & _T_629; // @[MemPrimitives.scala 125:64:@13252.4]
  assign StickySelects_io_ins_2 = io_rPort_6_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13253.4]
  assign StickySelects_io_ins_3 = io_rPort_7_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13254.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13255.4]
  assign StickySelects_io_ins_5 = io_rPort_9_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13256.4]
  assign StickySelects_1_clock = clock; // @[:@13311.4]
  assign StickySelects_1_reset = reset; // @[:@13312.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@13313.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@13314.4]
  assign StickySelects_1_io_ins_2 = io_rPort_4_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@13315.4]
  assign StickySelects_1_io_ins_3 = io_rPort_5_en_0 & _T_703; // @[MemPrimitives.scala 125:64:@13316.4]
  assign StickySelects_1_io_ins_4 = io_rPort_10_en_0 & _T_709; // @[MemPrimitives.scala 125:64:@13317.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_715; // @[MemPrimitives.scala 125:64:@13318.4]
  assign StickySelects_2_clock = clock; // @[:@13373.4]
  assign StickySelects_2_reset = reset; // @[:@13374.4]
  assign StickySelects_2_io_ins_0 = io_rPort_2_en_0 & _T_747; // @[MemPrimitives.scala 125:64:@13375.4]
  assign StickySelects_2_io_ins_1 = io_rPort_3_en_0 & _T_753; // @[MemPrimitives.scala 125:64:@13376.4]
  assign StickySelects_2_io_ins_2 = io_rPort_6_en_0 & _T_759; // @[MemPrimitives.scala 125:64:@13377.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_765; // @[MemPrimitives.scala 125:64:@13378.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_771; // @[MemPrimitives.scala 125:64:@13379.4]
  assign StickySelects_2_io_ins_5 = io_rPort_9_en_0 & _T_777; // @[MemPrimitives.scala 125:64:@13380.4]
  assign StickySelects_3_clock = clock; // @[:@13435.4]
  assign StickySelects_3_reset = reset; // @[:@13436.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_809; // @[MemPrimitives.scala 125:64:@13437.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_815; // @[MemPrimitives.scala 125:64:@13438.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_821; // @[MemPrimitives.scala 125:64:@13439.4]
  assign StickySelects_3_io_ins_3 = io_rPort_5_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@13440.4]
  assign StickySelects_3_io_ins_4 = io_rPort_10_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@13441.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_839; // @[MemPrimitives.scala 125:64:@13442.4]
  assign StickySelects_4_clock = clock; // @[:@13497.4]
  assign StickySelects_4_reset = reset; // @[:@13498.4]
  assign StickySelects_4_io_ins_0 = io_rPort_2_en_0 & _T_871; // @[MemPrimitives.scala 125:64:@13499.4]
  assign StickySelects_4_io_ins_1 = io_rPort_3_en_0 & _T_877; // @[MemPrimitives.scala 125:64:@13500.4]
  assign StickySelects_4_io_ins_2 = io_rPort_6_en_0 & _T_883; // @[MemPrimitives.scala 125:64:@13501.4]
  assign StickySelects_4_io_ins_3 = io_rPort_7_en_0 & _T_889; // @[MemPrimitives.scala 125:64:@13502.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_895; // @[MemPrimitives.scala 125:64:@13503.4]
  assign StickySelects_4_io_ins_5 = io_rPort_9_en_0 & _T_901; // @[MemPrimitives.scala 125:64:@13504.4]
  assign StickySelects_5_clock = clock; // @[:@13559.4]
  assign StickySelects_5_reset = reset; // @[:@13560.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_933; // @[MemPrimitives.scala 125:64:@13561.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_939; // @[MemPrimitives.scala 125:64:@13562.4]
  assign StickySelects_5_io_ins_2 = io_rPort_4_en_0 & _T_945; // @[MemPrimitives.scala 125:64:@13563.4]
  assign StickySelects_5_io_ins_3 = io_rPort_5_en_0 & _T_951; // @[MemPrimitives.scala 125:64:@13564.4]
  assign StickySelects_5_io_ins_4 = io_rPort_10_en_0 & _T_957; // @[MemPrimitives.scala 125:64:@13565.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_963; // @[MemPrimitives.scala 125:64:@13566.4]
  assign StickySelects_6_clock = clock; // @[:@13621.4]
  assign StickySelects_6_reset = reset; // @[:@13622.4]
  assign StickySelects_6_io_ins_0 = io_rPort_2_en_0 & _T_995; // @[MemPrimitives.scala 125:64:@13623.4]
  assign StickySelects_6_io_ins_1 = io_rPort_3_en_0 & _T_1001; // @[MemPrimitives.scala 125:64:@13624.4]
  assign StickySelects_6_io_ins_2 = io_rPort_6_en_0 & _T_1007; // @[MemPrimitives.scala 125:64:@13625.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1013; // @[MemPrimitives.scala 125:64:@13626.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1019; // @[MemPrimitives.scala 125:64:@13627.4]
  assign StickySelects_6_io_ins_5 = io_rPort_9_en_0 & _T_1025; // @[MemPrimitives.scala 125:64:@13628.4]
  assign StickySelects_7_clock = clock; // @[:@13683.4]
  assign StickySelects_7_reset = reset; // @[:@13684.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1057; // @[MemPrimitives.scala 125:64:@13685.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1063; // @[MemPrimitives.scala 125:64:@13686.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_1069; // @[MemPrimitives.scala 125:64:@13687.4]
  assign StickySelects_7_io_ins_3 = io_rPort_5_en_0 & _T_1075; // @[MemPrimitives.scala 125:64:@13688.4]
  assign StickySelects_7_io_ins_4 = io_rPort_10_en_0 & _T_1081; // @[MemPrimitives.scala 125:64:@13689.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1087; // @[MemPrimitives.scala 125:64:@13690.4]
  assign StickySelects_8_clock = clock; // @[:@13745.4]
  assign StickySelects_8_reset = reset; // @[:@13746.4]
  assign StickySelects_8_io_ins_0 = io_rPort_2_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13747.4]
  assign StickySelects_8_io_ins_1 = io_rPort_3_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13748.4]
  assign StickySelects_8_io_ins_2 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13749.4]
  assign StickySelects_8_io_ins_3 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13750.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13751.4]
  assign StickySelects_8_io_ins_5 = io_rPort_9_en_0 & _T_1149; // @[MemPrimitives.scala 125:64:@13752.4]
  assign StickySelects_9_clock = clock; // @[:@13807.4]
  assign StickySelects_9_reset = reset; // @[:@13808.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1181; // @[MemPrimitives.scala 125:64:@13809.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13810.4]
  assign StickySelects_9_io_ins_2 = io_rPort_4_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13811.4]
  assign StickySelects_9_io_ins_3 = io_rPort_5_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13812.4]
  assign StickySelects_9_io_ins_4 = io_rPort_10_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13813.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13814.4]
  assign StickySelects_10_clock = clock; // @[:@13869.4]
  assign StickySelects_10_reset = reset; // @[:@13870.4]
  assign StickySelects_10_io_ins_0 = io_rPort_2_en_0 & _T_1243; // @[MemPrimitives.scala 125:64:@13871.4]
  assign StickySelects_10_io_ins_1 = io_rPort_3_en_0 & _T_1249; // @[MemPrimitives.scala 125:64:@13872.4]
  assign StickySelects_10_io_ins_2 = io_rPort_6_en_0 & _T_1255; // @[MemPrimitives.scala 125:64:@13873.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_1261; // @[MemPrimitives.scala 125:64:@13874.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_1267; // @[MemPrimitives.scala 125:64:@13875.4]
  assign StickySelects_10_io_ins_5 = io_rPort_9_en_0 & _T_1273; // @[MemPrimitives.scala 125:64:@13876.4]
  assign StickySelects_11_clock = clock; // @[:@13931.4]
  assign StickySelects_11_reset = reset; // @[:@13932.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@13933.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@13934.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@13935.4]
  assign StickySelects_11_io_ins_3 = io_rPort_5_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@13936.4]
  assign StickySelects_11_io_ins_4 = io_rPort_10_en_0 & _T_1329; // @[MemPrimitives.scala 125:64:@13937.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1335; // @[MemPrimitives.scala 125:64:@13938.4]
  assign StickySelects_12_clock = clock; // @[:@13993.4]
  assign StickySelects_12_reset = reset; // @[:@13994.4]
  assign StickySelects_12_io_ins_0 = io_rPort_2_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@13995.4]
  assign StickySelects_12_io_ins_1 = io_rPort_3_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@13996.4]
  assign StickySelects_12_io_ins_2 = io_rPort_6_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@13997.4]
  assign StickySelects_12_io_ins_3 = io_rPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@13998.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@13999.4]
  assign StickySelects_12_io_ins_5 = io_rPort_9_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@14000.4]
  assign StickySelects_13_clock = clock; // @[:@14055.4]
  assign StickySelects_13_reset = reset; // @[:@14056.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1429; // @[MemPrimitives.scala 125:64:@14057.4]
  assign StickySelects_13_io_ins_1 = io_rPort_1_en_0 & _T_1435; // @[MemPrimitives.scala 125:64:@14058.4]
  assign StickySelects_13_io_ins_2 = io_rPort_4_en_0 & _T_1441; // @[MemPrimitives.scala 125:64:@14059.4]
  assign StickySelects_13_io_ins_3 = io_rPort_5_en_0 & _T_1447; // @[MemPrimitives.scala 125:64:@14060.4]
  assign StickySelects_13_io_ins_4 = io_rPort_10_en_0 & _T_1453; // @[MemPrimitives.scala 125:64:@14061.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@14062.4]
  assign StickySelects_14_clock = clock; // @[:@14117.4]
  assign StickySelects_14_reset = reset; // @[:@14118.4]
  assign StickySelects_14_io_ins_0 = io_rPort_2_en_0 & _T_1491; // @[MemPrimitives.scala 125:64:@14119.4]
  assign StickySelects_14_io_ins_1 = io_rPort_3_en_0 & _T_1497; // @[MemPrimitives.scala 125:64:@14120.4]
  assign StickySelects_14_io_ins_2 = io_rPort_6_en_0 & _T_1503; // @[MemPrimitives.scala 125:64:@14121.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_1509; // @[MemPrimitives.scala 125:64:@14122.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_1515; // @[MemPrimitives.scala 125:64:@14123.4]
  assign StickySelects_14_io_ins_5 = io_rPort_9_en_0 & _T_1521; // @[MemPrimitives.scala 125:64:@14124.4]
  assign StickySelects_15_clock = clock; // @[:@14179.4]
  assign StickySelects_15_reset = reset; // @[:@14180.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1553; // @[MemPrimitives.scala 125:64:@14181.4]
  assign StickySelects_15_io_ins_1 = io_rPort_1_en_0 & _T_1559; // @[MemPrimitives.scala 125:64:@14182.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_1565; // @[MemPrimitives.scala 125:64:@14183.4]
  assign StickySelects_15_io_ins_3 = io_rPort_5_en_0 & _T_1571; // @[MemPrimitives.scala 125:64:@14184.4]
  assign StickySelects_15_io_ins_4 = io_rPort_10_en_0 & _T_1577; // @[MemPrimitives.scala 125:64:@14185.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1583; // @[MemPrimitives.scala 125:64:@14186.4]
  assign RetimeWrapper_clock = clock; // @[:@14242.4]
  assign RetimeWrapper_reset = reset; // @[:@14243.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14245.4]
  assign RetimeWrapper_io_in = _T_685 & io_rPort_0_en_0; // @[package.scala 94:16:@14244.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14250.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14251.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14253.4]
  assign RetimeWrapper_1_io_in = _T_809 & io_rPort_0_en_0; // @[package.scala 94:16:@14252.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14258.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14259.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14261.4]
  assign RetimeWrapper_2_io_in = _T_933 & io_rPort_0_en_0; // @[package.scala 94:16:@14260.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14266.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14267.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14269.4]
  assign RetimeWrapper_3_io_in = _T_1057 & io_rPort_0_en_0; // @[package.scala 94:16:@14268.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14274.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14275.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14277.4]
  assign RetimeWrapper_4_io_in = _T_1181 & io_rPort_0_en_0; // @[package.scala 94:16:@14276.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14282.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14283.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14285.4]
  assign RetimeWrapper_5_io_in = _T_1305 & io_rPort_0_en_0; // @[package.scala 94:16:@14284.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14290.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14291.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14293.4]
  assign RetimeWrapper_6_io_in = _T_1429 & io_rPort_0_en_0; // @[package.scala 94:16:@14292.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14298.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14299.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14301.4]
  assign RetimeWrapper_7_io_in = _T_1553 & io_rPort_0_en_0; // @[package.scala 94:16:@14300.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14338.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14339.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14341.4]
  assign RetimeWrapper_8_io_in = _T_691 & io_rPort_1_en_0; // @[package.scala 94:16:@14340.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14346.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14347.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14349.4]
  assign RetimeWrapper_9_io_in = _T_815 & io_rPort_1_en_0; // @[package.scala 94:16:@14348.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14354.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14355.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14357.4]
  assign RetimeWrapper_10_io_in = _T_939 & io_rPort_1_en_0; // @[package.scala 94:16:@14356.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14362.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14363.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14365.4]
  assign RetimeWrapper_11_io_in = _T_1063 & io_rPort_1_en_0; // @[package.scala 94:16:@14364.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14370.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14371.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14373.4]
  assign RetimeWrapper_12_io_in = _T_1187 & io_rPort_1_en_0; // @[package.scala 94:16:@14372.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14378.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14379.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14381.4]
  assign RetimeWrapper_13_io_in = _T_1311 & io_rPort_1_en_0; // @[package.scala 94:16:@14380.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14386.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14387.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14389.4]
  assign RetimeWrapper_14_io_in = _T_1435 & io_rPort_1_en_0; // @[package.scala 94:16:@14388.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14394.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14395.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14397.4]
  assign RetimeWrapper_15_io_in = _T_1559 & io_rPort_1_en_0; // @[package.scala 94:16:@14396.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14434.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14435.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14437.4]
  assign RetimeWrapper_16_io_in = _T_623 & io_rPort_2_en_0; // @[package.scala 94:16:@14436.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14442.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14443.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14445.4]
  assign RetimeWrapper_17_io_in = _T_747 & io_rPort_2_en_0; // @[package.scala 94:16:@14444.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14450.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14451.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14453.4]
  assign RetimeWrapper_18_io_in = _T_871 & io_rPort_2_en_0; // @[package.scala 94:16:@14452.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14458.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14459.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14461.4]
  assign RetimeWrapper_19_io_in = _T_995 & io_rPort_2_en_0; // @[package.scala 94:16:@14460.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14466.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14467.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14469.4]
  assign RetimeWrapper_20_io_in = _T_1119 & io_rPort_2_en_0; // @[package.scala 94:16:@14468.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14474.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14475.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14477.4]
  assign RetimeWrapper_21_io_in = _T_1243 & io_rPort_2_en_0; // @[package.scala 94:16:@14476.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14482.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14483.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14485.4]
  assign RetimeWrapper_22_io_in = _T_1367 & io_rPort_2_en_0; // @[package.scala 94:16:@14484.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14490.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14491.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14493.4]
  assign RetimeWrapper_23_io_in = _T_1491 & io_rPort_2_en_0; // @[package.scala 94:16:@14492.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14530.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14531.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14533.4]
  assign RetimeWrapper_24_io_in = _T_629 & io_rPort_3_en_0; // @[package.scala 94:16:@14532.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14538.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14539.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14541.4]
  assign RetimeWrapper_25_io_in = _T_753 & io_rPort_3_en_0; // @[package.scala 94:16:@14540.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14546.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14547.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14549.4]
  assign RetimeWrapper_26_io_in = _T_877 & io_rPort_3_en_0; // @[package.scala 94:16:@14548.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14554.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14555.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14557.4]
  assign RetimeWrapper_27_io_in = _T_1001 & io_rPort_3_en_0; // @[package.scala 94:16:@14556.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14562.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14563.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14565.4]
  assign RetimeWrapper_28_io_in = _T_1125 & io_rPort_3_en_0; // @[package.scala 94:16:@14564.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14570.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14571.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14573.4]
  assign RetimeWrapper_29_io_in = _T_1249 & io_rPort_3_en_0; // @[package.scala 94:16:@14572.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14578.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14579.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14581.4]
  assign RetimeWrapper_30_io_in = _T_1373 & io_rPort_3_en_0; // @[package.scala 94:16:@14580.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14586.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14587.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14589.4]
  assign RetimeWrapper_31_io_in = _T_1497 & io_rPort_3_en_0; // @[package.scala 94:16:@14588.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14626.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14627.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14629.4]
  assign RetimeWrapper_32_io_in = _T_697 & io_rPort_4_en_0; // @[package.scala 94:16:@14628.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14634.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14635.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14637.4]
  assign RetimeWrapper_33_io_in = _T_821 & io_rPort_4_en_0; // @[package.scala 94:16:@14636.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14642.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14643.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14645.4]
  assign RetimeWrapper_34_io_in = _T_945 & io_rPort_4_en_0; // @[package.scala 94:16:@14644.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14650.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14651.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14653.4]
  assign RetimeWrapper_35_io_in = _T_1069 & io_rPort_4_en_0; // @[package.scala 94:16:@14652.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14658.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14659.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14661.4]
  assign RetimeWrapper_36_io_in = _T_1193 & io_rPort_4_en_0; // @[package.scala 94:16:@14660.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14666.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14667.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14669.4]
  assign RetimeWrapper_37_io_in = _T_1317 & io_rPort_4_en_0; // @[package.scala 94:16:@14668.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14674.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14675.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14677.4]
  assign RetimeWrapper_38_io_in = _T_1441 & io_rPort_4_en_0; // @[package.scala 94:16:@14676.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14682.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14683.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14685.4]
  assign RetimeWrapper_39_io_in = _T_1565 & io_rPort_4_en_0; // @[package.scala 94:16:@14684.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14722.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14723.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14725.4]
  assign RetimeWrapper_40_io_in = _T_703 & io_rPort_5_en_0; // @[package.scala 94:16:@14724.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14730.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14731.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14733.4]
  assign RetimeWrapper_41_io_in = _T_827 & io_rPort_5_en_0; // @[package.scala 94:16:@14732.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14738.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14739.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14741.4]
  assign RetimeWrapper_42_io_in = _T_951 & io_rPort_5_en_0; // @[package.scala 94:16:@14740.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14746.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14747.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14749.4]
  assign RetimeWrapper_43_io_in = _T_1075 & io_rPort_5_en_0; // @[package.scala 94:16:@14748.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14754.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14755.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14757.4]
  assign RetimeWrapper_44_io_in = _T_1199 & io_rPort_5_en_0; // @[package.scala 94:16:@14756.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14762.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14763.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14765.4]
  assign RetimeWrapper_45_io_in = _T_1323 & io_rPort_5_en_0; // @[package.scala 94:16:@14764.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14770.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14771.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14773.4]
  assign RetimeWrapper_46_io_in = _T_1447 & io_rPort_5_en_0; // @[package.scala 94:16:@14772.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14778.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14779.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14781.4]
  assign RetimeWrapper_47_io_in = _T_1571 & io_rPort_5_en_0; // @[package.scala 94:16:@14780.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14818.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14819.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14821.4]
  assign RetimeWrapper_48_io_in = _T_635 & io_rPort_6_en_0; // @[package.scala 94:16:@14820.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14826.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14827.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14829.4]
  assign RetimeWrapper_49_io_in = _T_759 & io_rPort_6_en_0; // @[package.scala 94:16:@14828.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14834.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14835.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14837.4]
  assign RetimeWrapper_50_io_in = _T_883 & io_rPort_6_en_0; // @[package.scala 94:16:@14836.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14842.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14843.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14845.4]
  assign RetimeWrapper_51_io_in = _T_1007 & io_rPort_6_en_0; // @[package.scala 94:16:@14844.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14850.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14851.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14853.4]
  assign RetimeWrapper_52_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@14852.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14858.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14859.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14861.4]
  assign RetimeWrapper_53_io_in = _T_1255 & io_rPort_6_en_0; // @[package.scala 94:16:@14860.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14866.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14867.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14869.4]
  assign RetimeWrapper_54_io_in = _T_1379 & io_rPort_6_en_0; // @[package.scala 94:16:@14868.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14874.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14875.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14877.4]
  assign RetimeWrapper_55_io_in = _T_1503 & io_rPort_6_en_0; // @[package.scala 94:16:@14876.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14914.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14915.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14917.4]
  assign RetimeWrapper_56_io_in = _T_641 & io_rPort_7_en_0; // @[package.scala 94:16:@14916.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14922.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14923.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14925.4]
  assign RetimeWrapper_57_io_in = _T_765 & io_rPort_7_en_0; // @[package.scala 94:16:@14924.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14930.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14931.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14933.4]
  assign RetimeWrapper_58_io_in = _T_889 & io_rPort_7_en_0; // @[package.scala 94:16:@14932.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14938.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14939.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14941.4]
  assign RetimeWrapper_59_io_in = _T_1013 & io_rPort_7_en_0; // @[package.scala 94:16:@14940.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14946.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14947.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14949.4]
  assign RetimeWrapper_60_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@14948.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14954.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14955.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14957.4]
  assign RetimeWrapper_61_io_in = _T_1261 & io_rPort_7_en_0; // @[package.scala 94:16:@14956.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14962.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14963.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14965.4]
  assign RetimeWrapper_62_io_in = _T_1385 & io_rPort_7_en_0; // @[package.scala 94:16:@14964.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14970.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14971.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14973.4]
  assign RetimeWrapper_63_io_in = _T_1509 & io_rPort_7_en_0; // @[package.scala 94:16:@14972.4]
  assign RetimeWrapper_64_clock = clock; // @[:@15010.4]
  assign RetimeWrapper_64_reset = reset; // @[:@15011.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15013.4]
  assign RetimeWrapper_64_io_in = _T_647 & io_rPort_8_en_0; // @[package.scala 94:16:@15012.4]
  assign RetimeWrapper_65_clock = clock; // @[:@15018.4]
  assign RetimeWrapper_65_reset = reset; // @[:@15019.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15021.4]
  assign RetimeWrapper_65_io_in = _T_771 & io_rPort_8_en_0; // @[package.scala 94:16:@15020.4]
  assign RetimeWrapper_66_clock = clock; // @[:@15026.4]
  assign RetimeWrapper_66_reset = reset; // @[:@15027.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15029.4]
  assign RetimeWrapper_66_io_in = _T_895 & io_rPort_8_en_0; // @[package.scala 94:16:@15028.4]
  assign RetimeWrapper_67_clock = clock; // @[:@15034.4]
  assign RetimeWrapper_67_reset = reset; // @[:@15035.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15037.4]
  assign RetimeWrapper_67_io_in = _T_1019 & io_rPort_8_en_0; // @[package.scala 94:16:@15036.4]
  assign RetimeWrapper_68_clock = clock; // @[:@15042.4]
  assign RetimeWrapper_68_reset = reset; // @[:@15043.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15045.4]
  assign RetimeWrapper_68_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15044.4]
  assign RetimeWrapper_69_clock = clock; // @[:@15050.4]
  assign RetimeWrapper_69_reset = reset; // @[:@15051.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15053.4]
  assign RetimeWrapper_69_io_in = _T_1267 & io_rPort_8_en_0; // @[package.scala 94:16:@15052.4]
  assign RetimeWrapper_70_clock = clock; // @[:@15058.4]
  assign RetimeWrapper_70_reset = reset; // @[:@15059.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15061.4]
  assign RetimeWrapper_70_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@15060.4]
  assign RetimeWrapper_71_clock = clock; // @[:@15066.4]
  assign RetimeWrapper_71_reset = reset; // @[:@15067.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15069.4]
  assign RetimeWrapper_71_io_in = _T_1515 & io_rPort_8_en_0; // @[package.scala 94:16:@15068.4]
  assign RetimeWrapper_72_clock = clock; // @[:@15106.4]
  assign RetimeWrapper_72_reset = reset; // @[:@15107.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15109.4]
  assign RetimeWrapper_72_io_in = _T_653 & io_rPort_9_en_0; // @[package.scala 94:16:@15108.4]
  assign RetimeWrapper_73_clock = clock; // @[:@15114.4]
  assign RetimeWrapper_73_reset = reset; // @[:@15115.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15117.4]
  assign RetimeWrapper_73_io_in = _T_777 & io_rPort_9_en_0; // @[package.scala 94:16:@15116.4]
  assign RetimeWrapper_74_clock = clock; // @[:@15122.4]
  assign RetimeWrapper_74_reset = reset; // @[:@15123.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15125.4]
  assign RetimeWrapper_74_io_in = _T_901 & io_rPort_9_en_0; // @[package.scala 94:16:@15124.4]
  assign RetimeWrapper_75_clock = clock; // @[:@15130.4]
  assign RetimeWrapper_75_reset = reset; // @[:@15131.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15133.4]
  assign RetimeWrapper_75_io_in = _T_1025 & io_rPort_9_en_0; // @[package.scala 94:16:@15132.4]
  assign RetimeWrapper_76_clock = clock; // @[:@15138.4]
  assign RetimeWrapper_76_reset = reset; // @[:@15139.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15141.4]
  assign RetimeWrapper_76_io_in = _T_1149 & io_rPort_9_en_0; // @[package.scala 94:16:@15140.4]
  assign RetimeWrapper_77_clock = clock; // @[:@15146.4]
  assign RetimeWrapper_77_reset = reset; // @[:@15147.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15149.4]
  assign RetimeWrapper_77_io_in = _T_1273 & io_rPort_9_en_0; // @[package.scala 94:16:@15148.4]
  assign RetimeWrapper_78_clock = clock; // @[:@15154.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15155.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15157.4]
  assign RetimeWrapper_78_io_in = _T_1397 & io_rPort_9_en_0; // @[package.scala 94:16:@15156.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15162.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15163.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15165.4]
  assign RetimeWrapper_79_io_in = _T_1521 & io_rPort_9_en_0; // @[package.scala 94:16:@15164.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15202.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15203.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15205.4]
  assign RetimeWrapper_80_io_in = _T_709 & io_rPort_10_en_0; // @[package.scala 94:16:@15204.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15210.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15211.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15213.4]
  assign RetimeWrapper_81_io_in = _T_833 & io_rPort_10_en_0; // @[package.scala 94:16:@15212.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15218.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15219.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15221.4]
  assign RetimeWrapper_82_io_in = _T_957 & io_rPort_10_en_0; // @[package.scala 94:16:@15220.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15226.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15227.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15229.4]
  assign RetimeWrapper_83_io_in = _T_1081 & io_rPort_10_en_0; // @[package.scala 94:16:@15228.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15234.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15235.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15237.4]
  assign RetimeWrapper_84_io_in = _T_1205 & io_rPort_10_en_0; // @[package.scala 94:16:@15236.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15242.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15243.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15245.4]
  assign RetimeWrapper_85_io_in = _T_1329 & io_rPort_10_en_0; // @[package.scala 94:16:@15244.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15250.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15251.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15253.4]
  assign RetimeWrapper_86_io_in = _T_1453 & io_rPort_10_en_0; // @[package.scala 94:16:@15252.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15258.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15259.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15261.4]
  assign RetimeWrapper_87_io_in = _T_1577 & io_rPort_10_en_0; // @[package.scala 94:16:@15260.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15298.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15299.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15301.4]
  assign RetimeWrapper_88_io_in = _T_715 & io_rPort_11_en_0; // @[package.scala 94:16:@15300.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15306.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15307.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15309.4]
  assign RetimeWrapper_89_io_in = _T_839 & io_rPort_11_en_0; // @[package.scala 94:16:@15308.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15314.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15315.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15317.4]
  assign RetimeWrapper_90_io_in = _T_963 & io_rPort_11_en_0; // @[package.scala 94:16:@15316.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15322.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15323.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15325.4]
  assign RetimeWrapper_91_io_in = _T_1087 & io_rPort_11_en_0; // @[package.scala 94:16:@15324.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15330.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15331.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15333.4]
  assign RetimeWrapper_92_io_in = _T_1211 & io_rPort_11_en_0; // @[package.scala 94:16:@15332.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15338.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15339.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15341.4]
  assign RetimeWrapper_93_io_in = _T_1335 & io_rPort_11_en_0; // @[package.scala 94:16:@15340.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15346.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15347.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15349.4]
  assign RetimeWrapper_94_io_in = _T_1459 & io_rPort_11_en_0; // @[package.scala 94:16:@15348.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15354.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15355.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15357.4]
  assign RetimeWrapper_95_io_in = _T_1583 & io_rPort_11_en_0; // @[package.scala 94:16:@15356.4]
endmodule
module RetimeWrapper_168( // @[:@15772.2]
  input         clock, // @[:@15773.4]
  input         reset, // @[:@15774.4]
  input         io_flow, // @[:@15775.4]
  input  [31:0] io_in, // @[:@15775.4]
  output [31:0] io_out // @[:@15775.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15777.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15790.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15789.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15788.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15787.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15786.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15784.4]
endmodule
module RetimeWrapper_169( // @[:@15804.2]
  input         clock, // @[:@15805.4]
  input         reset, // @[:@15806.4]
  input         io_flow, // @[:@15807.4]
  input  [31:0] io_in, // @[:@15807.4]
  output [31:0] io_out // @[:@15807.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15809.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15822.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15821.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15820.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15819.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15818.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15816.4]
endmodule
module RetimeWrapper_170( // @[:@15836.2]
  input   clock, // @[:@15837.4]
  input   reset, // @[:@15838.4]
  input   io_flow, // @[:@15839.4]
  input   io_in, // @[:@15839.4]
  output  io_out // @[:@15839.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15841.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15841.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15854.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15853.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15852.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15851.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15850.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15848.4]
endmodule
module RetimeWrapper_181( // @[:@16482.2]
  input         clock, // @[:@16483.4]
  input         reset, // @[:@16484.4]
  input         io_flow, // @[:@16485.4]
  input  [31:0] io_in, // @[:@16485.4]
  output [31:0] io_out // @[:@16485.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@16487.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16500.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16499.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16498.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16497.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16496.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16494.4]
endmodule
module RetimeWrapper_184( // @[:@16578.2]
  input         clock, // @[:@16579.4]
  input         reset, // @[:@16580.4]
  input         io_flow, // @[:@16581.4]
  input  [31:0] io_in, // @[:@16581.4]
  output [31:0] io_out // @[:@16581.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16583.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16596.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16595.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16594.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16593.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16592.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16590.4]
endmodule
module RetimeWrapper_186( // @[:@16642.2]
  input   clock, // @[:@16643.4]
  input   reset, // @[:@16644.4]
  input   io_flow, // @[:@16645.4]
  input   io_in, // @[:@16645.4]
  output  io_out // @[:@16645.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16647.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16660.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16659.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@16658.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16657.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16656.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16654.4]
endmodule
module RetimeWrapper_187( // @[:@16674.2]
  input         clock, // @[:@16675.4]
  input         reset, // @[:@16676.4]
  input         io_flow, // @[:@16677.4]
  input  [31:0] io_in, // @[:@16677.4]
  output [31:0] io_out // @[:@16677.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@16679.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16692.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16691.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16690.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16689.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16688.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16686.4]
endmodule
module RetimeWrapper_189( // @[:@16738.2]
  input         clock, // @[:@16739.4]
  input         reset, // @[:@16740.4]
  input         io_flow, // @[:@16741.4]
  input  [31:0] io_in, // @[:@16741.4]
  output [31:0] io_out // @[:@16741.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16743.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@16743.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16756.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16755.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16754.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16753.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16752.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16750.4]
endmodule
module RetimeWrapper_244( // @[:@20854.2]
  input         clock, // @[:@20855.4]
  input         reset, // @[:@20856.4]
  input         io_flow, // @[:@20857.4]
  input  [32:0] io_in, // @[:@20857.4]
  output [32:0] io_out // @[:@20857.4]
);
  wire [32:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20859.4]
  wire [32:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20859.4]
  wire [32:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20859.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20859.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20859.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20859.4]
  RetimeShiftRegister #(.WIDTH(33), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@20859.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20872.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20871.4]
  assign sr_init = 33'h0; // @[RetimeShiftRegister.scala 19:16:@20870.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20869.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20868.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20866.4]
endmodule
module RetimeWrapper_246( // @[:@20918.2]
  input         clock, // @[:@20919.4]
  input         reset, // @[:@20920.4]
  input         io_flow, // @[:@20921.4]
  input  [33:0] io_in, // @[:@20921.4]
  output [33:0] io_out // @[:@20921.4]
);
  wire [33:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20923.4]
  wire [33:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20923.4]
  wire [33:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20923.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20923.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20923.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20923.4]
  RetimeShiftRegister #(.WIDTH(34), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@20923.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20936.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20935.4]
  assign sr_init = 34'h0; // @[RetimeShiftRegister.scala 19:16:@20934.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20933.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20932.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20930.4]
endmodule
module fix2fixBox_84( // @[:@21034.2]
  input  [31:0] io_a, // @[:@21037.4]
  output [32:0] io_b // @[:@21037.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@21051.4]
endmodule
module __56( // @[:@21053.2]
  input  [31:0] io_b, // @[:@21056.4]
  output [32:0] io_result // @[:@21056.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@21061.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@21061.4]
  fix2fixBox_84 fix2fixBox ( // @[BigIPZynq.scala 219:30:@21061.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@21069.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@21064.4]
endmodule
module x394_x13( // @[:@21165.2]
  input         clock, // @[:@21166.4]
  input         reset, // @[:@21167.4]
  input  [31:0] io_a, // @[:@21168.4]
  input  [31:0] io_b, // @[:@21168.4]
  input         io_flow, // @[:@21168.4]
  output [31:0] io_result // @[:@21168.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@21176.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@21176.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@21183.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@21183.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@21193.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@21193.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@21193.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@21193.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@21193.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@21181.4 Math.scala 724:14:@21182.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@21188.4 Math.scala 724:14:@21189.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@21190.4]
  __56 _ ( // @[Math.scala 720:24:@21176.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __56 __1 ( // @[Math.scala 720:24:@21183.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@21193.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@21181.4 Math.scala 724:14:@21182.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@21188.4 Math.scala 724:14:@21189.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@21190.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@21201.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@21179.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@21186.4]
  assign fix2fixBox_clock = clock; // @[:@21194.4]
  assign fix2fixBox_reset = reset; // @[:@21195.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@21196.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@21199.4]
endmodule
module RetimeWrapper_259( // @[:@22293.2]
  input         clock, // @[:@22294.4]
  input         reset, // @[:@22295.4]
  input         io_flow, // @[:@22296.4]
  input  [31:0] io_in, // @[:@22296.4]
  output [31:0] io_out // @[:@22296.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22298.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22298.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22298.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22298.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22298.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22298.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@22298.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22311.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22310.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22309.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22308.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22307.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22305.4]
endmodule
module fix2fixBox_108( // @[:@22482.2]
  input  [31:0] io_a, // @[:@22485.4]
  output [31:0] io_b // @[:@22485.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@22495.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@22495.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@22498.4]
endmodule
module x402( // @[:@22500.2]
  input  [31:0] io_b, // @[:@22503.4]
  output [31:0] io_result // @[:@22503.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@22508.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@22508.4]
  fix2fixBox_108 fix2fixBox ( // @[BigIPZynq.scala 219:30:@22508.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@22516.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@22511.4]
endmodule
module Multiplier( // @[:@22528.2]
  input         clock, // @[:@22529.4]
  input         io_flow, // @[:@22531.4]
  input  [38:0] io_a, // @[:@22531.4]
  input  [38:0] io_b, // @[:@22531.4]
  output [38:0] io_out // @[:@22531.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@22533.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@22533.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@22533.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@22533.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@22533.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@22533.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@22543.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@22541.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@22540.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@22542.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@22539.4]
endmodule
module fix2fixBox_109( // @[:@22545.2]
  input  [38:0] io_a, // @[:@22548.4]
  output [31:0] io_b // @[:@22548.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@22556.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@22559.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@22556.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@22559.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@22562.4]
endmodule
module x403_mul( // @[:@22564.2]
  input         clock, // @[:@22565.4]
  input  [31:0] io_a, // @[:@22567.4]
  input  [31:0] io_b, // @[:@22567.4]
  input         io_flow, // @[:@22567.4]
  output [31:0] io_result // @[:@22567.4]
);
  wire  x403_mul_clock; // @[BigIPZynq.scala 63:21:@22582.4]
  wire  x403_mul_io_flow; // @[BigIPZynq.scala 63:21:@22582.4]
  wire [38:0] x403_mul_io_a; // @[BigIPZynq.scala 63:21:@22582.4]
  wire [38:0] x403_mul_io_b; // @[BigIPZynq.scala 63:21:@22582.4]
  wire [38:0] x403_mul_io_out; // @[BigIPZynq.scala 63:21:@22582.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@22590.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@22590.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@22574.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@22576.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@22578.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@22580.4]
  Multiplier x403_mul ( // @[BigIPZynq.scala 63:21:@22582.4]
    .clock(x403_mul_clock),
    .io_flow(x403_mul_io_flow),
    .io_a(x403_mul_io_a),
    .io_b(x403_mul_io_b),
    .io_out(x403_mul_io_out)
  );
  fix2fixBox_109 fix2fixBox ( // @[Math.scala 253:30:@22590.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@22574.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@22576.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@22578.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@22580.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@22598.4]
  assign x403_mul_clock = clock; // @[:@22583.4]
  assign x403_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@22587.4]
  assign x403_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@22585.4]
  assign x403_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@22586.4]
  assign fix2fixBox_io_a = x403_mul_io_out; // @[Math.scala 254:23:@22593.4]
endmodule
module fix2fixBox_110( // @[:@22600.2]
  input  [31:0] io_a, // @[:@22603.4]
  output [31:0] io_b // @[:@22603.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@22615.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@22615.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@22618.4]
endmodule
module x404( // @[:@22620.2]
  input  [31:0] io_b, // @[:@22623.4]
  output [31:0] io_result // @[:@22623.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@22628.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@22628.4]
  fix2fixBox_110 fix2fixBox ( // @[BigIPZynq.scala 219:30:@22628.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@22636.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@22631.4]
endmodule
module RetimeWrapper_261( // @[:@22650.2]
  input         clock, // @[:@22651.4]
  input         reset, // @[:@22652.4]
  input         io_flow, // @[:@22653.4]
  input  [31:0] io_in, // @[:@22653.4]
  output [31:0] io_out // @[:@22653.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22655.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22655.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22655.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22655.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22655.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22655.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@22655.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22668.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22667.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22666.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22665.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22664.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22662.4]
endmodule
module x405_sub( // @[:@22801.2]
  input         clock, // @[:@22802.4]
  input         reset, // @[:@22803.4]
  input  [31:0] io_a, // @[:@22804.4]
  input  [31:0] io_b, // @[:@22804.4]
  input         io_flow, // @[:@22804.4]
  output [31:0] io_result // @[:@22804.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@22812.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@22812.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@22819.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@22819.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@22830.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@22830.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@22830.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@22830.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@22830.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@22817.4 Math.scala 724:14:@22818.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@22824.4 Math.scala 724:14:@22825.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@22826.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@22827.4]
  __56 _ ( // @[Math.scala 720:24:@22812.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __56 __1 ( // @[Math.scala 720:24:@22819.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@22830.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@22817.4 Math.scala 724:14:@22818.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@22824.4 Math.scala 724:14:@22825.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@22826.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@22827.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@22838.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@22815.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@22822.4]
  assign fix2fixBox_clock = clock; // @[:@22831.4]
  assign fix2fixBox_reset = reset; // @[:@22832.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@22833.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@22836.4]
endmodule
module RetimeWrapper_265( // @[:@23210.2]
  input         clock, // @[:@23211.4]
  input         reset, // @[:@23212.4]
  input         io_flow, // @[:@23213.4]
  input  [31:0] io_in, // @[:@23213.4]
  output [31:0] io_out // @[:@23213.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23215.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23215.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23215.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23215.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23215.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23215.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@23215.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23228.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23227.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@23226.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23225.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23224.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23222.4]
endmodule
module RetimeWrapper_290( // @[:@25968.2]
  input         clock, // @[:@25969.4]
  input         reset, // @[:@25970.4]
  input         io_flow, // @[:@25971.4]
  input  [63:0] io_in, // @[:@25971.4]
  output [63:0] io_out // @[:@25971.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25973.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25973.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25973.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@25973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25985.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@25984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25980.4]
endmodule
module x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@26084.2]
  input          clock, // @[:@26085.4]
  input          reset, // @[:@26086.4]
  output         io_in_x253_TREADY, // @[:@26087.4]
  input  [255:0] io_in_x253_TDATA, // @[:@26087.4]
  input  [7:0]   io_in_x253_TID, // @[:@26087.4]
  input  [7:0]   io_in_x253_TDEST, // @[:@26087.4]
  output         io_in_x254_TVALID, // @[:@26087.4]
  input          io_in_x254_TREADY, // @[:@26087.4]
  output [255:0] io_in_x254_TDATA, // @[:@26087.4]
  input          io_sigsIn_backpressure, // @[:@26087.4]
  input          io_sigsIn_datapathEn, // @[:@26087.4]
  input          io_sigsIn_break, // @[:@26087.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@26087.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@26087.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@26087.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@26087.4]
  input          io_rr // @[:@26087.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@26101.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@26101.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@26113.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@26113.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26136.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26136.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26136.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@26136.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@26136.4]
  wire  x290_lb_0_clock; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_reset; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_11_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_11_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_11_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_11_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_11_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_11_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_10_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_10_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_10_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_10_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_10_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_10_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_9_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_9_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_9_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_9_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_9_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_9_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_8_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_8_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_8_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_8_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_8_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_8_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_7_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_7_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_7_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_7_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_7_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_7_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_6_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_6_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_6_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_6_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_6_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_6_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_5_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_5_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_5_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_5_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_5_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_5_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_4_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_4_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_4_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_4_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_4_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_4_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_3_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_3_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_3_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_3_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_3_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_3_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_2_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_2_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_2_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_2_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_2_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_2_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_1_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_1_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_1_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_1_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_1_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_1_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_0_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_rPort_0_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_rPort_0_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_0_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_rPort_0_backpressure; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_rPort_0_output_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_wPort_1_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_wPort_1_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_wPort_1_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_wPort_1_data_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_wPort_1_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_wPort_0_banks_1; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [2:0] x290_lb_0_io_wPort_0_banks_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [8:0] x290_lb_0_io_wPort_0_ofs_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire [31:0] x290_lb_0_io_wPort_0_data_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x290_lb_0_io_wPort_0_en_0; // @[m_x290_lb_0.scala 39:17:@26146.4]
  wire  x508_sub_1_clock; // @[Math.scala 191:24:@26309.4]
  wire  x508_sub_1_reset; // @[Math.scala 191:24:@26309.4]
  wire [31:0] x508_sub_1_io_a; // @[Math.scala 191:24:@26309.4]
  wire [31:0] x508_sub_1_io_b; // @[Math.scala 191:24:@26309.4]
  wire  x508_sub_1_io_flow; // @[Math.scala 191:24:@26309.4]
  wire [31:0] x508_sub_1_io_result; // @[Math.scala 191:24:@26309.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@26336.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@26336.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@26336.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@26336.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@26336.4]
  wire  x299_sum_1_clock; // @[Math.scala 150:24:@26345.4]
  wire  x299_sum_1_reset; // @[Math.scala 150:24:@26345.4]
  wire [31:0] x299_sum_1_io_a; // @[Math.scala 150:24:@26345.4]
  wire [31:0] x299_sum_1_io_b; // @[Math.scala 150:24:@26345.4]
  wire  x299_sum_1_io_flow; // @[Math.scala 150:24:@26345.4]
  wire [31:0] x299_sum_1_io_result; // @[Math.scala 150:24:@26345.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@26355.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@26355.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@26355.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@26355.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@26355.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@26364.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@26364.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@26364.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@26364.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@26364.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@26373.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@26373.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@26373.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@26373.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@26373.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@26382.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@26382.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@26382.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@26382.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@26382.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@26391.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@26391.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@26391.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@26391.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@26391.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@26400.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@26400.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@26400.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@26400.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@26400.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@26411.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@26411.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@26411.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@26411.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@26411.4]
  wire  x301_rdcol_1_clock; // @[Math.scala 150:24:@26434.4]
  wire  x301_rdcol_1_reset; // @[Math.scala 150:24:@26434.4]
  wire [31:0] x301_rdcol_1_io_a; // @[Math.scala 150:24:@26434.4]
  wire [31:0] x301_rdcol_1_io_b; // @[Math.scala 150:24:@26434.4]
  wire  x301_rdcol_1_io_flow; // @[Math.scala 150:24:@26434.4]
  wire [31:0] x301_rdcol_1_io_result; // @[Math.scala 150:24:@26434.4]
  wire  x305_sum_1_clock; // @[Math.scala 150:24:@26474.4]
  wire  x305_sum_1_reset; // @[Math.scala 150:24:@26474.4]
  wire [31:0] x305_sum_1_io_a; // @[Math.scala 150:24:@26474.4]
  wire [31:0] x305_sum_1_io_b; // @[Math.scala 150:24:@26474.4]
  wire  x305_sum_1_io_flow; // @[Math.scala 150:24:@26474.4]
  wire [31:0] x305_sum_1_io_result; // @[Math.scala 150:24:@26474.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@26484.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@26484.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@26484.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@26484.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@26484.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@26493.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@26493.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@26493.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@26493.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@26493.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@26502.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@26502.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@26502.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@26502.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@26502.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@26513.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@26513.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@26513.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@26513.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@26513.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@26534.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@26534.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@26534.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@26534.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@26534.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@26550.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@26550.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@26550.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@26550.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@26550.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@26581.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@26581.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@26581.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@26581.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@26581.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@26590.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@26590.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@26590.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@26590.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@26590.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@26599.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@26599.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@26599.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@26599.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@26599.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@26608.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@26608.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@26608.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@26608.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@26608.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@26626.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@26626.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@26626.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@26626.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@26626.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@26638.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@26638.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@26638.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@26638.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@26638.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@26659.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@26659.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@26659.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@26659.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@26659.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@26683.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@26683.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@26683.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@26683.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@26683.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@26692.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@26692.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@26692.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@26692.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@26692.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@26701.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@26701.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@26701.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@26701.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@26701.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@26713.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@26713.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@26713.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@26713.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@26713.4]
  wire  x319_rdcol_1_clock; // @[Math.scala 150:24:@26736.4]
  wire  x319_rdcol_1_reset; // @[Math.scala 150:24:@26736.4]
  wire [31:0] x319_rdcol_1_io_a; // @[Math.scala 150:24:@26736.4]
  wire [31:0] x319_rdcol_1_io_b; // @[Math.scala 150:24:@26736.4]
  wire  x319_rdcol_1_io_flow; // @[Math.scala 150:24:@26736.4]
  wire [31:0] x319_rdcol_1_io_result; // @[Math.scala 150:24:@26736.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@26787.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@26787.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@26787.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@26787.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@26787.4]
  wire  x325_sum_1_clock; // @[Math.scala 150:24:@26796.4]
  wire  x325_sum_1_reset; // @[Math.scala 150:24:@26796.4]
  wire [31:0] x325_sum_1_io_a; // @[Math.scala 150:24:@26796.4]
  wire [31:0] x325_sum_1_io_b; // @[Math.scala 150:24:@26796.4]
  wire  x325_sum_1_io_flow; // @[Math.scala 150:24:@26796.4]
  wire [31:0] x325_sum_1_io_result; // @[Math.scala 150:24:@26796.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@26806.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@26806.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@26806.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@26806.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@26806.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@26815.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@26815.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@26815.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@26815.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@26815.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@26824.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@26824.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@26824.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@26824.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@26824.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@26836.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@26836.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@26836.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@26836.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@26836.4]
  wire  x328_rdcol_1_clock; // @[Math.scala 150:24:@26859.4]
  wire  x328_rdcol_1_reset; // @[Math.scala 150:24:@26859.4]
  wire [31:0] x328_rdcol_1_io_a; // @[Math.scala 150:24:@26859.4]
  wire [31:0] x328_rdcol_1_io_b; // @[Math.scala 150:24:@26859.4]
  wire  x328_rdcol_1_io_flow; // @[Math.scala 150:24:@26859.4]
  wire [31:0] x328_rdcol_1_io_result; // @[Math.scala 150:24:@26859.4]
  wire  x334_sum_1_clock; // @[Math.scala 150:24:@26910.4]
  wire  x334_sum_1_reset; // @[Math.scala 150:24:@26910.4]
  wire [31:0] x334_sum_1_io_a; // @[Math.scala 150:24:@26910.4]
  wire [31:0] x334_sum_1_io_b; // @[Math.scala 150:24:@26910.4]
  wire  x334_sum_1_io_flow; // @[Math.scala 150:24:@26910.4]
  wire [31:0] x334_sum_1_io_result; // @[Math.scala 150:24:@26910.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@26920.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@26920.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@26920.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@26920.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@26920.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@26929.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@26929.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@26929.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@26929.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@26929.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@26938.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@26938.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@26938.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@26938.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@26938.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@26950.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@26950.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@26950.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@26950.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@26950.4]
  wire  x337_rdrow_1_clock; // @[Math.scala 191:24:@26973.4]
  wire  x337_rdrow_1_reset; // @[Math.scala 191:24:@26973.4]
  wire [31:0] x337_rdrow_1_io_a; // @[Math.scala 191:24:@26973.4]
  wire [31:0] x337_rdrow_1_io_b; // @[Math.scala 191:24:@26973.4]
  wire  x337_rdrow_1_io_flow; // @[Math.scala 191:24:@26973.4]
  wire [31:0] x337_rdrow_1_io_result; // @[Math.scala 191:24:@26973.4]
  wire  x516_sub_1_clock; // @[Math.scala 191:24:@27045.4]
  wire  x516_sub_1_reset; // @[Math.scala 191:24:@27045.4]
  wire [31:0] x516_sub_1_io_a; // @[Math.scala 191:24:@27045.4]
  wire [31:0] x516_sub_1_io_b; // @[Math.scala 191:24:@27045.4]
  wire  x516_sub_1_io_flow; // @[Math.scala 191:24:@27045.4]
  wire [31:0] x516_sub_1_io_result; // @[Math.scala 191:24:@27045.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@27055.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@27055.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@27055.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@27055.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@27055.4]
  wire  x345_sum_1_clock; // @[Math.scala 150:24:@27064.4]
  wire  x345_sum_1_reset; // @[Math.scala 150:24:@27064.4]
  wire [31:0] x345_sum_1_io_a; // @[Math.scala 150:24:@27064.4]
  wire [31:0] x345_sum_1_io_b; // @[Math.scala 150:24:@27064.4]
  wire  x345_sum_1_io_flow; // @[Math.scala 150:24:@27064.4]
  wire [31:0] x345_sum_1_io_result; // @[Math.scala 150:24:@27064.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@27074.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@27074.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@27074.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@27074.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@27074.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@27083.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@27083.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@27083.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@27083.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@27083.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@27095.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@27095.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@27095.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@27095.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@27095.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@27116.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@27116.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@27116.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@27116.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@27116.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@27131.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@27131.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@27131.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@27131.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@27131.4]
  wire  x350_sum_1_clock; // @[Math.scala 150:24:@27142.4]
  wire  x350_sum_1_reset; // @[Math.scala 150:24:@27142.4]
  wire [31:0] x350_sum_1_io_a; // @[Math.scala 150:24:@27142.4]
  wire [31:0] x350_sum_1_io_b; // @[Math.scala 150:24:@27142.4]
  wire  x350_sum_1_io_flow; // @[Math.scala 150:24:@27142.4]
  wire [31:0] x350_sum_1_io_result; // @[Math.scala 150:24:@27142.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@27152.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@27164.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@27164.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@27164.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@27164.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@27164.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@27191.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@27191.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@27191.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@27191.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@27191.4]
  wire  x355_sum_1_clock; // @[Math.scala 150:24:@27200.4]
  wire  x355_sum_1_reset; // @[Math.scala 150:24:@27200.4]
  wire [31:0] x355_sum_1_io_a; // @[Math.scala 150:24:@27200.4]
  wire [31:0] x355_sum_1_io_b; // @[Math.scala 150:24:@27200.4]
  wire  x355_sum_1_io_flow; // @[Math.scala 150:24:@27200.4]
  wire [31:0] x355_sum_1_io_result; // @[Math.scala 150:24:@27200.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@27210.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@27210.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@27210.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@27210.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@27210.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@27222.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@27222.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@27222.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@27222.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@27222.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@27249.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@27249.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@27249.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@27249.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@27249.4]
  wire  x360_sum_1_clock; // @[Math.scala 150:24:@27258.4]
  wire  x360_sum_1_reset; // @[Math.scala 150:24:@27258.4]
  wire [31:0] x360_sum_1_io_a; // @[Math.scala 150:24:@27258.4]
  wire [31:0] x360_sum_1_io_b; // @[Math.scala 150:24:@27258.4]
  wire  x360_sum_1_io_flow; // @[Math.scala 150:24:@27258.4]
  wire [31:0] x360_sum_1_io_result; // @[Math.scala 150:24:@27258.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@27268.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@27268.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@27268.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@27268.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@27268.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@27280.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@27280.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@27280.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@27280.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@27280.4]
  wire  x363_rdrow_1_clock; // @[Math.scala 191:24:@27303.4]
  wire  x363_rdrow_1_reset; // @[Math.scala 191:24:@27303.4]
  wire [31:0] x363_rdrow_1_io_a; // @[Math.scala 191:24:@27303.4]
  wire [31:0] x363_rdrow_1_io_b; // @[Math.scala 191:24:@27303.4]
  wire  x363_rdrow_1_io_flow; // @[Math.scala 191:24:@27303.4]
  wire [31:0] x363_rdrow_1_io_result; // @[Math.scala 191:24:@27303.4]
  wire  x521_sub_1_clock; // @[Math.scala 191:24:@27375.4]
  wire  x521_sub_1_reset; // @[Math.scala 191:24:@27375.4]
  wire [31:0] x521_sub_1_io_a; // @[Math.scala 191:24:@27375.4]
  wire [31:0] x521_sub_1_io_b; // @[Math.scala 191:24:@27375.4]
  wire  x521_sub_1_io_flow; // @[Math.scala 191:24:@27375.4]
  wire [31:0] x521_sub_1_io_result; // @[Math.scala 191:24:@27375.4]
  wire  x371_sum_1_clock; // @[Math.scala 150:24:@27385.4]
  wire  x371_sum_1_reset; // @[Math.scala 150:24:@27385.4]
  wire [31:0] x371_sum_1_io_a; // @[Math.scala 150:24:@27385.4]
  wire [31:0] x371_sum_1_io_b; // @[Math.scala 150:24:@27385.4]
  wire  x371_sum_1_io_flow; // @[Math.scala 150:24:@27385.4]
  wire [31:0] x371_sum_1_io_result; // @[Math.scala 150:24:@27385.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@27395.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@27395.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@27395.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@27395.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@27395.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@27404.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@27404.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@27404.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@27404.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@27404.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@27416.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@27416.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@27416.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@27416.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@27416.4]
  wire  x376_sum_1_clock; // @[Math.scala 150:24:@27443.4]
  wire  x376_sum_1_reset; // @[Math.scala 150:24:@27443.4]
  wire [31:0] x376_sum_1_io_a; // @[Math.scala 150:24:@27443.4]
  wire [31:0] x376_sum_1_io_b; // @[Math.scala 150:24:@27443.4]
  wire  x376_sum_1_io_flow; // @[Math.scala 150:24:@27443.4]
  wire [31:0] x376_sum_1_io_result; // @[Math.scala 150:24:@27443.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@27453.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@27453.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@27453.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@27453.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@27453.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@27465.4]
  wire  x381_sum_1_clock; // @[Math.scala 150:24:@27492.4]
  wire  x381_sum_1_reset; // @[Math.scala 150:24:@27492.4]
  wire [31:0] x381_sum_1_io_a; // @[Math.scala 150:24:@27492.4]
  wire [31:0] x381_sum_1_io_b; // @[Math.scala 150:24:@27492.4]
  wire  x381_sum_1_io_flow; // @[Math.scala 150:24:@27492.4]
  wire [31:0] x381_sum_1_io_result; // @[Math.scala 150:24:@27492.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@27502.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@27502.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@27502.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@27502.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@27502.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@27514.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@27514.4]
  wire  x386_sum_1_clock; // @[Math.scala 150:24:@27543.4]
  wire  x386_sum_1_reset; // @[Math.scala 150:24:@27543.4]
  wire [31:0] x386_sum_1_io_a; // @[Math.scala 150:24:@27543.4]
  wire [31:0] x386_sum_1_io_b; // @[Math.scala 150:24:@27543.4]
  wire  x386_sum_1_io_flow; // @[Math.scala 150:24:@27543.4]
  wire [31:0] x386_sum_1_io_result; // @[Math.scala 150:24:@27543.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@27553.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@27553.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@27553.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@27553.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@27553.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@27565.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@27588.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@27588.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@27588.4]
  wire [32:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@27588.4]
  wire [32:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@27588.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@27600.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@27600.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@27600.4]
  wire [32:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@27600.4]
  wire [32:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@27600.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@27612.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@27612.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@27612.4]
  wire [33:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@27612.4]
  wire [33:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@27612.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@27624.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@27624.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@27624.4]
  wire [32:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@27624.4]
  wire [32:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@27624.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@27636.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@27636.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@27636.4]
  wire [32:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@27636.4]
  wire [32:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@27636.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@27646.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@27646.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@27646.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@27646.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@27646.4]
  wire  x394_x13_1_clock; // @[Math.scala 150:24:@27655.4]
  wire  x394_x13_1_reset; // @[Math.scala 150:24:@27655.4]
  wire [31:0] x394_x13_1_io_a; // @[Math.scala 150:24:@27655.4]
  wire [31:0] x394_x13_1_io_b; // @[Math.scala 150:24:@27655.4]
  wire  x394_x13_1_io_flow; // @[Math.scala 150:24:@27655.4]
  wire [31:0] x394_x13_1_io_result; // @[Math.scala 150:24:@27655.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@27665.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@27665.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@27665.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@27665.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@27665.4]
  wire  x395_x14_1_clock; // @[Math.scala 150:24:@27674.4]
  wire  x395_x14_1_reset; // @[Math.scala 150:24:@27674.4]
  wire [31:0] x395_x14_1_io_a; // @[Math.scala 150:24:@27674.4]
  wire [31:0] x395_x14_1_io_b; // @[Math.scala 150:24:@27674.4]
  wire  x395_x14_1_io_flow; // @[Math.scala 150:24:@27674.4]
  wire [31:0] x395_x14_1_io_result; // @[Math.scala 150:24:@27674.4]
  wire  x396_x13_1_clock; // @[Math.scala 150:24:@27684.4]
  wire  x396_x13_1_reset; // @[Math.scala 150:24:@27684.4]
  wire [31:0] x396_x13_1_io_a; // @[Math.scala 150:24:@27684.4]
  wire [31:0] x396_x13_1_io_b; // @[Math.scala 150:24:@27684.4]
  wire  x396_x13_1_io_flow; // @[Math.scala 150:24:@27684.4]
  wire [31:0] x396_x13_1_io_result; // @[Math.scala 150:24:@27684.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@27694.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@27694.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@27694.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@27694.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@27694.4]
  wire  x397_x14_1_clock; // @[Math.scala 150:24:@27703.4]
  wire  x397_x14_1_reset; // @[Math.scala 150:24:@27703.4]
  wire [31:0] x397_x14_1_io_a; // @[Math.scala 150:24:@27703.4]
  wire [31:0] x397_x14_1_io_b; // @[Math.scala 150:24:@27703.4]
  wire  x397_x14_1_io_flow; // @[Math.scala 150:24:@27703.4]
  wire [31:0] x397_x14_1_io_result; // @[Math.scala 150:24:@27703.4]
  wire  x398_x13_1_clock; // @[Math.scala 150:24:@27713.4]
  wire  x398_x13_1_reset; // @[Math.scala 150:24:@27713.4]
  wire [31:0] x398_x13_1_io_a; // @[Math.scala 150:24:@27713.4]
  wire [31:0] x398_x13_1_io_b; // @[Math.scala 150:24:@27713.4]
  wire  x398_x13_1_io_flow; // @[Math.scala 150:24:@27713.4]
  wire [31:0] x398_x13_1_io_result; // @[Math.scala 150:24:@27713.4]
  wire  x399_x14_1_clock; // @[Math.scala 150:24:@27723.4]
  wire  x399_x14_1_reset; // @[Math.scala 150:24:@27723.4]
  wire [31:0] x399_x14_1_io_a; // @[Math.scala 150:24:@27723.4]
  wire [31:0] x399_x14_1_io_b; // @[Math.scala 150:24:@27723.4]
  wire  x399_x14_1_io_flow; // @[Math.scala 150:24:@27723.4]
  wire [31:0] x399_x14_1_io_result; // @[Math.scala 150:24:@27723.4]
  wire  x400_x13_1_clock; // @[Math.scala 150:24:@27733.4]
  wire  x400_x13_1_reset; // @[Math.scala 150:24:@27733.4]
  wire [31:0] x400_x13_1_io_a; // @[Math.scala 150:24:@27733.4]
  wire [31:0] x400_x13_1_io_b; // @[Math.scala 150:24:@27733.4]
  wire  x400_x13_1_io_flow; // @[Math.scala 150:24:@27733.4]
  wire [31:0] x400_x13_1_io_result; // @[Math.scala 150:24:@27733.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@27743.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@27743.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@27743.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@27743.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@27743.4]
  wire  x401_sum_1_clock; // @[Math.scala 150:24:@27752.4]
  wire  x401_sum_1_reset; // @[Math.scala 150:24:@27752.4]
  wire [31:0] x401_sum_1_io_a; // @[Math.scala 150:24:@27752.4]
  wire [31:0] x401_sum_1_io_b; // @[Math.scala 150:24:@27752.4]
  wire  x401_sum_1_io_flow; // @[Math.scala 150:24:@27752.4]
  wire [31:0] x401_sum_1_io_result; // @[Math.scala 150:24:@27752.4]
  wire [31:0] x402_1_io_b; // @[Math.scala 720:24:@27762.4]
  wire [31:0] x402_1_io_result; // @[Math.scala 720:24:@27762.4]
  wire  x403_mul_1_clock; // @[Math.scala 262:24:@27773.4]
  wire [31:0] x403_mul_1_io_a; // @[Math.scala 262:24:@27773.4]
  wire [31:0] x403_mul_1_io_b; // @[Math.scala 262:24:@27773.4]
  wire  x403_mul_1_io_flow; // @[Math.scala 262:24:@27773.4]
  wire [31:0] x403_mul_1_io_result; // @[Math.scala 262:24:@27773.4]
  wire [31:0] x404_1_io_b; // @[Math.scala 720:24:@27783.4]
  wire [31:0] x404_1_io_result; // @[Math.scala 720:24:@27783.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@27792.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@27792.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@27792.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@27792.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@27792.4]
  wire  x405_sub_1_clock; // @[Math.scala 191:24:@27801.4]
  wire  x405_sub_1_reset; // @[Math.scala 191:24:@27801.4]
  wire [31:0] x405_sub_1_io_a; // @[Math.scala 191:24:@27801.4]
  wire [31:0] x405_sub_1_io_b; // @[Math.scala 191:24:@27801.4]
  wire  x405_sub_1_io_flow; // @[Math.scala 191:24:@27801.4]
  wire [31:0] x405_sub_1_io_result; // @[Math.scala 191:24:@27801.4]
  wire  x407_sub_1_clock; // @[Math.scala 191:24:@27816.4]
  wire  x407_sub_1_reset; // @[Math.scala 191:24:@27816.4]
  wire [31:0] x407_sub_1_io_a; // @[Math.scala 191:24:@27816.4]
  wire [31:0] x407_sub_1_io_b; // @[Math.scala 191:24:@27816.4]
  wire  x407_sub_1_io_flow; // @[Math.scala 191:24:@27816.4]
  wire [31:0] x407_sub_1_io_result; // @[Math.scala 191:24:@27816.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@27839.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@27839.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@27839.4]
  wire [31:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@27839.4]
  wire [31:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@27839.4]
  wire [31:0] x411_1_io_b; // @[Math.scala 720:24:@27848.4]
  wire [31:0] x411_1_io_result; // @[Math.scala 720:24:@27848.4]
  wire  x412_mul_1_clock; // @[Math.scala 262:24:@27859.4]
  wire [31:0] x412_mul_1_io_a; // @[Math.scala 262:24:@27859.4]
  wire [31:0] x412_mul_1_io_b; // @[Math.scala 262:24:@27859.4]
  wire  x412_mul_1_io_flow; // @[Math.scala 262:24:@27859.4]
  wire [31:0] x412_mul_1_io_result; // @[Math.scala 262:24:@27859.4]
  wire [31:0] x413_1_io_b; // @[Math.scala 720:24:@27869.4]
  wire [31:0] x413_1_io_result; // @[Math.scala 720:24:@27869.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@27878.4]
  wire [31:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@27878.4]
  wire [31:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@27878.4]
  wire  x414_sum_1_clock; // @[Math.scala 150:24:@27887.4]
  wire  x414_sum_1_reset; // @[Math.scala 150:24:@27887.4]
  wire [31:0] x414_sum_1_io_a; // @[Math.scala 150:24:@27887.4]
  wire [31:0] x414_sum_1_io_b; // @[Math.scala 150:24:@27887.4]
  wire  x414_sum_1_io_flow; // @[Math.scala 150:24:@27887.4]
  wire [31:0] x414_sum_1_io_result; // @[Math.scala 150:24:@27887.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@27899.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@27899.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@27899.4]
  wire [32:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@27899.4]
  wire [32:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@27899.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@27911.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@27911.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@27911.4]
  wire [32:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@27911.4]
  wire [32:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@27911.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@27923.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@27923.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@27923.4]
  wire [33:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@27923.4]
  wire [33:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@27923.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@27935.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@27935.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@27935.4]
  wire [32:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@27935.4]
  wire [32:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@27935.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@27947.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@27947.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@27947.4]
  wire [32:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@27947.4]
  wire [32:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@27947.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@27957.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@27957.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@27957.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@27957.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@27957.4]
  wire  x420_x13_1_clock; // @[Math.scala 150:24:@27966.4]
  wire  x420_x13_1_reset; // @[Math.scala 150:24:@27966.4]
  wire [31:0] x420_x13_1_io_a; // @[Math.scala 150:24:@27966.4]
  wire [31:0] x420_x13_1_io_b; // @[Math.scala 150:24:@27966.4]
  wire  x420_x13_1_io_flow; // @[Math.scala 150:24:@27966.4]
  wire [31:0] x420_x13_1_io_result; // @[Math.scala 150:24:@27966.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@27976.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@27976.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@27976.4]
  wire [31:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@27976.4]
  wire [31:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@27976.4]
  wire  x421_x14_1_clock; // @[Math.scala 150:24:@27985.4]
  wire  x421_x14_1_reset; // @[Math.scala 150:24:@27985.4]
  wire [31:0] x421_x14_1_io_a; // @[Math.scala 150:24:@27985.4]
  wire [31:0] x421_x14_1_io_b; // @[Math.scala 150:24:@27985.4]
  wire  x421_x14_1_io_flow; // @[Math.scala 150:24:@27985.4]
  wire [31:0] x421_x14_1_io_result; // @[Math.scala 150:24:@27985.4]
  wire  x422_x13_1_clock; // @[Math.scala 150:24:@27995.4]
  wire  x422_x13_1_reset; // @[Math.scala 150:24:@27995.4]
  wire [31:0] x422_x13_1_io_a; // @[Math.scala 150:24:@27995.4]
  wire [31:0] x422_x13_1_io_b; // @[Math.scala 150:24:@27995.4]
  wire  x422_x13_1_io_flow; // @[Math.scala 150:24:@27995.4]
  wire [31:0] x422_x13_1_io_result; // @[Math.scala 150:24:@27995.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@28005.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@28005.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@28005.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@28005.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@28005.4]
  wire  x423_x14_1_clock; // @[Math.scala 150:24:@28016.4]
  wire  x423_x14_1_reset; // @[Math.scala 150:24:@28016.4]
  wire [31:0] x423_x14_1_io_a; // @[Math.scala 150:24:@28016.4]
  wire [31:0] x423_x14_1_io_b; // @[Math.scala 150:24:@28016.4]
  wire  x423_x14_1_io_flow; // @[Math.scala 150:24:@28016.4]
  wire [31:0] x423_x14_1_io_result; // @[Math.scala 150:24:@28016.4]
  wire  x424_x13_1_clock; // @[Math.scala 150:24:@28026.4]
  wire  x424_x13_1_reset; // @[Math.scala 150:24:@28026.4]
  wire [31:0] x424_x13_1_io_a; // @[Math.scala 150:24:@28026.4]
  wire [31:0] x424_x13_1_io_b; // @[Math.scala 150:24:@28026.4]
  wire  x424_x13_1_io_flow; // @[Math.scala 150:24:@28026.4]
  wire [31:0] x424_x13_1_io_result; // @[Math.scala 150:24:@28026.4]
  wire  x425_x14_1_clock; // @[Math.scala 150:24:@28036.4]
  wire  x425_x14_1_reset; // @[Math.scala 150:24:@28036.4]
  wire [31:0] x425_x14_1_io_a; // @[Math.scala 150:24:@28036.4]
  wire [31:0] x425_x14_1_io_b; // @[Math.scala 150:24:@28036.4]
  wire  x425_x14_1_io_flow; // @[Math.scala 150:24:@28036.4]
  wire [31:0] x425_x14_1_io_result; // @[Math.scala 150:24:@28036.4]
  wire  x426_x13_1_clock; // @[Math.scala 150:24:@28046.4]
  wire  x426_x13_1_reset; // @[Math.scala 150:24:@28046.4]
  wire [31:0] x426_x13_1_io_a; // @[Math.scala 150:24:@28046.4]
  wire [31:0] x426_x13_1_io_b; // @[Math.scala 150:24:@28046.4]
  wire  x426_x13_1_io_flow; // @[Math.scala 150:24:@28046.4]
  wire [31:0] x426_x13_1_io_result; // @[Math.scala 150:24:@28046.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@28056.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@28056.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@28056.4]
  wire [31:0] RetimeWrapper_80_io_in; // @[package.scala 93:22:@28056.4]
  wire [31:0] RetimeWrapper_80_io_out; // @[package.scala 93:22:@28056.4]
  wire  x427_sum_1_clock; // @[Math.scala 150:24:@28065.4]
  wire  x427_sum_1_reset; // @[Math.scala 150:24:@28065.4]
  wire [31:0] x427_sum_1_io_a; // @[Math.scala 150:24:@28065.4]
  wire [31:0] x427_sum_1_io_b; // @[Math.scala 150:24:@28065.4]
  wire  x427_sum_1_io_flow; // @[Math.scala 150:24:@28065.4]
  wire [31:0] x427_sum_1_io_result; // @[Math.scala 150:24:@28065.4]
  wire [31:0] x428_1_io_b; // @[Math.scala 720:24:@28075.4]
  wire [31:0] x428_1_io_result; // @[Math.scala 720:24:@28075.4]
  wire  x429_mul_1_clock; // @[Math.scala 262:24:@28086.4]
  wire [31:0] x429_mul_1_io_a; // @[Math.scala 262:24:@28086.4]
  wire [31:0] x429_mul_1_io_b; // @[Math.scala 262:24:@28086.4]
  wire  x429_mul_1_io_flow; // @[Math.scala 262:24:@28086.4]
  wire [31:0] x429_mul_1_io_result; // @[Math.scala 262:24:@28086.4]
  wire [31:0] x430_1_io_b; // @[Math.scala 720:24:@28096.4]
  wire [31:0] x430_1_io_result; // @[Math.scala 720:24:@28096.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@28105.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@28105.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@28105.4]
  wire [31:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@28105.4]
  wire [31:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@28105.4]
  wire  x431_sub_1_clock; // @[Math.scala 191:24:@28114.4]
  wire  x431_sub_1_reset; // @[Math.scala 191:24:@28114.4]
  wire [31:0] x431_sub_1_io_a; // @[Math.scala 191:24:@28114.4]
  wire [31:0] x431_sub_1_io_b; // @[Math.scala 191:24:@28114.4]
  wire  x431_sub_1_io_flow; // @[Math.scala 191:24:@28114.4]
  wire [31:0] x431_sub_1_io_result; // @[Math.scala 191:24:@28114.4]
  wire  x433_sub_1_clock; // @[Math.scala 191:24:@28129.4]
  wire  x433_sub_1_reset; // @[Math.scala 191:24:@28129.4]
  wire [31:0] x433_sub_1_io_a; // @[Math.scala 191:24:@28129.4]
  wire [31:0] x433_sub_1_io_b; // @[Math.scala 191:24:@28129.4]
  wire  x433_sub_1_io_flow; // @[Math.scala 191:24:@28129.4]
  wire [31:0] x433_sub_1_io_result; // @[Math.scala 191:24:@28129.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@28152.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@28152.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@28152.4]
  wire [31:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@28152.4]
  wire [31:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@28152.4]
  wire [31:0] x437_1_io_b; // @[Math.scala 720:24:@28161.4]
  wire [31:0] x437_1_io_result; // @[Math.scala 720:24:@28161.4]
  wire  x438_mul_1_clock; // @[Math.scala 262:24:@28172.4]
  wire [31:0] x438_mul_1_io_a; // @[Math.scala 262:24:@28172.4]
  wire [31:0] x438_mul_1_io_b; // @[Math.scala 262:24:@28172.4]
  wire  x438_mul_1_io_flow; // @[Math.scala 262:24:@28172.4]
  wire [31:0] x438_mul_1_io_result; // @[Math.scala 262:24:@28172.4]
  wire [31:0] x439_1_io_b; // @[Math.scala 720:24:@28182.4]
  wire [31:0] x439_1_io_result; // @[Math.scala 720:24:@28182.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@28191.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@28191.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@28191.4]
  wire [31:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@28191.4]
  wire [31:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@28191.4]
  wire  x440_sum_1_clock; // @[Math.scala 150:24:@28200.4]
  wire  x440_sum_1_reset; // @[Math.scala 150:24:@28200.4]
  wire [31:0] x440_sum_1_io_a; // @[Math.scala 150:24:@28200.4]
  wire [31:0] x440_sum_1_io_b; // @[Math.scala 150:24:@28200.4]
  wire  x440_sum_1_io_flow; // @[Math.scala 150:24:@28200.4]
  wire [31:0] x440_sum_1_io_result; // @[Math.scala 150:24:@28200.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@28216.4]
  wire [63:0] RetimeWrapper_84_io_in; // @[package.scala 93:22:@28216.4]
  wire [63:0] RetimeWrapper_84_io_out; // @[package.scala 93:22:@28216.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@28225.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@28225.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@28225.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@28225.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@28225.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@28234.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@28234.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@28234.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@28234.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@28234.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@28243.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@28243.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@28243.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@28243.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@28243.4]
  wire  b286; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 62:18:@26121.4]
  wire  b287; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 63:18:@26122.4]
  wire  _T_205; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 67:30:@26124.4]
  wire  _T_206; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 67:37:@26125.4]
  wire  _T_210; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:76:@26130.4]
  wire  _T_211; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:62:@26131.4]
  wire  _T_213; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:101:@26132.4]
  wire [63:0] x527_x288_D1_0_number; // @[package.scala 96:25:@26141.4 package.scala 96:25:@26142.4]
  wire [31:0] b284_number; // @[Math.scala 723:22:@26106.4 Math.scala 724:14:@26107.4]
  wire [31:0] _T_243; // @[Math.scala 406:49:@26250.4]
  wire [31:0] _T_245; // @[Math.scala 406:56:@26252.4]
  wire [31:0] _T_246; // @[Math.scala 406:56:@26253.4]
  wire [31:0] x503_number; // @[implicits.scala 133:21:@26254.4]
  wire [31:0] _T_256; // @[Math.scala 406:49:@26263.4]
  wire [31:0] _T_258; // @[Math.scala 406:56:@26265.4]
  wire [31:0] _T_259; // @[Math.scala 406:56:@26266.4]
  wire [31:0] b285_number; // @[Math.scala 723:22:@26118.4 Math.scala 724:14:@26119.4]
  wire [31:0] _T_268; // @[Math.scala 406:49:@26274.4]
  wire [31:0] _T_270; // @[Math.scala 406:56:@26276.4]
  wire [31:0] _T_271; // @[Math.scala 406:56:@26277.4]
  wire  _T_275; // @[FixedPoint.scala 50:25:@26283.4]
  wire [1:0] _T_279; // @[Bitwise.scala 72:12:@26285.4]
  wire [29:0] _T_280; // @[FixedPoint.scala 18:52:@26286.4]
  wire  _T_286; // @[Math.scala 451:55:@26288.4]
  wire [1:0] _T_287; // @[FixedPoint.scala 18:52:@26289.4]
  wire  _T_293; // @[Math.scala 451:110:@26291.4]
  wire  _T_294; // @[Math.scala 451:94:@26292.4]
  wire [31:0] _T_296; // @[Cat.scala 30:58:@26294.4]
  wire [31:0] x296_1_number; // @[Math.scala 454:20:@26295.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@26300.4]
  wire [40:0] _T_301; // @[Math.scala 461:32:@26300.4]
  wire [36:0] _GEN_1; // @[Math.scala 461:32:@26305.4]
  wire [36:0] _T_304; // @[Math.scala 461:32:@26305.4]
  wire  _T_310; // @[FixedPoint.scala 50:25:@26320.4]
  wire [1:0] _T_314; // @[Bitwise.scala 72:12:@26322.4]
  wire [29:0] _T_315; // @[FixedPoint.scala 18:52:@26323.4]
  wire  _T_321; // @[Math.scala 451:55:@26325.4]
  wire [1:0] _T_322; // @[FixedPoint.scala 18:52:@26326.4]
  wire  _T_328; // @[Math.scala 451:110:@26328.4]
  wire  _T_329; // @[Math.scala 451:94:@26329.4]
  wire [31:0] _T_331; // @[Cat.scala 30:58:@26331.4]
  wire  _T_359; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:101:@26408.4]
  wire  _T_363; // @[package.scala 96:25:@26416.4 package.scala 96:25:@26417.4]
  wire  _T_365; // @[implicits.scala 55:10:@26418.4]
  wire  _T_366; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:118:@26419.4]
  wire  _T_368; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:206:@26421.4]
  wire  _T_369; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:225:@26422.4]
  wire  x531_b286_D3; // @[package.scala 96:25:@26378.4 package.scala 96:25:@26379.4]
  wire  _T_370; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:251:@26423.4]
  wire  x534_b287_D3; // @[package.scala 96:25:@26405.4 package.scala 96:25:@26406.4]
  wire [31:0] x301_rdcol_number; // @[Math.scala 154:22:@26440.4 Math.scala 155:14:@26441.4]
  wire [31:0] _T_387; // @[Math.scala 406:49:@26449.4]
  wire [31:0] _T_389; // @[Math.scala 406:56:@26451.4]
  wire [31:0] _T_390; // @[Math.scala 406:56:@26452.4]
  wire  _T_394; // @[FixedPoint.scala 50:25:@26458.4]
  wire [1:0] _T_398; // @[Bitwise.scala 72:12:@26460.4]
  wire [29:0] _T_399; // @[FixedPoint.scala 18:52:@26461.4]
  wire  _T_405; // @[Math.scala 451:55:@26463.4]
  wire [1:0] _T_406; // @[FixedPoint.scala 18:52:@26464.4]
  wire  _T_412; // @[Math.scala 451:110:@26466.4]
  wire  _T_413; // @[Math.scala 451:94:@26467.4]
  wire [31:0] _T_415; // @[Cat.scala 30:58:@26469.4]
  wire  _T_435; // @[package.scala 96:25:@26518.4 package.scala 96:25:@26519.4]
  wire  _T_437; // @[implicits.scala 55:10:@26520.4]
  wire  _T_438; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:118:@26521.4]
  wire  _T_440; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:206:@26523.4]
  wire  _T_441; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:225:@26524.4]
  wire  _T_442; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:251:@26525.4]
  wire [31:0] x538_b284_D6_number; // @[package.scala 96:25:@26539.4 package.scala 96:25:@26540.4]
  wire [31:0] _T_452; // @[Math.scala 476:37:@26545.4]
  wire  x308; // @[Math.scala 476:44:@26547.4]
  wire [31:0] x539_x301_rdcol_D6_number; // @[package.scala 96:25:@26555.4 package.scala 96:25:@26556.4]
  wire [31:0] _T_463; // @[Math.scala 476:37:@26561.4]
  wire  x309; // @[Math.scala 476:44:@26563.4]
  wire  x540_x308_D1; // @[package.scala 96:25:@26571.4 package.scala 96:25:@26572.4]
  wire  x310; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 151:24:@26575.4]
  wire  _T_502; // @[package.scala 96:25:@26643.4 package.scala 96:25:@26644.4]
  wire  _T_504; // @[implicits.scala 55:10:@26645.4]
  wire  _T_505; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 170:146:@26646.4]
  wire  x542_x311_D2; // @[package.scala 96:25:@26595.4 package.scala 96:25:@26596.4]
  wire  _T_506; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 170:234:@26647.4]
  wire  x543_b286_D9; // @[package.scala 96:25:@26604.4 package.scala 96:25:@26605.4]
  wire  _T_507; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 170:242:@26648.4]
  wire  x545_b287_D9; // @[package.scala 96:25:@26622.4 package.scala 96:25:@26623.4]
  wire [31:0] x547_b285_D6_number; // @[package.scala 96:25:@26664.4 package.scala 96:25:@26665.4]
  wire [31:0] _T_520; // @[Math.scala 476:37:@26672.4]
  wire  x314; // @[Math.scala 476:44:@26674.4]
  wire  x315; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 186:59:@26677.4]
  wire  _T_547; // @[package.scala 96:25:@26718.4 package.scala 96:25:@26719.4]
  wire  _T_549; // @[implicits.scala 55:10:@26720.4]
  wire  _T_550; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:194:@26721.4]
  wire  x548_x316_D3; // @[package.scala 96:25:@26688.4 package.scala 96:25:@26689.4]
  wire  _T_551; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:282:@26722.4]
  wire  _T_552; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:290:@26723.4]
  wire [31:0] x319_rdcol_number; // @[Math.scala 154:22:@26742.4 Math.scala 155:14:@26743.4]
  wire [31:0] _T_567; // @[Math.scala 476:37:@26748.4]
  wire  x320; // @[Math.scala 476:44:@26750.4]
  wire  x321; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 207:59:@26753.4]
  wire [31:0] _T_583; // @[Math.scala 406:56:@26764.4]
  wire [31:0] _T_584; // @[Math.scala 406:56:@26765.4]
  wire  _T_588; // @[FixedPoint.scala 50:25:@26771.4]
  wire [1:0] _T_592; // @[Bitwise.scala 72:12:@26773.4]
  wire [29:0] _T_593; // @[FixedPoint.scala 18:52:@26774.4]
  wire  _T_599; // @[Math.scala 451:55:@26776.4]
  wire [1:0] _T_600; // @[FixedPoint.scala 18:52:@26777.4]
  wire  _T_606; // @[Math.scala 451:110:@26779.4]
  wire  _T_607; // @[Math.scala 451:94:@26780.4]
  wire [31:0] _T_609; // @[Cat.scala 30:58:@26782.4]
  wire  _T_638; // @[package.scala 96:25:@26841.4 package.scala 96:25:@26842.4]
  wire  _T_640; // @[implicits.scala 55:10:@26843.4]
  wire  _T_641; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:194:@26844.4]
  wire  x554_x322_D2; // @[package.scala 96:25:@26829.4 package.scala 96:25:@26830.4]
  wire  _T_642; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:282:@26845.4]
  wire  _T_643; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:290:@26846.4]
  wire [31:0] x328_rdcol_number; // @[Math.scala 154:22:@26865.4 Math.scala 155:14:@26866.4]
  wire [31:0] _T_658; // @[Math.scala 476:37:@26871.4]
  wire  x329; // @[Math.scala 476:44:@26873.4]
  wire  x330; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 236:59:@26876.4]
  wire [31:0] _T_674; // @[Math.scala 406:56:@26887.4]
  wire [31:0] _T_675; // @[Math.scala 406:56:@26888.4]
  wire  _T_679; // @[FixedPoint.scala 50:25:@26894.4]
  wire [1:0] _T_683; // @[Bitwise.scala 72:12:@26896.4]
  wire [29:0] _T_684; // @[FixedPoint.scala 18:52:@26897.4]
  wire  _T_690; // @[Math.scala 451:55:@26899.4]
  wire [1:0] _T_691; // @[FixedPoint.scala 18:52:@26900.4]
  wire  _T_697; // @[Math.scala 451:110:@26902.4]
  wire  _T_698; // @[Math.scala 451:94:@26903.4]
  wire [31:0] _T_700; // @[Cat.scala 30:58:@26905.4]
  wire  _T_726; // @[package.scala 96:25:@26955.4 package.scala 96:25:@26956.4]
  wire  _T_728; // @[implicits.scala 55:10:@26957.4]
  wire  _T_729; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 255:194:@26958.4]
  wire  x557_x331_D2; // @[package.scala 96:25:@26943.4 package.scala 96:25:@26944.4]
  wire  _T_730; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 255:282:@26959.4]
  wire  _T_731; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 255:290:@26960.4]
  wire [31:0] x337_rdrow_number; // @[Math.scala 195:22:@26979.4 Math.scala 196:14:@26980.4]
  wire [31:0] _T_748; // @[Math.scala 406:49:@26986.4]
  wire [31:0] _T_750; // @[Math.scala 406:56:@26988.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@26989.4]
  wire [31:0] x512_number; // @[implicits.scala 133:21:@26990.4]
  wire  x339; // @[Math.scala 476:44:@26998.4]
  wire  x340; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 265:24:@27001.4]
  wire [31:0] _T_772; // @[Math.scala 406:49:@27010.4]
  wire [31:0] _T_774; // @[Math.scala 406:56:@27012.4]
  wire [31:0] _T_775; // @[Math.scala 406:56:@27013.4]
  wire  _T_779; // @[FixedPoint.scala 50:25:@27019.4]
  wire [1:0] _T_783; // @[Bitwise.scala 72:12:@27021.4]
  wire [29:0] _T_784; // @[FixedPoint.scala 18:52:@27022.4]
  wire  _T_790; // @[Math.scala 451:55:@27024.4]
  wire [1:0] _T_791; // @[FixedPoint.scala 18:52:@27025.4]
  wire  _T_797; // @[Math.scala 451:110:@27027.4]
  wire  _T_798; // @[Math.scala 451:94:@27028.4]
  wire [31:0] _T_800; // @[Cat.scala 30:58:@27030.4]
  wire [31:0] x343_1_number; // @[Math.scala 454:20:@27031.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@27036.4]
  wire [40:0] _T_805; // @[Math.scala 461:32:@27036.4]
  wire [36:0] _GEN_3; // @[Math.scala 461:32:@27041.4]
  wire [36:0] _T_808; // @[Math.scala 461:32:@27041.4]
  wire  _T_835; // @[package.scala 96:25:@27100.4 package.scala 96:25:@27101.4]
  wire  _T_837; // @[implicits.scala 55:10:@27102.4]
  wire  _T_838; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:194:@27103.4]
  wire  x560_x341_D2; // @[package.scala 96:25:@27088.4 package.scala 96:25:@27089.4]
  wire  _T_839; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:282:@27104.4]
  wire  _T_840; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:290:@27105.4]
  wire  x561_x314_D1; // @[package.scala 96:25:@27121.4 package.scala 96:25:@27122.4]
  wire  x348; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 302:59:@27125.4]
  wire  _T_872; // @[package.scala 96:25:@27169.4 package.scala 96:25:@27170.4]
  wire  _T_874; // @[implicits.scala 55:10:@27171.4]
  wire  _T_875; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:194:@27172.4]
  wire  x563_x349_D2; // @[package.scala 96:25:@27157.4 package.scala 96:25:@27158.4]
  wire  _T_876; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:282:@27173.4]
  wire  _T_877; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:290:@27174.4]
  wire  x353; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 321:59:@27185.4]
  wire  _T_904; // @[package.scala 96:25:@27227.4 package.scala 96:25:@27228.4]
  wire  _T_906; // @[implicits.scala 55:10:@27229.4]
  wire  _T_907; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:194:@27230.4]
  wire  x565_x354_D2; // @[package.scala 96:25:@27215.4 package.scala 96:25:@27216.4]
  wire  _T_908; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:282:@27231.4]
  wire  _T_909; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:290:@27232.4]
  wire  x358; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 338:59:@27243.4]
  wire  _T_936; // @[package.scala 96:25:@27285.4 package.scala 96:25:@27286.4]
  wire  _T_938; // @[implicits.scala 55:10:@27287.4]
  wire  _T_939; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:194:@27288.4]
  wire  x567_x359_D2; // @[package.scala 96:25:@27273.4 package.scala 96:25:@27274.4]
  wire  _T_940; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:282:@27289.4]
  wire  _T_941; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:290:@27290.4]
  wire [31:0] x363_rdrow_number; // @[Math.scala 195:22:@27309.4 Math.scala 196:14:@27310.4]
  wire [31:0] _T_958; // @[Math.scala 406:49:@27316.4]
  wire [31:0] _T_960; // @[Math.scala 406:56:@27318.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@27319.4]
  wire [31:0] x517_number; // @[implicits.scala 133:21:@27320.4]
  wire  x365; // @[Math.scala 476:44:@27328.4]
  wire  x366; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 361:24:@27331.4]
  wire [31:0] _T_982; // @[Math.scala 406:49:@27340.4]
  wire [31:0] _T_984; // @[Math.scala 406:56:@27342.4]
  wire [31:0] _T_985; // @[Math.scala 406:56:@27343.4]
  wire  _T_989; // @[FixedPoint.scala 50:25:@27349.4]
  wire [1:0] _T_993; // @[Bitwise.scala 72:12:@27351.4]
  wire [29:0] _T_994; // @[FixedPoint.scala 18:52:@27352.4]
  wire  _T_1000; // @[Math.scala 451:55:@27354.4]
  wire [1:0] _T_1001; // @[FixedPoint.scala 18:52:@27355.4]
  wire  _T_1007; // @[Math.scala 451:110:@27357.4]
  wire  _T_1008; // @[Math.scala 451:94:@27358.4]
  wire [31:0] _T_1010; // @[Cat.scala 30:58:@27360.4]
  wire [31:0] x369_1_number; // @[Math.scala 454:20:@27361.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@27366.4]
  wire [40:0] _T_1015; // @[Math.scala 461:32:@27366.4]
  wire [36:0] _GEN_5; // @[Math.scala 461:32:@27371.4]
  wire [36:0] _T_1018; // @[Math.scala 461:32:@27371.4]
  wire  _T_1042; // @[package.scala 96:25:@27421.4 package.scala 96:25:@27422.4]
  wire  _T_1044; // @[implicits.scala 55:10:@27423.4]
  wire  _T_1045; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 384:194:@27424.4]
  wire  x569_x367_D2; // @[package.scala 96:25:@27409.4 package.scala 96:25:@27410.4]
  wire  _T_1046; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 384:282:@27425.4]
  wire  _T_1047; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 384:290:@27426.4]
  wire  x374; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 388:24:@27437.4]
  wire  _T_1071; // @[package.scala 96:25:@27470.4 package.scala 96:25:@27471.4]
  wire  _T_1073; // @[implicits.scala 55:10:@27472.4]
  wire  _T_1074; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:194:@27473.4]
  wire  x570_x375_D2; // @[package.scala 96:25:@27458.4 package.scala 96:25:@27459.4]
  wire  _T_1075; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:282:@27474.4]
  wire  _T_1076; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:290:@27475.4]
  wire  x379; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 403:24:@27486.4]
  wire  _T_1100; // @[package.scala 96:25:@27519.4 package.scala 96:25:@27520.4]
  wire  _T_1102; // @[implicits.scala 55:10:@27521.4]
  wire  _T_1103; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:194:@27522.4]
  wire  x571_x380_D2; // @[package.scala 96:25:@27507.4 package.scala 96:25:@27508.4]
  wire  _T_1104; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:282:@27523.4]
  wire  _T_1105; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:290:@27524.4]
  wire  x384; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 424:59:@27535.4]
  wire  _T_1131; // @[package.scala 96:25:@27570.4 package.scala 96:25:@27571.4]
  wire  _T_1133; // @[implicits.scala 55:10:@27572.4]
  wire  _T_1134; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 437:194:@27573.4]
  wire  x572_x385_D2; // @[package.scala 96:25:@27558.4 package.scala 96:25:@27559.4]
  wire  _T_1135; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 437:282:@27574.4]
  wire  _T_1136; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 437:290:@27575.4]
  wire [31:0] x317_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 195:29:@26709.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:407:@26730.4]
  wire [32:0] _GEN_6; // @[Math.scala 461:32:@27587.4]
  wire [31:0] x346_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 286:29:@27091.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:407:@27112.4]
  wire [32:0] _GEN_7; // @[Math.scala 461:32:@27599.4]
  wire [31:0] x351_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 313:29:@27160.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:407:@27181.4]
  wire [33:0] _GEN_8; // @[Math.scala 461:32:@27611.4]
  wire [31:0] x356_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 330:29:@27218.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:407:@27239.4]
  wire [32:0] _GEN_9; // @[Math.scala 461:32:@27623.4]
  wire [31:0] x377_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 395:29:@27461.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:407:@27482.4]
  wire [32:0] _GEN_10; // @[Math.scala 461:32:@27635.4]
  wire [31:0] x405_sub_number; // @[Math.scala 195:22:@27807.4 Math.scala 196:14:@27808.4]
  wire  x406; // @[Math.scala 477:37:@27813.4]
  wire [31:0] x407_sub_number; // @[Math.scala 195:22:@27822.4 Math.scala 196:14:@27823.4]
  wire  x408; // @[Math.scala 477:37:@27828.4]
  wire  x409; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 491:24:@27831.4]
  wire [31:0] x326_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 224:29:@26832.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:407:@26853.4]
  wire [32:0] _GEN_11; // @[Math.scala 461:32:@27898.4]
  wire [32:0] _GEN_12; // @[Math.scala 461:32:@27910.4]
  wire [33:0] _GEN_13; // @[Math.scala 461:32:@27922.4]
  wire [31:0] x361_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 347:29:@27276.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:407:@27297.4]
  wire [32:0] _GEN_14; // @[Math.scala 461:32:@27934.4]
  wire [31:0] x382_rd_0_number; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 410:29:@27510.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:407:@27531.4]
  wire [32:0] _GEN_15; // @[Math.scala 461:32:@27946.4]
  wire [31:0] x431_sub_number; // @[Math.scala 195:22:@28120.4 Math.scala 196:14:@28121.4]
  wire  x432; // @[Math.scala 477:37:@28126.4]
  wire [31:0] x433_sub_number; // @[Math.scala 195:22:@28135.4 Math.scala 196:14:@28136.4]
  wire  x434; // @[Math.scala 477:37:@28141.4]
  wire  x435; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 565:24:@28144.4]
  wire [31:0] x414_sum_number; // @[Math.scala 154:22:@27893.4 Math.scala 155:14:@27894.4]
  wire [31:0] x440_sum_number; // @[Math.scala 154:22:@28206.4 Math.scala 155:14:@28207.4]
  wire  _T_1412; // @[package.scala 96:25:@28248.4 package.scala 96:25:@28249.4]
  wire  _T_1414; // @[implicits.scala 55:10:@28250.4]
  wire  x588_b286_D34; // @[package.scala 96:25:@28239.4 package.scala 96:25:@28240.4]
  wire  _T_1415; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 589:117:@28251.4]
  wire  x587_b287_D34; // @[package.scala 96:25:@28230.4 package.scala 96:25:@28231.4]
  wire  _T_1416; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 589:123:@28252.4]
  wire [31:0] x529_x504_D3_number; // @[package.scala 96:25:@26360.4 package.scala 96:25:@26361.4]
  wire [31:0] x532_x299_sum_D1_number; // @[package.scala 96:25:@26387.4 package.scala 96:25:@26388.4]
  wire [31:0] x533_x505_D3_number; // @[package.scala 96:25:@26396.4 package.scala 96:25:@26397.4]
  wire [31:0] x536_x509_D2_number; // @[package.scala 96:25:@26498.4 package.scala 96:25:@26499.4]
  wire [31:0] x537_x305_sum_D1_number; // @[package.scala 96:25:@26507.4 package.scala 96:25:@26508.4]
  wire [31:0] x541_x504_D9_number; // @[package.scala 96:25:@26586.4 package.scala 96:25:@26587.4]
  wire [31:0] x544_x509_D8_number; // @[package.scala 96:25:@26613.4 package.scala 96:25:@26614.4]
  wire [31:0] x546_x305_sum_D7_number; // @[package.scala 96:25:@26631.4 package.scala 96:25:@26632.4]
  wire [31:0] x549_x299_sum_D7_number; // @[package.scala 96:25:@26697.4 package.scala 96:25:@26698.4]
  wire [31:0] x550_x505_D9_number; // @[package.scala 96:25:@26706.4 package.scala 96:25:@26707.4]
  wire [31:0] x552_x325_sum_D1_number; // @[package.scala 96:25:@26811.4 package.scala 96:25:@26812.4]
  wire [31:0] x553_x510_D2_number; // @[package.scala 96:25:@26820.4 package.scala 96:25:@26821.4]
  wire [31:0] x555_x511_D2_number; // @[package.scala 96:25:@26925.4 package.scala 96:25:@26926.4]
  wire [31:0] x556_x334_sum_D1_number; // @[package.scala 96:25:@26934.4 package.scala 96:25:@26935.4]
  wire [31:0] x345_sum_number; // @[Math.scala 154:22:@27070.4 Math.scala 155:14:@27071.4]
  wire [31:0] x559_x513_D2_number; // @[package.scala 96:25:@27079.4 package.scala 96:25:@27080.4]
  wire [31:0] x350_sum_number; // @[Math.scala 154:22:@27148.4 Math.scala 155:14:@27149.4]
  wire [31:0] x355_sum_number; // @[Math.scala 154:22:@27206.4 Math.scala 155:14:@27207.4]
  wire [31:0] x360_sum_number; // @[Math.scala 154:22:@27264.4 Math.scala 155:14:@27265.4]
  wire [31:0] x371_sum_number; // @[Math.scala 154:22:@27391.4 Math.scala 155:14:@27392.4]
  wire [31:0] x568_x518_D2_number; // @[package.scala 96:25:@27400.4 package.scala 96:25:@27401.4]
  wire [31:0] x376_sum_number; // @[Math.scala 154:22:@27449.4 Math.scala 155:14:@27450.4]
  wire [31:0] x381_sum_number; // @[Math.scala 154:22:@27498.4 Math.scala 155:14:@27499.4]
  wire [31:0] x386_sum_number; // @[Math.scala 154:22:@27549.4 Math.scala 155:14:@27550.4]
  wire [32:0] _T_1143; // @[package.scala 96:25:@27593.4 package.scala 96:25:@27594.4]
  wire [32:0] _T_1148; // @[package.scala 96:25:@27605.4 package.scala 96:25:@27606.4]
  wire [33:0] _T_1153; // @[package.scala 96:25:@27617.4 package.scala 96:25:@27618.4]
  wire [32:0] _T_1158; // @[package.scala 96:25:@27629.4 package.scala 96:25:@27630.4]
  wire [32:0] _T_1163; // @[package.scala 96:25:@27641.4 package.scala 96:25:@27642.4]
  wire [32:0] _T_1268; // @[package.scala 96:25:@27904.4 package.scala 96:25:@27905.4]
  wire [32:0] _T_1273; // @[package.scala 96:25:@27916.4 package.scala 96:25:@27917.4]
  wire [33:0] _T_1278; // @[package.scala 96:25:@27928.4 package.scala 96:25:@27929.4]
  wire [32:0] _T_1283; // @[package.scala 96:25:@27940.4 package.scala 96:25:@27941.4]
  wire [32:0] _T_1288; // @[package.scala 96:25:@27952.4 package.scala 96:25:@27953.4]
  _ _ ( // @[Math.scala 720:24:@26101.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@26113.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@26136.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x290_lb_0 x290_lb_0 ( // @[m_x290_lb_0.scala 39:17:@26146.4]
    .clock(x290_lb_0_clock),
    .reset(x290_lb_0_reset),
    .io_rPort_11_banks_1(x290_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x290_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x290_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x290_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x290_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x290_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x290_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x290_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x290_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x290_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x290_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x290_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x290_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x290_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x290_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x290_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x290_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x290_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x290_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x290_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x290_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x290_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x290_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x290_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x290_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x290_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x290_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x290_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x290_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x290_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x290_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x290_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x290_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x290_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x290_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x290_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x290_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x290_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x290_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x290_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x290_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x290_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x290_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x290_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x290_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x290_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x290_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x290_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x290_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x290_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x290_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x290_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x290_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x290_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x290_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x290_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x290_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x290_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x290_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x290_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x290_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x290_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x290_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x290_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x290_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x290_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x290_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x290_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x290_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x290_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x290_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x290_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x290_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x290_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x290_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x290_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x290_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x290_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x290_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x290_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x290_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x290_lb_0_io_wPort_0_en_0)
  );
  x496_sub x508_sub_1 ( // @[Math.scala 191:24:@26309.4]
    .clock(x508_sub_1_clock),
    .reset(x508_sub_1_reset),
    .io_a(x508_sub_1_io_a),
    .io_b(x508_sub_1_io_b),
    .io_flow(x508_sub_1_io_flow),
    .io_result(x508_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@26336.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x267_sum x299_sum_1 ( // @[Math.scala 150:24:@26345.4]
    .clock(x299_sum_1_clock),
    .reset(x299_sum_1_reset),
    .io_a(x299_sum_1_io_a),
    .io_b(x299_sum_1_io_b),
    .io_flow(x299_sum_1_io_flow),
    .io_result(x299_sum_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_2 ( // @[package.scala 93:22:@26355.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_3 ( // @[package.scala 93:22:@26364.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_4 ( // @[package.scala 93:22:@26373.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@26382.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_168 RetimeWrapper_6 ( // @[package.scala 93:22:@26391.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_7 ( // @[package.scala 93:22:@26400.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_8 ( // @[package.scala 93:22:@26411.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x267_sum x301_rdcol_1 ( // @[Math.scala 150:24:@26434.4]
    .clock(x301_rdcol_1_clock),
    .reset(x301_rdcol_1_reset),
    .io_a(x301_rdcol_1_io_a),
    .io_b(x301_rdcol_1_io_b),
    .io_flow(x301_rdcol_1_io_flow),
    .io_result(x301_rdcol_1_io_result)
  );
  x267_sum x305_sum_1 ( // @[Math.scala 150:24:@26474.4]
    .clock(x305_sum_1_clock),
    .reset(x305_sum_1_reset),
    .io_a(x305_sum_1_io_a),
    .io_b(x305_sum_1_io_b),
    .io_flow(x305_sum_1_io_flow),
    .io_result(x305_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_9 ( // @[package.scala 93:22:@26484.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_10 ( // @[package.scala 93:22:@26493.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_11 ( // @[package.scala 93:22:@26502.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_12 ( // @[package.scala 93:22:@26513.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_13 ( // @[package.scala 93:22:@26534.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_14 ( // @[package.scala 93:22:@26550.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@26566.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_184 RetimeWrapper_16 ( // @[package.scala 93:22:@26581.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@26590.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_18 ( // @[package.scala 93:22:@26599.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_19 ( // @[package.scala 93:22:@26608.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_20 ( // @[package.scala 93:22:@26617.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_21 ( // @[package.scala 93:22:@26626.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_22 ( // @[package.scala 93:22:@26638.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_23 ( // @[package.scala 93:22:@26659.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_24 ( // @[package.scala 93:22:@26683.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_25 ( // @[package.scala 93:22:@26692.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_184 RetimeWrapper_26 ( // @[package.scala 93:22:@26701.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_27 ( // @[package.scala 93:22:@26713.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x267_sum x319_rdcol_1 ( // @[Math.scala 150:24:@26736.4]
    .clock(x319_rdcol_1_clock),
    .reset(x319_rdcol_1_reset),
    .io_a(x319_rdcol_1_io_a),
    .io_b(x319_rdcol_1_io_b),
    .io_flow(x319_rdcol_1_io_flow),
    .io_result(x319_rdcol_1_io_result)
  );
  RetimeWrapper_181 RetimeWrapper_28 ( // @[package.scala 93:22:@26787.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x267_sum x325_sum_1 ( // @[Math.scala 150:24:@26796.4]
    .clock(x325_sum_1_clock),
    .reset(x325_sum_1_reset),
    .io_a(x325_sum_1_io_a),
    .io_b(x325_sum_1_io_b),
    .io_flow(x325_sum_1_io_flow),
    .io_result(x325_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_29 ( // @[package.scala 93:22:@26806.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_30 ( // @[package.scala 93:22:@26815.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@26824.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_32 ( // @[package.scala 93:22:@26836.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x267_sum x328_rdcol_1 ( // @[Math.scala 150:24:@26859.4]
    .clock(x328_rdcol_1_clock),
    .reset(x328_rdcol_1_reset),
    .io_a(x328_rdcol_1_io_a),
    .io_b(x328_rdcol_1_io_b),
    .io_flow(x328_rdcol_1_io_flow),
    .io_result(x328_rdcol_1_io_result)
  );
  x267_sum x334_sum_1 ( // @[Math.scala 150:24:@26910.4]
    .clock(x334_sum_1_clock),
    .reset(x334_sum_1_reset),
    .io_a(x334_sum_1_io_a),
    .io_b(x334_sum_1_io_b),
    .io_flow(x334_sum_1_io_flow),
    .io_result(x334_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_33 ( // @[package.scala 93:22:@26920.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_34 ( // @[package.scala 93:22:@26929.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@26938.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_36 ( // @[package.scala 93:22:@26950.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x496_sub x337_rdrow_1 ( // @[Math.scala 191:24:@26973.4]
    .clock(x337_rdrow_1_clock),
    .reset(x337_rdrow_1_reset),
    .io_a(x337_rdrow_1_io_a),
    .io_b(x337_rdrow_1_io_b),
    .io_flow(x337_rdrow_1_io_flow),
    .io_result(x337_rdrow_1_io_result)
  );
  x496_sub x516_sub_1 ( // @[Math.scala 191:24:@27045.4]
    .clock(x516_sub_1_clock),
    .reset(x516_sub_1_reset),
    .io_a(x516_sub_1_io_a),
    .io_b(x516_sub_1_io_b),
    .io_flow(x516_sub_1_io_flow),
    .io_result(x516_sub_1_io_result)
  );
  RetimeWrapper_189 RetimeWrapper_37 ( // @[package.scala 93:22:@27055.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x267_sum x345_sum_1 ( // @[Math.scala 150:24:@27064.4]
    .clock(x345_sum_1_clock),
    .reset(x345_sum_1_reset),
    .io_a(x345_sum_1_io_a),
    .io_b(x345_sum_1_io_b),
    .io_flow(x345_sum_1_io_flow),
    .io_result(x345_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_38 ( // @[package.scala 93:22:@27074.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@27083.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_40 ( // @[package.scala 93:22:@27095.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@27116.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_42 ( // @[package.scala 93:22:@27131.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  x267_sum x350_sum_1 ( // @[Math.scala 150:24:@27142.4]
    .clock(x350_sum_1_clock),
    .reset(x350_sum_1_reset),
    .io_a(x350_sum_1_io_a),
    .io_b(x350_sum_1_io_b),
    .io_flow(x350_sum_1_io_flow),
    .io_result(x350_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@27152.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_44 ( // @[package.scala 93:22:@27164.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_45 ( // @[package.scala 93:22:@27191.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x267_sum x355_sum_1 ( // @[Math.scala 150:24:@27200.4]
    .clock(x355_sum_1_clock),
    .reset(x355_sum_1_reset),
    .io_a(x355_sum_1_io_a),
    .io_b(x355_sum_1_io_b),
    .io_flow(x355_sum_1_io_flow),
    .io_result(x355_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@27210.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_47 ( // @[package.scala 93:22:@27222.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_48 ( // @[package.scala 93:22:@27249.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x267_sum x360_sum_1 ( // @[Math.scala 150:24:@27258.4]
    .clock(x360_sum_1_clock),
    .reset(x360_sum_1_reset),
    .io_a(x360_sum_1_io_a),
    .io_b(x360_sum_1_io_b),
    .io_flow(x360_sum_1_io_flow),
    .io_result(x360_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@27268.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_50 ( // @[package.scala 93:22:@27280.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x496_sub x363_rdrow_1 ( // @[Math.scala 191:24:@27303.4]
    .clock(x363_rdrow_1_clock),
    .reset(x363_rdrow_1_reset),
    .io_a(x363_rdrow_1_io_a),
    .io_b(x363_rdrow_1_io_b),
    .io_flow(x363_rdrow_1_io_flow),
    .io_result(x363_rdrow_1_io_result)
  );
  x496_sub x521_sub_1 ( // @[Math.scala 191:24:@27375.4]
    .clock(x521_sub_1_clock),
    .reset(x521_sub_1_reset),
    .io_a(x521_sub_1_io_a),
    .io_b(x521_sub_1_io_b),
    .io_flow(x521_sub_1_io_flow),
    .io_result(x521_sub_1_io_result)
  );
  x267_sum x371_sum_1 ( // @[Math.scala 150:24:@27385.4]
    .clock(x371_sum_1_clock),
    .reset(x371_sum_1_reset),
    .io_a(x371_sum_1_io_a),
    .io_b(x371_sum_1_io_b),
    .io_flow(x371_sum_1_io_flow),
    .io_result(x371_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_51 ( // @[package.scala 93:22:@27395.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@27404.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_53 ( // @[package.scala 93:22:@27416.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x267_sum x376_sum_1 ( // @[Math.scala 150:24:@27443.4]
    .clock(x376_sum_1_clock),
    .reset(x376_sum_1_reset),
    .io_a(x376_sum_1_io_a),
    .io_b(x376_sum_1_io_b),
    .io_flow(x376_sum_1_io_flow),
    .io_result(x376_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@27453.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_55 ( // @[package.scala 93:22:@27465.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x267_sum x381_sum_1 ( // @[Math.scala 150:24:@27492.4]
    .clock(x381_sum_1_clock),
    .reset(x381_sum_1_reset),
    .io_a(x381_sum_1_io_a),
    .io_b(x381_sum_1_io_b),
    .io_flow(x381_sum_1_io_flow),
    .io_result(x381_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@27502.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_57 ( // @[package.scala 93:22:@27514.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x267_sum x386_sum_1 ( // @[Math.scala 150:24:@27543.4]
    .clock(x386_sum_1_clock),
    .reset(x386_sum_1_reset),
    .io_a(x386_sum_1_io_a),
    .io_b(x386_sum_1_io_b),
    .io_flow(x386_sum_1_io_flow),
    .io_result(x386_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@27553.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_59 ( // @[package.scala 93:22:@27565.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_60 ( // @[package.scala 93:22:@27588.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_61 ( // @[package.scala 93:22:@27600.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_62 ( // @[package.scala 93:22:@27612.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_63 ( // @[package.scala 93:22:@27624.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_64 ( // @[package.scala 93:22:@27636.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_65 ( // @[package.scala 93:22:@27646.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x394_x13 x394_x13_1 ( // @[Math.scala 150:24:@27655.4]
    .clock(x394_x13_1_clock),
    .reset(x394_x13_1_reset),
    .io_a(x394_x13_1_io_a),
    .io_b(x394_x13_1_io_b),
    .io_flow(x394_x13_1_io_flow),
    .io_result(x394_x13_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_66 ( // @[package.scala 93:22:@27665.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x394_x13 x395_x14_1 ( // @[Math.scala 150:24:@27674.4]
    .clock(x395_x14_1_clock),
    .reset(x395_x14_1_reset),
    .io_a(x395_x14_1_io_a),
    .io_b(x395_x14_1_io_b),
    .io_flow(x395_x14_1_io_flow),
    .io_result(x395_x14_1_io_result)
  );
  x394_x13 x396_x13_1 ( // @[Math.scala 150:24:@27684.4]
    .clock(x396_x13_1_clock),
    .reset(x396_x13_1_reset),
    .io_a(x396_x13_1_io_a),
    .io_b(x396_x13_1_io_b),
    .io_flow(x396_x13_1_io_flow),
    .io_result(x396_x13_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_67 ( // @[package.scala 93:22:@27694.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x394_x13 x397_x14_1 ( // @[Math.scala 150:24:@27703.4]
    .clock(x397_x14_1_clock),
    .reset(x397_x14_1_reset),
    .io_a(x397_x14_1_io_a),
    .io_b(x397_x14_1_io_b),
    .io_flow(x397_x14_1_io_flow),
    .io_result(x397_x14_1_io_result)
  );
  x394_x13 x398_x13_1 ( // @[Math.scala 150:24:@27713.4]
    .clock(x398_x13_1_clock),
    .reset(x398_x13_1_reset),
    .io_a(x398_x13_1_io_a),
    .io_b(x398_x13_1_io_b),
    .io_flow(x398_x13_1_io_flow),
    .io_result(x398_x13_1_io_result)
  );
  x394_x13 x399_x14_1 ( // @[Math.scala 150:24:@27723.4]
    .clock(x399_x14_1_clock),
    .reset(x399_x14_1_reset),
    .io_a(x399_x14_1_io_a),
    .io_b(x399_x14_1_io_b),
    .io_flow(x399_x14_1_io_flow),
    .io_result(x399_x14_1_io_result)
  );
  x394_x13 x400_x13_1 ( // @[Math.scala 150:24:@27733.4]
    .clock(x400_x13_1_clock),
    .reset(x400_x13_1_reset),
    .io_a(x400_x13_1_io_a),
    .io_b(x400_x13_1_io_b),
    .io_flow(x400_x13_1_io_flow),
    .io_result(x400_x13_1_io_result)
  );
  RetimeWrapper_259 RetimeWrapper_68 ( // @[package.scala 93:22:@27743.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  x394_x13 x401_sum_1 ( // @[Math.scala 150:24:@27752.4]
    .clock(x401_sum_1_clock),
    .reset(x401_sum_1_reset),
    .io_a(x401_sum_1_io_a),
    .io_b(x401_sum_1_io_b),
    .io_flow(x401_sum_1_io_flow),
    .io_result(x401_sum_1_io_result)
  );
  x402 x402_1 ( // @[Math.scala 720:24:@27762.4]
    .io_b(x402_1_io_b),
    .io_result(x402_1_io_result)
  );
  x403_mul x403_mul_1 ( // @[Math.scala 262:24:@27773.4]
    .clock(x403_mul_1_clock),
    .io_a(x403_mul_1_io_a),
    .io_b(x403_mul_1_io_b),
    .io_flow(x403_mul_1_io_flow),
    .io_result(x403_mul_1_io_result)
  );
  x404 x404_1 ( // @[Math.scala 720:24:@27783.4]
    .io_b(x404_1_io_b),
    .io_result(x404_1_io_result)
  );
  RetimeWrapper_261 RetimeWrapper_69 ( // @[package.scala 93:22:@27792.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x405_sub x405_sub_1 ( // @[Math.scala 191:24:@27801.4]
    .clock(x405_sub_1_clock),
    .reset(x405_sub_1_reset),
    .io_a(x405_sub_1_io_a),
    .io_b(x405_sub_1_io_b),
    .io_flow(x405_sub_1_io_flow),
    .io_result(x405_sub_1_io_result)
  );
  x405_sub x407_sub_1 ( // @[Math.scala 191:24:@27816.4]
    .clock(x407_sub_1_clock),
    .reset(x407_sub_1_reset),
    .io_a(x407_sub_1_io_a),
    .io_b(x407_sub_1_io_b),
    .io_flow(x407_sub_1_io_flow),
    .io_result(x407_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_70 ( // @[package.scala 93:22:@27839.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  x402 x411_1 ( // @[Math.scala 720:24:@27848.4]
    .io_b(x411_1_io_b),
    .io_result(x411_1_io_result)
  );
  x403_mul x412_mul_1 ( // @[Math.scala 262:24:@27859.4]
    .clock(x412_mul_1_clock),
    .io_a(x412_mul_1_io_a),
    .io_b(x412_mul_1_io_b),
    .io_flow(x412_mul_1_io_flow),
    .io_result(x412_mul_1_io_result)
  );
  x404 x413_1 ( // @[Math.scala 720:24:@27869.4]
    .io_b(x413_1_io_b),
    .io_result(x413_1_io_result)
  );
  RetimeWrapper_265 RetimeWrapper_71 ( // @[package.scala 93:22:@27878.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x394_x13 x414_sum_1 ( // @[Math.scala 150:24:@27887.4]
    .clock(x414_sum_1_clock),
    .reset(x414_sum_1_reset),
    .io_a(x414_sum_1_io_a),
    .io_b(x414_sum_1_io_b),
    .io_flow(x414_sum_1_io_flow),
    .io_result(x414_sum_1_io_result)
  );
  RetimeWrapper_244 RetimeWrapper_72 ( // @[package.scala 93:22:@27899.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_73 ( // @[package.scala 93:22:@27911.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_74 ( // @[package.scala 93:22:@27923.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_75 ( // @[package.scala 93:22:@27935.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_244 RetimeWrapper_76 ( // @[package.scala 93:22:@27947.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_77 ( // @[package.scala 93:22:@27957.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x394_x13 x420_x13_1 ( // @[Math.scala 150:24:@27966.4]
    .clock(x420_x13_1_clock),
    .reset(x420_x13_1_reset),
    .io_a(x420_x13_1_io_a),
    .io_b(x420_x13_1_io_b),
    .io_flow(x420_x13_1_io_flow),
    .io_result(x420_x13_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_78 ( // @[package.scala 93:22:@27976.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x394_x13 x421_x14_1 ( // @[Math.scala 150:24:@27985.4]
    .clock(x421_x14_1_clock),
    .reset(x421_x14_1_reset),
    .io_a(x421_x14_1_io_a),
    .io_b(x421_x14_1_io_b),
    .io_flow(x421_x14_1_io_flow),
    .io_result(x421_x14_1_io_result)
  );
  x394_x13 x422_x13_1 ( // @[Math.scala 150:24:@27995.4]
    .clock(x422_x13_1_clock),
    .reset(x422_x13_1_reset),
    .io_a(x422_x13_1_io_a),
    .io_b(x422_x13_1_io_b),
    .io_flow(x422_x13_1_io_flow),
    .io_result(x422_x13_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_79 ( // @[package.scala 93:22:@28005.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  x394_x13 x423_x14_1 ( // @[Math.scala 150:24:@28016.4]
    .clock(x423_x14_1_clock),
    .reset(x423_x14_1_reset),
    .io_a(x423_x14_1_io_a),
    .io_b(x423_x14_1_io_b),
    .io_flow(x423_x14_1_io_flow),
    .io_result(x423_x14_1_io_result)
  );
  x394_x13 x424_x13_1 ( // @[Math.scala 150:24:@28026.4]
    .clock(x424_x13_1_clock),
    .reset(x424_x13_1_reset),
    .io_a(x424_x13_1_io_a),
    .io_b(x424_x13_1_io_b),
    .io_flow(x424_x13_1_io_flow),
    .io_result(x424_x13_1_io_result)
  );
  x394_x13 x425_x14_1 ( // @[Math.scala 150:24:@28036.4]
    .clock(x425_x14_1_clock),
    .reset(x425_x14_1_reset),
    .io_a(x425_x14_1_io_a),
    .io_b(x425_x14_1_io_b),
    .io_flow(x425_x14_1_io_flow),
    .io_result(x425_x14_1_io_result)
  );
  x394_x13 x426_x13_1 ( // @[Math.scala 150:24:@28046.4]
    .clock(x426_x13_1_clock),
    .reset(x426_x13_1_reset),
    .io_a(x426_x13_1_io_a),
    .io_b(x426_x13_1_io_b),
    .io_flow(x426_x13_1_io_flow),
    .io_result(x426_x13_1_io_result)
  );
  RetimeWrapper_259 RetimeWrapper_80 ( // @[package.scala 93:22:@28056.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x394_x13 x427_sum_1 ( // @[Math.scala 150:24:@28065.4]
    .clock(x427_sum_1_clock),
    .reset(x427_sum_1_reset),
    .io_a(x427_sum_1_io_a),
    .io_b(x427_sum_1_io_b),
    .io_flow(x427_sum_1_io_flow),
    .io_result(x427_sum_1_io_result)
  );
  x402 x428_1 ( // @[Math.scala 720:24:@28075.4]
    .io_b(x428_1_io_b),
    .io_result(x428_1_io_result)
  );
  x403_mul x429_mul_1 ( // @[Math.scala 262:24:@28086.4]
    .clock(x429_mul_1_clock),
    .io_a(x429_mul_1_io_a),
    .io_b(x429_mul_1_io_b),
    .io_flow(x429_mul_1_io_flow),
    .io_result(x429_mul_1_io_result)
  );
  x404 x430_1 ( // @[Math.scala 720:24:@28096.4]
    .io_b(x430_1_io_b),
    .io_result(x430_1_io_result)
  );
  RetimeWrapper_261 RetimeWrapper_81 ( // @[package.scala 93:22:@28105.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  x405_sub x431_sub_1 ( // @[Math.scala 191:24:@28114.4]
    .clock(x431_sub_1_clock),
    .reset(x431_sub_1_reset),
    .io_a(x431_sub_1_io_a),
    .io_b(x431_sub_1_io_b),
    .io_flow(x431_sub_1_io_flow),
    .io_result(x431_sub_1_io_result)
  );
  x405_sub x433_sub_1 ( // @[Math.scala 191:24:@28129.4]
    .clock(x433_sub_1_clock),
    .reset(x433_sub_1_reset),
    .io_a(x433_sub_1_io_a),
    .io_b(x433_sub_1_io_b),
    .io_flow(x433_sub_1_io_flow),
    .io_result(x433_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_82 ( // @[package.scala 93:22:@28152.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x402 x437_1 ( // @[Math.scala 720:24:@28161.4]
    .io_b(x437_1_io_b),
    .io_result(x437_1_io_result)
  );
  x403_mul x438_mul_1 ( // @[Math.scala 262:24:@28172.4]
    .clock(x438_mul_1_clock),
    .io_a(x438_mul_1_io_a),
    .io_b(x438_mul_1_io_b),
    .io_flow(x438_mul_1_io_flow),
    .io_result(x438_mul_1_io_result)
  );
  x404 x439_1 ( // @[Math.scala 720:24:@28182.4]
    .io_b(x439_1_io_b),
    .io_result(x439_1_io_result)
  );
  RetimeWrapper_265 RetimeWrapper_83 ( // @[package.scala 93:22:@28191.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  x394_x13 x440_sum_1 ( // @[Math.scala 150:24:@28200.4]
    .clock(x440_sum_1_clock),
    .reset(x440_sum_1_reset),
    .io_a(x440_sum_1_io_a),
    .io_b(x440_sum_1_io_b),
    .io_flow(x440_sum_1_io_flow),
    .io_result(x440_sum_1_io_result)
  );
  RetimeWrapper_290 RetimeWrapper_84 ( // @[package.scala 93:22:@28216.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_85 ( // @[package.scala 93:22:@28225.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_86 ( // @[package.scala 93:22:@28234.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_87 ( // @[package.scala 93:22:@28243.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  assign b286 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 62:18:@26121.4]
  assign b287 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 63:18:@26122.4]
  assign _T_205 = b286 & b287; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 67:30:@26124.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 67:37:@26125.4]
  assign _T_210 = io_in_x253_TID == 8'h0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:76:@26130.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:62:@26131.4]
  assign _T_213 = io_in_x253_TDEST == 8'h0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:101:@26132.4]
  assign x527_x288_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@26141.4 package.scala 96:25:@26142.4]
  assign b284_number = __io_result; // @[Math.scala 723:22:@26106.4 Math.scala 724:14:@26107.4]
  assign _T_243 = $signed(b284_number); // @[Math.scala 406:49:@26250.4]
  assign _T_245 = $signed(_T_243) & $signed(32'sh3); // @[Math.scala 406:56:@26252.4]
  assign _T_246 = $signed(_T_245); // @[Math.scala 406:56:@26253.4]
  assign x503_number = $unsigned(_T_246); // @[implicits.scala 133:21:@26254.4]
  assign _T_256 = $signed(x503_number); // @[Math.scala 406:49:@26263.4]
  assign _T_258 = $signed(_T_256) & $signed(32'sh3); // @[Math.scala 406:56:@26265.4]
  assign _T_259 = $signed(_T_258); // @[Math.scala 406:56:@26266.4]
  assign b285_number = __1_io_result; // @[Math.scala 723:22:@26118.4 Math.scala 724:14:@26119.4]
  assign _T_268 = $signed(b285_number); // @[Math.scala 406:49:@26274.4]
  assign _T_270 = $signed(_T_268) & $signed(32'sh3); // @[Math.scala 406:56:@26276.4]
  assign _T_271 = $signed(_T_270); // @[Math.scala 406:56:@26277.4]
  assign _T_275 = x503_number[31]; // @[FixedPoint.scala 50:25:@26283.4]
  assign _T_279 = _T_275 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26285.4]
  assign _T_280 = x503_number[31:2]; // @[FixedPoint.scala 18:52:@26286.4]
  assign _T_286 = _T_280 == 30'h3fffffff; // @[Math.scala 451:55:@26288.4]
  assign _T_287 = x503_number[1:0]; // @[FixedPoint.scala 18:52:@26289.4]
  assign _T_293 = _T_287 != 2'h0; // @[Math.scala 451:110:@26291.4]
  assign _T_294 = _T_286 & _T_293; // @[Math.scala 451:94:@26292.4]
  assign _T_296 = {_T_279,_T_280}; // @[Cat.scala 30:58:@26294.4]
  assign x296_1_number = _T_294 ? 32'h0 : _T_296; // @[Math.scala 454:20:@26295.4]
  assign _GEN_0 = {{9'd0}, x296_1_number}; // @[Math.scala 461:32:@26300.4]
  assign _T_301 = _GEN_0 << 9; // @[Math.scala 461:32:@26300.4]
  assign _GEN_1 = {{5'd0}, x296_1_number}; // @[Math.scala 461:32:@26305.4]
  assign _T_304 = _GEN_1 << 5; // @[Math.scala 461:32:@26305.4]
  assign _T_310 = b285_number[31]; // @[FixedPoint.scala 50:25:@26320.4]
  assign _T_314 = _T_310 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26322.4]
  assign _T_315 = b285_number[31:2]; // @[FixedPoint.scala 18:52:@26323.4]
  assign _T_321 = _T_315 == 30'h3fffffff; // @[Math.scala 451:55:@26325.4]
  assign _T_322 = b285_number[1:0]; // @[FixedPoint.scala 18:52:@26326.4]
  assign _T_328 = _T_322 != 2'h0; // @[Math.scala 451:110:@26328.4]
  assign _T_329 = _T_321 & _T_328; // @[Math.scala 451:94:@26329.4]
  assign _T_331 = {_T_314,_T_315}; // @[Cat.scala 30:58:@26331.4]
  assign _T_359 = ~ io_sigsIn_break; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:101:@26408.4]
  assign _T_363 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@26416.4 package.scala 96:25:@26417.4]
  assign _T_365 = io_rr ? _T_363 : 1'h0; // @[implicits.scala 55:10:@26418.4]
  assign _T_366 = _T_359 & _T_365; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:118:@26419.4]
  assign _T_368 = _T_366 & _T_359; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:206:@26421.4]
  assign _T_369 = _T_368 & io_sigsIn_backpressure; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:225:@26422.4]
  assign x531_b286_D3 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@26378.4 package.scala 96:25:@26379.4]
  assign _T_370 = _T_369 & x531_b286_D3; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 117:251:@26423.4]
  assign x534_b287_D3 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@26405.4 package.scala 96:25:@26406.4]
  assign x301_rdcol_number = x301_rdcol_1_io_result; // @[Math.scala 154:22:@26440.4 Math.scala 155:14:@26441.4]
  assign _T_387 = $signed(x301_rdcol_number); // @[Math.scala 406:49:@26449.4]
  assign _T_389 = $signed(_T_387) & $signed(32'sh3); // @[Math.scala 406:56:@26451.4]
  assign _T_390 = $signed(_T_389); // @[Math.scala 406:56:@26452.4]
  assign _T_394 = x301_rdcol_number[31]; // @[FixedPoint.scala 50:25:@26458.4]
  assign _T_398 = _T_394 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26460.4]
  assign _T_399 = x301_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@26461.4]
  assign _T_405 = _T_399 == 30'h3fffffff; // @[Math.scala 451:55:@26463.4]
  assign _T_406 = x301_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@26464.4]
  assign _T_412 = _T_406 != 2'h0; // @[Math.scala 451:110:@26466.4]
  assign _T_413 = _T_405 & _T_412; // @[Math.scala 451:94:@26467.4]
  assign _T_415 = {_T_398,_T_399}; // @[Cat.scala 30:58:@26469.4]
  assign _T_435 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@26518.4 package.scala 96:25:@26519.4]
  assign _T_437 = io_rr ? _T_435 : 1'h0; // @[implicits.scala 55:10:@26520.4]
  assign _T_438 = _T_359 & _T_437; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:118:@26521.4]
  assign _T_440 = _T_438 & _T_359; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:206:@26523.4]
  assign _T_441 = _T_440 & io_sigsIn_backpressure; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:225:@26524.4]
  assign _T_442 = _T_441 & x531_b286_D3; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 138:251:@26525.4]
  assign x538_b284_D6_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@26539.4 package.scala 96:25:@26540.4]
  assign _T_452 = $signed(x538_b284_D6_number); // @[Math.scala 476:37:@26545.4]
  assign x308 = $signed(_T_452) < $signed(32'sh0); // @[Math.scala 476:44:@26547.4]
  assign x539_x301_rdcol_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@26555.4 package.scala 96:25:@26556.4]
  assign _T_463 = $signed(x539_x301_rdcol_D6_number); // @[Math.scala 476:37:@26561.4]
  assign x309 = $signed(_T_463) < $signed(32'sh0); // @[Math.scala 476:44:@26563.4]
  assign x540_x308_D1 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@26571.4 package.scala 96:25:@26572.4]
  assign x310 = x540_x308_D1 | x309; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 151:24:@26575.4]
  assign _T_502 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@26643.4 package.scala 96:25:@26644.4]
  assign _T_504 = io_rr ? _T_502 : 1'h0; // @[implicits.scala 55:10:@26645.4]
  assign _T_505 = _T_359 & _T_504; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 170:146:@26646.4]
  assign x542_x311_D2 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@26595.4 package.scala 96:25:@26596.4]
  assign _T_506 = _T_505 & x542_x311_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 170:234:@26647.4]
  assign x543_b286_D9 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@26604.4 package.scala 96:25:@26605.4]
  assign _T_507 = _T_506 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 170:242:@26648.4]
  assign x545_b287_D9 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@26622.4 package.scala 96:25:@26623.4]
  assign x547_b285_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@26664.4 package.scala 96:25:@26665.4]
  assign _T_520 = $signed(x547_b285_D6_number); // @[Math.scala 476:37:@26672.4]
  assign x314 = $signed(_T_520) < $signed(32'sh0); // @[Math.scala 476:44:@26674.4]
  assign x315 = x308 | x314; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 186:59:@26677.4]
  assign _T_547 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@26718.4 package.scala 96:25:@26719.4]
  assign _T_549 = io_rr ? _T_547 : 1'h0; // @[implicits.scala 55:10:@26720.4]
  assign _T_550 = _T_359 & _T_549; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:194:@26721.4]
  assign x548_x316_D3 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@26688.4 package.scala 96:25:@26689.4]
  assign _T_551 = _T_550 & x548_x316_D3; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:282:@26722.4]
  assign _T_552 = _T_551 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:290:@26723.4]
  assign x319_rdcol_number = x319_rdcol_1_io_result; // @[Math.scala 154:22:@26742.4 Math.scala 155:14:@26743.4]
  assign _T_567 = $signed(x319_rdcol_number); // @[Math.scala 476:37:@26748.4]
  assign x320 = $signed(_T_567) < $signed(32'sh0); // @[Math.scala 476:44:@26750.4]
  assign x321 = x540_x308_D1 | x320; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 207:59:@26753.4]
  assign _T_583 = $signed(_T_567) & $signed(32'sh3); // @[Math.scala 406:56:@26764.4]
  assign _T_584 = $signed(_T_583); // @[Math.scala 406:56:@26765.4]
  assign _T_588 = x319_rdcol_number[31]; // @[FixedPoint.scala 50:25:@26771.4]
  assign _T_592 = _T_588 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26773.4]
  assign _T_593 = x319_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@26774.4]
  assign _T_599 = _T_593 == 30'h3fffffff; // @[Math.scala 451:55:@26776.4]
  assign _T_600 = x319_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@26777.4]
  assign _T_606 = _T_600 != 2'h0; // @[Math.scala 451:110:@26779.4]
  assign _T_607 = _T_599 & _T_606; // @[Math.scala 451:94:@26780.4]
  assign _T_609 = {_T_592,_T_593}; // @[Cat.scala 30:58:@26782.4]
  assign _T_638 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@26841.4 package.scala 96:25:@26842.4]
  assign _T_640 = io_rr ? _T_638 : 1'h0; // @[implicits.scala 55:10:@26843.4]
  assign _T_641 = _T_359 & _T_640; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:194:@26844.4]
  assign x554_x322_D2 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@26829.4 package.scala 96:25:@26830.4]
  assign _T_642 = _T_641 & x554_x322_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:282:@26845.4]
  assign _T_643 = _T_642 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:290:@26846.4]
  assign x328_rdcol_number = x328_rdcol_1_io_result; // @[Math.scala 154:22:@26865.4 Math.scala 155:14:@26866.4]
  assign _T_658 = $signed(x328_rdcol_number); // @[Math.scala 476:37:@26871.4]
  assign x329 = $signed(_T_658) < $signed(32'sh0); // @[Math.scala 476:44:@26873.4]
  assign x330 = x540_x308_D1 | x329; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 236:59:@26876.4]
  assign _T_674 = $signed(_T_658) & $signed(32'sh3); // @[Math.scala 406:56:@26887.4]
  assign _T_675 = $signed(_T_674); // @[Math.scala 406:56:@26888.4]
  assign _T_679 = x328_rdcol_number[31]; // @[FixedPoint.scala 50:25:@26894.4]
  assign _T_683 = _T_679 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26896.4]
  assign _T_684 = x328_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@26897.4]
  assign _T_690 = _T_684 == 30'h3fffffff; // @[Math.scala 451:55:@26899.4]
  assign _T_691 = x328_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@26900.4]
  assign _T_697 = _T_691 != 2'h0; // @[Math.scala 451:110:@26902.4]
  assign _T_698 = _T_690 & _T_697; // @[Math.scala 451:94:@26903.4]
  assign _T_700 = {_T_683,_T_684}; // @[Cat.scala 30:58:@26905.4]
  assign _T_726 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@26955.4 package.scala 96:25:@26956.4]
  assign _T_728 = io_rr ? _T_726 : 1'h0; // @[implicits.scala 55:10:@26957.4]
  assign _T_729 = _T_359 & _T_728; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 255:194:@26958.4]
  assign x557_x331_D2 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@26943.4 package.scala 96:25:@26944.4]
  assign _T_730 = _T_729 & x557_x331_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 255:282:@26959.4]
  assign _T_731 = _T_730 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 255:290:@26960.4]
  assign x337_rdrow_number = x337_rdrow_1_io_result; // @[Math.scala 195:22:@26979.4 Math.scala 196:14:@26980.4]
  assign _T_748 = $signed(x337_rdrow_number); // @[Math.scala 406:49:@26986.4]
  assign _T_750 = $signed(_T_748) & $signed(32'sh3); // @[Math.scala 406:56:@26988.4]
  assign _T_751 = $signed(_T_750); // @[Math.scala 406:56:@26989.4]
  assign x512_number = $unsigned(_T_751); // @[implicits.scala 133:21:@26990.4]
  assign x339 = $signed(_T_748) < $signed(32'sh0); // @[Math.scala 476:44:@26998.4]
  assign x340 = x339 | x309; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 265:24:@27001.4]
  assign _T_772 = $signed(x512_number); // @[Math.scala 406:49:@27010.4]
  assign _T_774 = $signed(_T_772) & $signed(32'sh3); // @[Math.scala 406:56:@27012.4]
  assign _T_775 = $signed(_T_774); // @[Math.scala 406:56:@27013.4]
  assign _T_779 = x512_number[31]; // @[FixedPoint.scala 50:25:@27019.4]
  assign _T_783 = _T_779 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27021.4]
  assign _T_784 = x512_number[31:2]; // @[FixedPoint.scala 18:52:@27022.4]
  assign _T_790 = _T_784 == 30'h3fffffff; // @[Math.scala 451:55:@27024.4]
  assign _T_791 = x512_number[1:0]; // @[FixedPoint.scala 18:52:@27025.4]
  assign _T_797 = _T_791 != 2'h0; // @[Math.scala 451:110:@27027.4]
  assign _T_798 = _T_790 & _T_797; // @[Math.scala 451:94:@27028.4]
  assign _T_800 = {_T_783,_T_784}; // @[Cat.scala 30:58:@27030.4]
  assign x343_1_number = _T_798 ? 32'h0 : _T_800; // @[Math.scala 454:20:@27031.4]
  assign _GEN_2 = {{9'd0}, x343_1_number}; // @[Math.scala 461:32:@27036.4]
  assign _T_805 = _GEN_2 << 9; // @[Math.scala 461:32:@27036.4]
  assign _GEN_3 = {{5'd0}, x343_1_number}; // @[Math.scala 461:32:@27041.4]
  assign _T_808 = _GEN_3 << 5; // @[Math.scala 461:32:@27041.4]
  assign _T_835 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@27100.4 package.scala 96:25:@27101.4]
  assign _T_837 = io_rr ? _T_835 : 1'h0; // @[implicits.scala 55:10:@27102.4]
  assign _T_838 = _T_359 & _T_837; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:194:@27103.4]
  assign x560_x341_D2 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@27088.4 package.scala 96:25:@27089.4]
  assign _T_839 = _T_838 & x560_x341_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:282:@27104.4]
  assign _T_840 = _T_839 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:290:@27105.4]
  assign x561_x314_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@27121.4 package.scala 96:25:@27122.4]
  assign x348 = x339 | x561_x314_D1; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 302:59:@27125.4]
  assign _T_872 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@27169.4 package.scala 96:25:@27170.4]
  assign _T_874 = io_rr ? _T_872 : 1'h0; // @[implicits.scala 55:10:@27171.4]
  assign _T_875 = _T_359 & _T_874; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:194:@27172.4]
  assign x563_x349_D2 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@27157.4 package.scala 96:25:@27158.4]
  assign _T_876 = _T_875 & x563_x349_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:282:@27173.4]
  assign _T_877 = _T_876 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:290:@27174.4]
  assign x353 = x339 | x320; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 321:59:@27185.4]
  assign _T_904 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@27227.4 package.scala 96:25:@27228.4]
  assign _T_906 = io_rr ? _T_904 : 1'h0; // @[implicits.scala 55:10:@27229.4]
  assign _T_907 = _T_359 & _T_906; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:194:@27230.4]
  assign x565_x354_D2 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@27215.4 package.scala 96:25:@27216.4]
  assign _T_908 = _T_907 & x565_x354_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:282:@27231.4]
  assign _T_909 = _T_908 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:290:@27232.4]
  assign x358 = x339 | x329; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 338:59:@27243.4]
  assign _T_936 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@27285.4 package.scala 96:25:@27286.4]
  assign _T_938 = io_rr ? _T_936 : 1'h0; // @[implicits.scala 55:10:@27287.4]
  assign _T_939 = _T_359 & _T_938; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:194:@27288.4]
  assign x567_x359_D2 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@27273.4 package.scala 96:25:@27274.4]
  assign _T_940 = _T_939 & x567_x359_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:282:@27289.4]
  assign _T_941 = _T_940 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:290:@27290.4]
  assign x363_rdrow_number = x363_rdrow_1_io_result; // @[Math.scala 195:22:@27309.4 Math.scala 196:14:@27310.4]
  assign _T_958 = $signed(x363_rdrow_number); // @[Math.scala 406:49:@27316.4]
  assign _T_960 = $signed(_T_958) & $signed(32'sh3); // @[Math.scala 406:56:@27318.4]
  assign _T_961 = $signed(_T_960); // @[Math.scala 406:56:@27319.4]
  assign x517_number = $unsigned(_T_961); // @[implicits.scala 133:21:@27320.4]
  assign x365 = $signed(_T_958) < $signed(32'sh0); // @[Math.scala 476:44:@27328.4]
  assign x366 = x365 | x309; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 361:24:@27331.4]
  assign _T_982 = $signed(x517_number); // @[Math.scala 406:49:@27340.4]
  assign _T_984 = $signed(_T_982) & $signed(32'sh3); // @[Math.scala 406:56:@27342.4]
  assign _T_985 = $signed(_T_984); // @[Math.scala 406:56:@27343.4]
  assign _T_989 = x517_number[31]; // @[FixedPoint.scala 50:25:@27349.4]
  assign _T_993 = _T_989 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27351.4]
  assign _T_994 = x517_number[31:2]; // @[FixedPoint.scala 18:52:@27352.4]
  assign _T_1000 = _T_994 == 30'h3fffffff; // @[Math.scala 451:55:@27354.4]
  assign _T_1001 = x517_number[1:0]; // @[FixedPoint.scala 18:52:@27355.4]
  assign _T_1007 = _T_1001 != 2'h0; // @[Math.scala 451:110:@27357.4]
  assign _T_1008 = _T_1000 & _T_1007; // @[Math.scala 451:94:@27358.4]
  assign _T_1010 = {_T_993,_T_994}; // @[Cat.scala 30:58:@27360.4]
  assign x369_1_number = _T_1008 ? 32'h0 : _T_1010; // @[Math.scala 454:20:@27361.4]
  assign _GEN_4 = {{9'd0}, x369_1_number}; // @[Math.scala 461:32:@27366.4]
  assign _T_1015 = _GEN_4 << 9; // @[Math.scala 461:32:@27366.4]
  assign _GEN_5 = {{5'd0}, x369_1_number}; // @[Math.scala 461:32:@27371.4]
  assign _T_1018 = _GEN_5 << 5; // @[Math.scala 461:32:@27371.4]
  assign _T_1042 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@27421.4 package.scala 96:25:@27422.4]
  assign _T_1044 = io_rr ? _T_1042 : 1'h0; // @[implicits.scala 55:10:@27423.4]
  assign _T_1045 = _T_359 & _T_1044; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 384:194:@27424.4]
  assign x569_x367_D2 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@27409.4 package.scala 96:25:@27410.4]
  assign _T_1046 = _T_1045 & x569_x367_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 384:282:@27425.4]
  assign _T_1047 = _T_1046 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 384:290:@27426.4]
  assign x374 = x365 | x561_x314_D1; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 388:24:@27437.4]
  assign _T_1071 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@27470.4 package.scala 96:25:@27471.4]
  assign _T_1073 = io_rr ? _T_1071 : 1'h0; // @[implicits.scala 55:10:@27472.4]
  assign _T_1074 = _T_359 & _T_1073; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:194:@27473.4]
  assign x570_x375_D2 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@27458.4 package.scala 96:25:@27459.4]
  assign _T_1075 = _T_1074 & x570_x375_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:282:@27474.4]
  assign _T_1076 = _T_1075 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:290:@27475.4]
  assign x379 = x365 | x320; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 403:24:@27486.4]
  assign _T_1100 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@27519.4 package.scala 96:25:@27520.4]
  assign _T_1102 = io_rr ? _T_1100 : 1'h0; // @[implicits.scala 55:10:@27521.4]
  assign _T_1103 = _T_359 & _T_1102; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:194:@27522.4]
  assign x571_x380_D2 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@27507.4 package.scala 96:25:@27508.4]
  assign _T_1104 = _T_1103 & x571_x380_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:282:@27523.4]
  assign _T_1105 = _T_1104 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:290:@27524.4]
  assign x384 = x365 | x329; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 424:59:@27535.4]
  assign _T_1131 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@27570.4 package.scala 96:25:@27571.4]
  assign _T_1133 = io_rr ? _T_1131 : 1'h0; // @[implicits.scala 55:10:@27572.4]
  assign _T_1134 = _T_359 & _T_1133; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 437:194:@27573.4]
  assign x572_x385_D2 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@27558.4 package.scala 96:25:@27559.4]
  assign _T_1135 = _T_1134 & x572_x385_D2; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 437:282:@27574.4]
  assign _T_1136 = _T_1135 & x543_b286_D9; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 437:290:@27575.4]
  assign x317_rd_0_number = x290_lb_0_io_rPort_3_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 195:29:@26709.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 199:407:@26730.4]
  assign _GEN_6 = {{1'd0}, x317_rd_0_number}; // @[Math.scala 461:32:@27587.4]
  assign x346_rd_0_number = x290_lb_0_io_rPort_10_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 286:29:@27091.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 290:407:@27112.4]
  assign _GEN_7 = {{1'd0}, x346_rd_0_number}; // @[Math.scala 461:32:@27599.4]
  assign x351_rd_0_number = x290_lb_0_io_rPort_9_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 313:29:@27160.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 317:407:@27181.4]
  assign _GEN_8 = {{2'd0}, x351_rd_0_number}; // @[Math.scala 461:32:@27611.4]
  assign x356_rd_0_number = x290_lb_0_io_rPort_4_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 330:29:@27218.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 334:407:@27239.4]
  assign _GEN_9 = {{1'd0}, x356_rd_0_number}; // @[Math.scala 461:32:@27623.4]
  assign x377_rd_0_number = x290_lb_0_io_rPort_7_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 395:29:@27461.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 399:407:@27482.4]
  assign _GEN_10 = {{1'd0}, x377_rd_0_number}; // @[Math.scala 461:32:@27635.4]
  assign x405_sub_number = x405_sub_1_io_result; // @[Math.scala 195:22:@27807.4 Math.scala 196:14:@27808.4]
  assign x406 = 32'hf < x405_sub_number; // @[Math.scala 477:37:@27813.4]
  assign x407_sub_number = x407_sub_1_io_result; // @[Math.scala 195:22:@27822.4 Math.scala 196:14:@27823.4]
  assign x408 = 32'hf < x407_sub_number; // @[Math.scala 477:37:@27828.4]
  assign x409 = x406 | x408; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 491:24:@27831.4]
  assign x326_rd_0_number = x290_lb_0_io_rPort_11_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 224:29:@26832.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 228:407:@26853.4]
  assign _GEN_11 = {{1'd0}, x326_rd_0_number}; // @[Math.scala 461:32:@27898.4]
  assign _GEN_12 = {{1'd0}, x351_rd_0_number}; // @[Math.scala 461:32:@27910.4]
  assign _GEN_13 = {{2'd0}, x356_rd_0_number}; // @[Math.scala 461:32:@27922.4]
  assign x361_rd_0_number = x290_lb_0_io_rPort_2_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 347:29:@27276.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 351:407:@27297.4]
  assign _GEN_14 = {{1'd0}, x361_rd_0_number}; // @[Math.scala 461:32:@27934.4]
  assign x382_rd_0_number = x290_lb_0_io_rPort_5_output_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 410:29:@27510.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 414:407:@27531.4]
  assign _GEN_15 = {{1'd0}, x382_rd_0_number}; // @[Math.scala 461:32:@27946.4]
  assign x431_sub_number = x431_sub_1_io_result; // @[Math.scala 195:22:@28120.4 Math.scala 196:14:@28121.4]
  assign x432 = 32'hf < x431_sub_number; // @[Math.scala 477:37:@28126.4]
  assign x433_sub_number = x433_sub_1_io_result; // @[Math.scala 195:22:@28135.4 Math.scala 196:14:@28136.4]
  assign x434 = 32'hf < x433_sub_number; // @[Math.scala 477:37:@28141.4]
  assign x435 = x432 | x434; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 565:24:@28144.4]
  assign x414_sum_number = x414_sum_1_io_result; // @[Math.scala 154:22:@27893.4 Math.scala 155:14:@27894.4]
  assign x440_sum_number = x440_sum_1_io_result; // @[Math.scala 154:22:@28206.4 Math.scala 155:14:@28207.4]
  assign _T_1412 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@28248.4 package.scala 96:25:@28249.4]
  assign _T_1414 = io_rr ? _T_1412 : 1'h0; // @[implicits.scala 55:10:@28250.4]
  assign x588_b286_D34 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@28239.4 package.scala 96:25:@28240.4]
  assign _T_1415 = _T_1414 & x588_b286_D34; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 589:117:@28251.4]
  assign x587_b287_D34 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@28230.4 package.scala 96:25:@28231.4]
  assign _T_1416 = _T_1415 & x587_b287_D34; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 589:123:@28252.4]
  assign x529_x504_D3_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@26360.4 package.scala 96:25:@26361.4]
  assign x532_x299_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@26387.4 package.scala 96:25:@26388.4]
  assign x533_x505_D3_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@26396.4 package.scala 96:25:@26397.4]
  assign x536_x509_D2_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@26498.4 package.scala 96:25:@26499.4]
  assign x537_x305_sum_D1_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@26507.4 package.scala 96:25:@26508.4]
  assign x541_x504_D9_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@26586.4 package.scala 96:25:@26587.4]
  assign x544_x509_D8_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@26613.4 package.scala 96:25:@26614.4]
  assign x546_x305_sum_D7_number = RetimeWrapper_21_io_out; // @[package.scala 96:25:@26631.4 package.scala 96:25:@26632.4]
  assign x549_x299_sum_D7_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@26697.4 package.scala 96:25:@26698.4]
  assign x550_x505_D9_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@26706.4 package.scala 96:25:@26707.4]
  assign x552_x325_sum_D1_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@26811.4 package.scala 96:25:@26812.4]
  assign x553_x510_D2_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@26820.4 package.scala 96:25:@26821.4]
  assign x555_x511_D2_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@26925.4 package.scala 96:25:@26926.4]
  assign x556_x334_sum_D1_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@26934.4 package.scala 96:25:@26935.4]
  assign x345_sum_number = x345_sum_1_io_result; // @[Math.scala 154:22:@27070.4 Math.scala 155:14:@27071.4]
  assign x559_x513_D2_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@27079.4 package.scala 96:25:@27080.4]
  assign x350_sum_number = x350_sum_1_io_result; // @[Math.scala 154:22:@27148.4 Math.scala 155:14:@27149.4]
  assign x355_sum_number = x355_sum_1_io_result; // @[Math.scala 154:22:@27206.4 Math.scala 155:14:@27207.4]
  assign x360_sum_number = x360_sum_1_io_result; // @[Math.scala 154:22:@27264.4 Math.scala 155:14:@27265.4]
  assign x371_sum_number = x371_sum_1_io_result; // @[Math.scala 154:22:@27391.4 Math.scala 155:14:@27392.4]
  assign x568_x518_D2_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@27400.4 package.scala 96:25:@27401.4]
  assign x376_sum_number = x376_sum_1_io_result; // @[Math.scala 154:22:@27449.4 Math.scala 155:14:@27450.4]
  assign x381_sum_number = x381_sum_1_io_result; // @[Math.scala 154:22:@27498.4 Math.scala 155:14:@27499.4]
  assign x386_sum_number = x386_sum_1_io_result; // @[Math.scala 154:22:@27549.4 Math.scala 155:14:@27550.4]
  assign _T_1143 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@27593.4 package.scala 96:25:@27594.4]
  assign _T_1148 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@27605.4 package.scala 96:25:@27606.4]
  assign _T_1153 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@27617.4 package.scala 96:25:@27618.4]
  assign _T_1158 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@27629.4 package.scala 96:25:@27630.4]
  assign _T_1163 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@27641.4 package.scala 96:25:@27642.4]
  assign _T_1268 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@27904.4 package.scala 96:25:@27905.4]
  assign _T_1273 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@27916.4 package.scala 96:25:@27917.4]
  assign _T_1278 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@27928.4 package.scala 96:25:@27929.4]
  assign _T_1283 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@27940.4 package.scala 96:25:@27941.4]
  assign _T_1288 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@27952.4 package.scala 96:25:@27953.4]
  assign io_in_x253_TREADY = _T_211 & _T_213; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 67:22:@26126.4 sm_x445_inr_Foreach_SAMPLER_BOX.scala 69:22:@26134.4]
  assign io_in_x254_TVALID = _T_1416 & io_sigsIn_backpressure; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 589:22:@28254.4]
  assign io_in_x254_TDATA = {{192'd0}, RetimeWrapper_84_io_out}; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 590:24:@28255.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@26104.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@26116.4]
  assign RetimeWrapper_clock = clock; // @[:@26137.4]
  assign RetimeWrapper_reset = reset; // @[:@26138.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26140.4]
  assign RetimeWrapper_io_in = io_in_x253_TDATA[63:0]; // @[package.scala 94:16:@26139.4]
  assign x290_lb_0_clock = clock; // @[:@26147.4]
  assign x290_lb_0_reset = reset; // @[:@26148.4]
  assign x290_lb_0_io_rPort_11_banks_1 = x553_x510_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26849.4]
  assign x290_lb_0_io_rPort_11_banks_0 = x541_x504_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26848.4]
  assign x290_lb_0_io_rPort_11_ofs_0 = x552_x325_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@26850.4]
  assign x290_lb_0_io_rPort_11_en_0 = _T_643 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@26852.4]
  assign x290_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26851.4]
  assign x290_lb_0_io_rPort_10_banks_1 = x544_x509_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@27108.4]
  assign x290_lb_0_io_rPort_10_banks_0 = x559_x513_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27107.4]
  assign x290_lb_0_io_rPort_10_ofs_0 = x345_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27109.4]
  assign x290_lb_0_io_rPort_10_en_0 = _T_840 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27111.4]
  assign x290_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27110.4]
  assign x290_lb_0_io_rPort_9_banks_1 = x550_x505_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27177.4]
  assign x290_lb_0_io_rPort_9_banks_0 = x559_x513_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27176.4]
  assign x290_lb_0_io_rPort_9_ofs_0 = x350_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27178.4]
  assign x290_lb_0_io_rPort_9_en_0 = _T_877 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27180.4]
  assign x290_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27179.4]
  assign x290_lb_0_io_rPort_8_banks_1 = x555_x511_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27578.4]
  assign x290_lb_0_io_rPort_8_banks_0 = x568_x518_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27577.4]
  assign x290_lb_0_io_rPort_8_ofs_0 = x386_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27579.4]
  assign x290_lb_0_io_rPort_8_en_0 = _T_1136 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27581.4]
  assign x290_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27580.4]
  assign x290_lb_0_io_rPort_7_banks_1 = x550_x505_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@27478.4]
  assign x290_lb_0_io_rPort_7_banks_0 = x568_x518_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27477.4]
  assign x290_lb_0_io_rPort_7_ofs_0 = x376_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27479.4]
  assign x290_lb_0_io_rPort_7_en_0 = _T_1076 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27481.4]
  assign x290_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27480.4]
  assign x290_lb_0_io_rPort_6_banks_1 = x555_x511_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26963.4]
  assign x290_lb_0_io_rPort_6_banks_0 = x541_x504_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26962.4]
  assign x290_lb_0_io_rPort_6_ofs_0 = x556_x334_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@26964.4]
  assign x290_lb_0_io_rPort_6_en_0 = _T_731 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@26966.4]
  assign x290_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26965.4]
  assign x290_lb_0_io_rPort_5_banks_1 = x553_x510_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27527.4]
  assign x290_lb_0_io_rPort_5_banks_0 = x568_x518_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27526.4]
  assign x290_lb_0_io_rPort_5_ofs_0 = x381_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27528.4]
  assign x290_lb_0_io_rPort_5_en_0 = _T_1105 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27530.4]
  assign x290_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27529.4]
  assign x290_lb_0_io_rPort_4_banks_1 = x553_x510_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27235.4]
  assign x290_lb_0_io_rPort_4_banks_0 = x559_x513_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27234.4]
  assign x290_lb_0_io_rPort_4_ofs_0 = x355_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27236.4]
  assign x290_lb_0_io_rPort_4_en_0 = _T_909 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27238.4]
  assign x290_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27237.4]
  assign x290_lb_0_io_rPort_3_banks_1 = x550_x505_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26726.4]
  assign x290_lb_0_io_rPort_3_banks_0 = x541_x504_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26725.4]
  assign x290_lb_0_io_rPort_3_ofs_0 = x549_x299_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@26727.4]
  assign x290_lb_0_io_rPort_3_en_0 = _T_552 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@26729.4]
  assign x290_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26728.4]
  assign x290_lb_0_io_rPort_2_banks_1 = x555_x511_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27293.4]
  assign x290_lb_0_io_rPort_2_banks_0 = x559_x513_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27292.4]
  assign x290_lb_0_io_rPort_2_ofs_0 = x360_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27294.4]
  assign x290_lb_0_io_rPort_2_en_0 = _T_941 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27296.4]
  assign x290_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27295.4]
  assign x290_lb_0_io_rPort_1_banks_1 = x544_x509_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@26651.4]
  assign x290_lb_0_io_rPort_1_banks_0 = x541_x504_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26650.4]
  assign x290_lb_0_io_rPort_1_ofs_0 = x546_x305_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@26652.4]
  assign x290_lb_0_io_rPort_1_en_0 = _T_507 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@26654.4]
  assign x290_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26653.4]
  assign x290_lb_0_io_rPort_0_banks_1 = x544_x509_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@27429.4]
  assign x290_lb_0_io_rPort_0_banks_0 = x568_x518_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@27428.4]
  assign x290_lb_0_io_rPort_0_ofs_0 = x371_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@27430.4]
  assign x290_lb_0_io_rPort_0_en_0 = _T_1047 & x545_b287_D9; // @[MemInterfaceType.scala 110:79:@27432.4]
  assign x290_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27431.4]
  assign x290_lb_0_io_wPort_1_banks_1 = x536_x509_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@26528.4]
  assign x290_lb_0_io_wPort_1_banks_0 = x529_x504_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@26527.4]
  assign x290_lb_0_io_wPort_1_ofs_0 = x537_x305_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@26529.4]
  assign x290_lb_0_io_wPort_1_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@26530.4]
  assign x290_lb_0_io_wPort_1_en_0 = _T_442 & x534_b287_D3; // @[MemInterfaceType.scala 93:57:@26532.4]
  assign x290_lb_0_io_wPort_0_banks_1 = x533_x505_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@26426.4]
  assign x290_lb_0_io_wPort_0_banks_0 = x529_x504_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@26425.4]
  assign x290_lb_0_io_wPort_0_ofs_0 = x532_x299_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@26427.4]
  assign x290_lb_0_io_wPort_0_data_0 = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 90:56:@26428.4]
  assign x290_lb_0_io_wPort_0_en_0 = _T_370 & x534_b287_D3; // @[MemInterfaceType.scala 93:57:@26430.4]
  assign x508_sub_1_clock = clock; // @[:@26310.4]
  assign x508_sub_1_reset = reset; // @[:@26311.4]
  assign x508_sub_1_io_a = _T_301[31:0]; // @[Math.scala 192:17:@26312.4]
  assign x508_sub_1_io_b = _T_304[31:0]; // @[Math.scala 193:17:@26313.4]
  assign x508_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@26314.4]
  assign RetimeWrapper_1_clock = clock; // @[:@26337.4]
  assign RetimeWrapper_1_reset = reset; // @[:@26338.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26340.4]
  assign RetimeWrapper_1_io_in = _T_329 ? 32'h0 : _T_331; // @[package.scala 94:16:@26339.4]
  assign x299_sum_1_clock = clock; // @[:@26346.4]
  assign x299_sum_1_reset = reset; // @[:@26347.4]
  assign x299_sum_1_io_a = x508_sub_1_io_result; // @[Math.scala 151:17:@26348.4]
  assign x299_sum_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 152:17:@26349.4]
  assign x299_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26350.4]
  assign RetimeWrapper_2_clock = clock; // @[:@26356.4]
  assign RetimeWrapper_2_reset = reset; // @[:@26357.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26359.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_259); // @[package.scala 94:16:@26358.4]
  assign RetimeWrapper_3_clock = clock; // @[:@26365.4]
  assign RetimeWrapper_3_reset = reset; // @[:@26366.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26368.4]
  assign RetimeWrapper_3_io_in = x527_x288_D1_0_number[31:0]; // @[package.scala 94:16:@26367.4]
  assign RetimeWrapper_4_clock = clock; // @[:@26374.4]
  assign RetimeWrapper_4_reset = reset; // @[:@26375.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26377.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@26376.4]
  assign RetimeWrapper_5_clock = clock; // @[:@26383.4]
  assign RetimeWrapper_5_reset = reset; // @[:@26384.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26386.4]
  assign RetimeWrapper_5_io_in = x299_sum_1_io_result; // @[package.scala 94:16:@26385.4]
  assign RetimeWrapper_6_clock = clock; // @[:@26392.4]
  assign RetimeWrapper_6_reset = reset; // @[:@26393.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26395.4]
  assign RetimeWrapper_6_io_in = $unsigned(_T_271); // @[package.scala 94:16:@26394.4]
  assign RetimeWrapper_7_clock = clock; // @[:@26401.4]
  assign RetimeWrapper_7_reset = reset; // @[:@26402.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26404.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@26403.4]
  assign RetimeWrapper_8_clock = clock; // @[:@26412.4]
  assign RetimeWrapper_8_reset = reset; // @[:@26413.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26415.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26414.4]
  assign x301_rdcol_1_clock = clock; // @[:@26435.4]
  assign x301_rdcol_1_reset = reset; // @[:@26436.4]
  assign x301_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@26437.4]
  assign x301_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@26438.4]
  assign x301_rdcol_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26439.4]
  assign x305_sum_1_clock = clock; // @[:@26475.4]
  assign x305_sum_1_reset = reset; // @[:@26476.4]
  assign x305_sum_1_io_a = x508_sub_1_io_result; // @[Math.scala 151:17:@26477.4]
  assign x305_sum_1_io_b = _T_413 ? 32'h0 : _T_415; // @[Math.scala 152:17:@26478.4]
  assign x305_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26479.4]
  assign RetimeWrapper_9_clock = clock; // @[:@26485.4]
  assign RetimeWrapper_9_reset = reset; // @[:@26486.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26488.4]
  assign RetimeWrapper_9_io_in = x527_x288_D1_0_number[63:32]; // @[package.scala 94:16:@26487.4]
  assign RetimeWrapper_10_clock = clock; // @[:@26494.4]
  assign RetimeWrapper_10_reset = reset; // @[:@26495.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26497.4]
  assign RetimeWrapper_10_io_in = $unsigned(_T_390); // @[package.scala 94:16:@26496.4]
  assign RetimeWrapper_11_clock = clock; // @[:@26503.4]
  assign RetimeWrapper_11_reset = reset; // @[:@26504.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26506.4]
  assign RetimeWrapper_11_io_in = x305_sum_1_io_result; // @[package.scala 94:16:@26505.4]
  assign RetimeWrapper_12_clock = clock; // @[:@26514.4]
  assign RetimeWrapper_12_reset = reset; // @[:@26515.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26517.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26516.4]
  assign RetimeWrapper_13_clock = clock; // @[:@26535.4]
  assign RetimeWrapper_13_reset = reset; // @[:@26536.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26538.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@26537.4]
  assign RetimeWrapper_14_clock = clock; // @[:@26551.4]
  assign RetimeWrapper_14_reset = reset; // @[:@26552.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26554.4]
  assign RetimeWrapper_14_io_in = x301_rdcol_1_io_result; // @[package.scala 94:16:@26553.4]
  assign RetimeWrapper_15_clock = clock; // @[:@26567.4]
  assign RetimeWrapper_15_reset = reset; // @[:@26568.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26570.4]
  assign RetimeWrapper_15_io_in = $signed(_T_452) < $signed(32'sh0); // @[package.scala 94:16:@26569.4]
  assign RetimeWrapper_16_clock = clock; // @[:@26582.4]
  assign RetimeWrapper_16_reset = reset; // @[:@26583.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26585.4]
  assign RetimeWrapper_16_io_in = $unsigned(_T_259); // @[package.scala 94:16:@26584.4]
  assign RetimeWrapper_17_clock = clock; // @[:@26591.4]
  assign RetimeWrapper_17_reset = reset; // @[:@26592.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26594.4]
  assign RetimeWrapper_17_io_in = ~ x310; // @[package.scala 94:16:@26593.4]
  assign RetimeWrapper_18_clock = clock; // @[:@26600.4]
  assign RetimeWrapper_18_reset = reset; // @[:@26601.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26603.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@26602.4]
  assign RetimeWrapper_19_clock = clock; // @[:@26609.4]
  assign RetimeWrapper_19_reset = reset; // @[:@26610.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26612.4]
  assign RetimeWrapper_19_io_in = $unsigned(_T_390); // @[package.scala 94:16:@26611.4]
  assign RetimeWrapper_20_clock = clock; // @[:@26618.4]
  assign RetimeWrapper_20_reset = reset; // @[:@26619.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26621.4]
  assign RetimeWrapper_20_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@26620.4]
  assign RetimeWrapper_21_clock = clock; // @[:@26627.4]
  assign RetimeWrapper_21_reset = reset; // @[:@26628.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26630.4]
  assign RetimeWrapper_21_io_in = x305_sum_1_io_result; // @[package.scala 94:16:@26629.4]
  assign RetimeWrapper_22_clock = clock; // @[:@26639.4]
  assign RetimeWrapper_22_reset = reset; // @[:@26640.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26642.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26641.4]
  assign RetimeWrapper_23_clock = clock; // @[:@26660.4]
  assign RetimeWrapper_23_reset = reset; // @[:@26661.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26663.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@26662.4]
  assign RetimeWrapper_24_clock = clock; // @[:@26684.4]
  assign RetimeWrapper_24_reset = reset; // @[:@26685.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26687.4]
  assign RetimeWrapper_24_io_in = ~ x315; // @[package.scala 94:16:@26686.4]
  assign RetimeWrapper_25_clock = clock; // @[:@26693.4]
  assign RetimeWrapper_25_reset = reset; // @[:@26694.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26696.4]
  assign RetimeWrapper_25_io_in = x299_sum_1_io_result; // @[package.scala 94:16:@26695.4]
  assign RetimeWrapper_26_clock = clock; // @[:@26702.4]
  assign RetimeWrapper_26_reset = reset; // @[:@26703.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26705.4]
  assign RetimeWrapper_26_io_in = $unsigned(_T_271); // @[package.scala 94:16:@26704.4]
  assign RetimeWrapper_27_clock = clock; // @[:@26714.4]
  assign RetimeWrapper_27_reset = reset; // @[:@26715.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26717.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26716.4]
  assign x319_rdcol_1_clock = clock; // @[:@26737.4]
  assign x319_rdcol_1_reset = reset; // @[:@26738.4]
  assign x319_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@26739.4]
  assign x319_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@26740.4]
  assign x319_rdcol_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26741.4]
  assign RetimeWrapper_28_clock = clock; // @[:@26788.4]
  assign RetimeWrapper_28_reset = reset; // @[:@26789.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26791.4]
  assign RetimeWrapper_28_io_in = x508_sub_1_io_result; // @[package.scala 94:16:@26790.4]
  assign x325_sum_1_clock = clock; // @[:@26797.4]
  assign x325_sum_1_reset = reset; // @[:@26798.4]
  assign x325_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@26799.4]
  assign x325_sum_1_io_b = _T_607 ? 32'h0 : _T_609; // @[Math.scala 152:17:@26800.4]
  assign x325_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26801.4]
  assign RetimeWrapper_29_clock = clock; // @[:@26807.4]
  assign RetimeWrapper_29_reset = reset; // @[:@26808.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26810.4]
  assign RetimeWrapper_29_io_in = x325_sum_1_io_result; // @[package.scala 94:16:@26809.4]
  assign RetimeWrapper_30_clock = clock; // @[:@26816.4]
  assign RetimeWrapper_30_reset = reset; // @[:@26817.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26819.4]
  assign RetimeWrapper_30_io_in = $unsigned(_T_584); // @[package.scala 94:16:@26818.4]
  assign RetimeWrapper_31_clock = clock; // @[:@26825.4]
  assign RetimeWrapper_31_reset = reset; // @[:@26826.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26828.4]
  assign RetimeWrapper_31_io_in = ~ x321; // @[package.scala 94:16:@26827.4]
  assign RetimeWrapper_32_clock = clock; // @[:@26837.4]
  assign RetimeWrapper_32_reset = reset; // @[:@26838.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26840.4]
  assign RetimeWrapper_32_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26839.4]
  assign x328_rdcol_1_clock = clock; // @[:@26860.4]
  assign x328_rdcol_1_reset = reset; // @[:@26861.4]
  assign x328_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@26862.4]
  assign x328_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@26863.4]
  assign x328_rdcol_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26864.4]
  assign x334_sum_1_clock = clock; // @[:@26911.4]
  assign x334_sum_1_reset = reset; // @[:@26912.4]
  assign x334_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@26913.4]
  assign x334_sum_1_io_b = _T_698 ? 32'h0 : _T_700; // @[Math.scala 152:17:@26914.4]
  assign x334_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@26915.4]
  assign RetimeWrapper_33_clock = clock; // @[:@26921.4]
  assign RetimeWrapper_33_reset = reset; // @[:@26922.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26924.4]
  assign RetimeWrapper_33_io_in = $unsigned(_T_675); // @[package.scala 94:16:@26923.4]
  assign RetimeWrapper_34_clock = clock; // @[:@26930.4]
  assign RetimeWrapper_34_reset = reset; // @[:@26931.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26933.4]
  assign RetimeWrapper_34_io_in = x334_sum_1_io_result; // @[package.scala 94:16:@26932.4]
  assign RetimeWrapper_35_clock = clock; // @[:@26939.4]
  assign RetimeWrapper_35_reset = reset; // @[:@26940.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26942.4]
  assign RetimeWrapper_35_io_in = ~ x330; // @[package.scala 94:16:@26941.4]
  assign RetimeWrapper_36_clock = clock; // @[:@26951.4]
  assign RetimeWrapper_36_reset = reset; // @[:@26952.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26954.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26953.4]
  assign x337_rdrow_1_clock = clock; // @[:@26974.4]
  assign x337_rdrow_1_reset = reset; // @[:@26975.4]
  assign x337_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@26976.4]
  assign x337_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@26977.4]
  assign x337_rdrow_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@26978.4]
  assign x516_sub_1_clock = clock; // @[:@27046.4]
  assign x516_sub_1_reset = reset; // @[:@27047.4]
  assign x516_sub_1_io_a = _T_805[31:0]; // @[Math.scala 192:17:@27048.4]
  assign x516_sub_1_io_b = _T_808[31:0]; // @[Math.scala 193:17:@27049.4]
  assign x516_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@27050.4]
  assign RetimeWrapper_37_clock = clock; // @[:@27056.4]
  assign RetimeWrapper_37_reset = reset; // @[:@27057.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27059.4]
  assign RetimeWrapper_37_io_in = _T_413 ? 32'h0 : _T_415; // @[package.scala 94:16:@27058.4]
  assign x345_sum_1_clock = clock; // @[:@27065.4]
  assign x345_sum_1_reset = reset; // @[:@27066.4]
  assign x345_sum_1_io_a = x516_sub_1_io_result; // @[Math.scala 151:17:@27067.4]
  assign x345_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@27068.4]
  assign x345_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27069.4]
  assign RetimeWrapper_38_clock = clock; // @[:@27075.4]
  assign RetimeWrapper_38_reset = reset; // @[:@27076.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27078.4]
  assign RetimeWrapper_38_io_in = $unsigned(_T_775); // @[package.scala 94:16:@27077.4]
  assign RetimeWrapper_39_clock = clock; // @[:@27084.4]
  assign RetimeWrapper_39_reset = reset; // @[:@27085.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27087.4]
  assign RetimeWrapper_39_io_in = ~ x340; // @[package.scala 94:16:@27086.4]
  assign RetimeWrapper_40_clock = clock; // @[:@27096.4]
  assign RetimeWrapper_40_reset = reset; // @[:@27097.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27099.4]
  assign RetimeWrapper_40_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27098.4]
  assign RetimeWrapper_41_clock = clock; // @[:@27117.4]
  assign RetimeWrapper_41_reset = reset; // @[:@27118.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27120.4]
  assign RetimeWrapper_41_io_in = $signed(_T_520) < $signed(32'sh0); // @[package.scala 94:16:@27119.4]
  assign RetimeWrapper_42_clock = clock; // @[:@27132.4]
  assign RetimeWrapper_42_reset = reset; // @[:@27133.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27135.4]
  assign RetimeWrapper_42_io_in = _T_329 ? 32'h0 : _T_331; // @[package.scala 94:16:@27134.4]
  assign x350_sum_1_clock = clock; // @[:@27143.4]
  assign x350_sum_1_reset = reset; // @[:@27144.4]
  assign x350_sum_1_io_a = x516_sub_1_io_result; // @[Math.scala 151:17:@27145.4]
  assign x350_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@27146.4]
  assign x350_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27147.4]
  assign RetimeWrapper_43_clock = clock; // @[:@27153.4]
  assign RetimeWrapper_43_reset = reset; // @[:@27154.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27156.4]
  assign RetimeWrapper_43_io_in = ~ x348; // @[package.scala 94:16:@27155.4]
  assign RetimeWrapper_44_clock = clock; // @[:@27165.4]
  assign RetimeWrapper_44_reset = reset; // @[:@27166.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27168.4]
  assign RetimeWrapper_44_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27167.4]
  assign RetimeWrapper_45_clock = clock; // @[:@27192.4]
  assign RetimeWrapper_45_reset = reset; // @[:@27193.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27195.4]
  assign RetimeWrapper_45_io_in = _T_607 ? 32'h0 : _T_609; // @[package.scala 94:16:@27194.4]
  assign x355_sum_1_clock = clock; // @[:@27201.4]
  assign x355_sum_1_reset = reset; // @[:@27202.4]
  assign x355_sum_1_io_a = x516_sub_1_io_result; // @[Math.scala 151:17:@27203.4]
  assign x355_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@27204.4]
  assign x355_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27205.4]
  assign RetimeWrapper_46_clock = clock; // @[:@27211.4]
  assign RetimeWrapper_46_reset = reset; // @[:@27212.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27214.4]
  assign RetimeWrapper_46_io_in = ~ x353; // @[package.scala 94:16:@27213.4]
  assign RetimeWrapper_47_clock = clock; // @[:@27223.4]
  assign RetimeWrapper_47_reset = reset; // @[:@27224.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27226.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27225.4]
  assign RetimeWrapper_48_clock = clock; // @[:@27250.4]
  assign RetimeWrapper_48_reset = reset; // @[:@27251.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27253.4]
  assign RetimeWrapper_48_io_in = _T_698 ? 32'h0 : _T_700; // @[package.scala 94:16:@27252.4]
  assign x360_sum_1_clock = clock; // @[:@27259.4]
  assign x360_sum_1_reset = reset; // @[:@27260.4]
  assign x360_sum_1_io_a = x516_sub_1_io_result; // @[Math.scala 151:17:@27261.4]
  assign x360_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@27262.4]
  assign x360_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27263.4]
  assign RetimeWrapper_49_clock = clock; // @[:@27269.4]
  assign RetimeWrapper_49_reset = reset; // @[:@27270.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27272.4]
  assign RetimeWrapper_49_io_in = ~ x358; // @[package.scala 94:16:@27271.4]
  assign RetimeWrapper_50_clock = clock; // @[:@27281.4]
  assign RetimeWrapper_50_reset = reset; // @[:@27282.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27284.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27283.4]
  assign x363_rdrow_1_clock = clock; // @[:@27304.4]
  assign x363_rdrow_1_reset = reset; // @[:@27305.4]
  assign x363_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@27306.4]
  assign x363_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@27307.4]
  assign x363_rdrow_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@27308.4]
  assign x521_sub_1_clock = clock; // @[:@27376.4]
  assign x521_sub_1_reset = reset; // @[:@27377.4]
  assign x521_sub_1_io_a = _T_1015[31:0]; // @[Math.scala 192:17:@27378.4]
  assign x521_sub_1_io_b = _T_1018[31:0]; // @[Math.scala 193:17:@27379.4]
  assign x521_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@27380.4]
  assign x371_sum_1_clock = clock; // @[:@27386.4]
  assign x371_sum_1_reset = reset; // @[:@27387.4]
  assign x371_sum_1_io_a = x521_sub_1_io_result; // @[Math.scala 151:17:@27388.4]
  assign x371_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@27389.4]
  assign x371_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27390.4]
  assign RetimeWrapper_51_clock = clock; // @[:@27396.4]
  assign RetimeWrapper_51_reset = reset; // @[:@27397.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27399.4]
  assign RetimeWrapper_51_io_in = $unsigned(_T_985); // @[package.scala 94:16:@27398.4]
  assign RetimeWrapper_52_clock = clock; // @[:@27405.4]
  assign RetimeWrapper_52_reset = reset; // @[:@27406.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27408.4]
  assign RetimeWrapper_52_io_in = ~ x366; // @[package.scala 94:16:@27407.4]
  assign RetimeWrapper_53_clock = clock; // @[:@27417.4]
  assign RetimeWrapper_53_reset = reset; // @[:@27418.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27420.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27419.4]
  assign x376_sum_1_clock = clock; // @[:@27444.4]
  assign x376_sum_1_reset = reset; // @[:@27445.4]
  assign x376_sum_1_io_a = x521_sub_1_io_result; // @[Math.scala 151:17:@27446.4]
  assign x376_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@27447.4]
  assign x376_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27448.4]
  assign RetimeWrapper_54_clock = clock; // @[:@27454.4]
  assign RetimeWrapper_54_reset = reset; // @[:@27455.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27457.4]
  assign RetimeWrapper_54_io_in = ~ x374; // @[package.scala 94:16:@27456.4]
  assign RetimeWrapper_55_clock = clock; // @[:@27466.4]
  assign RetimeWrapper_55_reset = reset; // @[:@27467.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27469.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27468.4]
  assign x381_sum_1_clock = clock; // @[:@27493.4]
  assign x381_sum_1_reset = reset; // @[:@27494.4]
  assign x381_sum_1_io_a = x521_sub_1_io_result; // @[Math.scala 151:17:@27495.4]
  assign x381_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@27496.4]
  assign x381_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27497.4]
  assign RetimeWrapper_56_clock = clock; // @[:@27503.4]
  assign RetimeWrapper_56_reset = reset; // @[:@27504.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27506.4]
  assign RetimeWrapper_56_io_in = ~ x379; // @[package.scala 94:16:@27505.4]
  assign RetimeWrapper_57_clock = clock; // @[:@27515.4]
  assign RetimeWrapper_57_reset = reset; // @[:@27516.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27518.4]
  assign RetimeWrapper_57_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27517.4]
  assign x386_sum_1_clock = clock; // @[:@27544.4]
  assign x386_sum_1_reset = reset; // @[:@27545.4]
  assign x386_sum_1_io_a = x521_sub_1_io_result; // @[Math.scala 151:17:@27546.4]
  assign x386_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@27547.4]
  assign x386_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27548.4]
  assign RetimeWrapper_58_clock = clock; // @[:@27554.4]
  assign RetimeWrapper_58_reset = reset; // @[:@27555.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27557.4]
  assign RetimeWrapper_58_io_in = ~ x384; // @[package.scala 94:16:@27556.4]
  assign RetimeWrapper_59_clock = clock; // @[:@27566.4]
  assign RetimeWrapper_59_reset = reset; // @[:@27567.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27569.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27568.4]
  assign RetimeWrapper_60_clock = clock; // @[:@27589.4]
  assign RetimeWrapper_60_reset = reset; // @[:@27590.4]
  assign RetimeWrapper_60_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27592.4]
  assign RetimeWrapper_60_io_in = _GEN_6 << 1; // @[package.scala 94:16:@27591.4]
  assign RetimeWrapper_61_clock = clock; // @[:@27601.4]
  assign RetimeWrapper_61_reset = reset; // @[:@27602.4]
  assign RetimeWrapper_61_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27604.4]
  assign RetimeWrapper_61_io_in = _GEN_7 << 1; // @[package.scala 94:16:@27603.4]
  assign RetimeWrapper_62_clock = clock; // @[:@27613.4]
  assign RetimeWrapper_62_reset = reset; // @[:@27614.4]
  assign RetimeWrapper_62_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27616.4]
  assign RetimeWrapper_62_io_in = _GEN_8 << 2; // @[package.scala 94:16:@27615.4]
  assign RetimeWrapper_63_clock = clock; // @[:@27625.4]
  assign RetimeWrapper_63_reset = reset; // @[:@27626.4]
  assign RetimeWrapper_63_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27628.4]
  assign RetimeWrapper_63_io_in = _GEN_9 << 1; // @[package.scala 94:16:@27627.4]
  assign RetimeWrapper_64_clock = clock; // @[:@27637.4]
  assign RetimeWrapper_64_reset = reset; // @[:@27638.4]
  assign RetimeWrapper_64_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27640.4]
  assign RetimeWrapper_64_io_in = _GEN_10 << 1; // @[package.scala 94:16:@27639.4]
  assign RetimeWrapper_65_clock = clock; // @[:@27647.4]
  assign RetimeWrapper_65_reset = reset; // @[:@27648.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27650.4]
  assign RetimeWrapper_65_io_in = x290_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@27649.4]
  assign x394_x13_1_clock = clock; // @[:@27656.4]
  assign x394_x13_1_reset = reset; // @[:@27657.4]
  assign x394_x13_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@27658.4]
  assign x394_x13_1_io_b = _T_1143[31:0]; // @[Math.scala 152:17:@27659.4]
  assign x394_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27660.4]
  assign RetimeWrapper_66_clock = clock; // @[:@27666.4]
  assign RetimeWrapper_66_reset = reset; // @[:@27667.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27669.4]
  assign RetimeWrapper_66_io_in = x290_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@27668.4]
  assign x395_x14_1_clock = clock; // @[:@27675.4]
  assign x395_x14_1_reset = reset; // @[:@27676.4]
  assign x395_x14_1_io_a = RetimeWrapper_66_io_out; // @[Math.scala 151:17:@27677.4]
  assign x395_x14_1_io_b = _T_1148[31:0]; // @[Math.scala 152:17:@27678.4]
  assign x395_x14_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27679.4]
  assign x396_x13_1_clock = clock; // @[:@27685.4]
  assign x396_x13_1_reset = reset; // @[:@27686.4]
  assign x396_x13_1_io_a = _T_1153[31:0]; // @[Math.scala 151:17:@27687.4]
  assign x396_x13_1_io_b = _T_1158[31:0]; // @[Math.scala 152:17:@27688.4]
  assign x396_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27689.4]
  assign RetimeWrapper_67_clock = clock; // @[:@27695.4]
  assign RetimeWrapper_67_reset = reset; // @[:@27696.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27698.4]
  assign RetimeWrapper_67_io_in = x290_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@27697.4]
  assign x397_x14_1_clock = clock; // @[:@27704.4]
  assign x397_x14_1_reset = reset; // @[:@27705.4]
  assign x397_x14_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@27706.4]
  assign x397_x14_1_io_b = _T_1163[31:0]; // @[Math.scala 152:17:@27707.4]
  assign x397_x14_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27708.4]
  assign x398_x13_1_clock = clock; // @[:@27714.4]
  assign x398_x13_1_reset = reset; // @[:@27715.4]
  assign x398_x13_1_io_a = x394_x13_1_io_result; // @[Math.scala 151:17:@27716.4]
  assign x398_x13_1_io_b = x395_x14_1_io_result; // @[Math.scala 152:17:@27717.4]
  assign x398_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27718.4]
  assign x399_x14_1_clock = clock; // @[:@27724.4]
  assign x399_x14_1_reset = reset; // @[:@27725.4]
  assign x399_x14_1_io_a = x396_x13_1_io_result; // @[Math.scala 151:17:@27726.4]
  assign x399_x14_1_io_b = x397_x14_1_io_result; // @[Math.scala 152:17:@27727.4]
  assign x399_x14_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27728.4]
  assign x400_x13_1_clock = clock; // @[:@27734.4]
  assign x400_x13_1_reset = reset; // @[:@27735.4]
  assign x400_x13_1_io_a = x398_x13_1_io_result; // @[Math.scala 151:17:@27736.4]
  assign x400_x13_1_io_b = x399_x14_1_io_result; // @[Math.scala 152:17:@27737.4]
  assign x400_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27738.4]
  assign RetimeWrapper_68_clock = clock; // @[:@27744.4]
  assign RetimeWrapper_68_reset = reset; // @[:@27745.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27747.4]
  assign RetimeWrapper_68_io_in = x290_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@27746.4]
  assign x401_sum_1_clock = clock; // @[:@27753.4]
  assign x401_sum_1_reset = reset; // @[:@27754.4]
  assign x401_sum_1_io_a = x400_x13_1_io_result; // @[Math.scala 151:17:@27755.4]
  assign x401_sum_1_io_b = RetimeWrapper_68_io_out; // @[Math.scala 152:17:@27756.4]
  assign x401_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27757.4]
  assign x402_1_io_b = x401_sum_1_io_result; // @[Math.scala 721:17:@27765.4]
  assign x403_mul_1_clock = clock; // @[:@27774.4]
  assign x403_mul_1_io_a = x402_1_io_result; // @[Math.scala 263:17:@27776.4]
  assign x403_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@27777.4]
  assign x403_mul_1_io_flow = io_in_x254_TREADY; // @[Math.scala 265:20:@27778.4]
  assign x404_1_io_b = x403_mul_1_io_result; // @[Math.scala 721:17:@27786.4]
  assign RetimeWrapper_69_clock = clock; // @[:@27793.4]
  assign RetimeWrapper_69_reset = reset; // @[:@27794.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27796.4]
  assign RetimeWrapper_69_io_in = x290_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@27795.4]
  assign x405_sub_1_clock = clock; // @[:@27802.4]
  assign x405_sub_1_reset = reset; // @[:@27803.4]
  assign x405_sub_1_io_a = RetimeWrapper_69_io_out; // @[Math.scala 192:17:@27804.4]
  assign x405_sub_1_io_b = x404_1_io_result; // @[Math.scala 193:17:@27805.4]
  assign x405_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@27806.4]
  assign x407_sub_1_clock = clock; // @[:@27817.4]
  assign x407_sub_1_reset = reset; // @[:@27818.4]
  assign x407_sub_1_io_a = x404_1_io_result; // @[Math.scala 192:17:@27819.4]
  assign x407_sub_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 193:17:@27820.4]
  assign x407_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@27821.4]
  assign RetimeWrapper_70_clock = clock; // @[:@27840.4]
  assign RetimeWrapper_70_reset = reset; // @[:@27841.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27843.4]
  assign RetimeWrapper_70_io_in = x409 ? x405_sub_number : 32'h0; // @[package.scala 94:16:@27842.4]
  assign x411_1_io_b = RetimeWrapper_70_io_out; // @[Math.scala 721:17:@27851.4]
  assign x412_mul_1_clock = clock; // @[:@27860.4]
  assign x412_mul_1_io_a = x411_1_io_result; // @[Math.scala 263:17:@27862.4]
  assign x412_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@27863.4]
  assign x412_mul_1_io_flow = io_in_x254_TREADY; // @[Math.scala 265:20:@27864.4]
  assign x413_1_io_b = x412_mul_1_io_result; // @[Math.scala 721:17:@27872.4]
  assign RetimeWrapper_71_clock = clock; // @[:@27879.4]
  assign RetimeWrapper_71_reset = reset; // @[:@27880.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27882.4]
  assign RetimeWrapper_71_io_in = x290_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@27881.4]
  assign x414_sum_1_clock = clock; // @[:@27888.4]
  assign x414_sum_1_reset = reset; // @[:@27889.4]
  assign x414_sum_1_io_a = RetimeWrapper_71_io_out; // @[Math.scala 151:17:@27890.4]
  assign x414_sum_1_io_b = x413_1_io_result; // @[Math.scala 152:17:@27891.4]
  assign x414_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27892.4]
  assign RetimeWrapper_72_clock = clock; // @[:@27900.4]
  assign RetimeWrapper_72_reset = reset; // @[:@27901.4]
  assign RetimeWrapper_72_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27903.4]
  assign RetimeWrapper_72_io_in = _GEN_11 << 1; // @[package.scala 94:16:@27902.4]
  assign RetimeWrapper_73_clock = clock; // @[:@27912.4]
  assign RetimeWrapper_73_reset = reset; // @[:@27913.4]
  assign RetimeWrapper_73_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27915.4]
  assign RetimeWrapper_73_io_in = _GEN_12 << 1; // @[package.scala 94:16:@27914.4]
  assign RetimeWrapper_74_clock = clock; // @[:@27924.4]
  assign RetimeWrapper_74_reset = reset; // @[:@27925.4]
  assign RetimeWrapper_74_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27927.4]
  assign RetimeWrapper_74_io_in = _GEN_13 << 2; // @[package.scala 94:16:@27926.4]
  assign RetimeWrapper_75_clock = clock; // @[:@27936.4]
  assign RetimeWrapper_75_reset = reset; // @[:@27937.4]
  assign RetimeWrapper_75_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27939.4]
  assign RetimeWrapper_75_io_in = _GEN_14 << 1; // @[package.scala 94:16:@27938.4]
  assign RetimeWrapper_76_clock = clock; // @[:@27948.4]
  assign RetimeWrapper_76_reset = reset; // @[:@27949.4]
  assign RetimeWrapper_76_io_flow = io_in_x254_TREADY; // @[package.scala 95:18:@27951.4]
  assign RetimeWrapper_76_io_in = _GEN_15 << 1; // @[package.scala 94:16:@27950.4]
  assign RetimeWrapper_77_clock = clock; // @[:@27958.4]
  assign RetimeWrapper_77_reset = reset; // @[:@27959.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27961.4]
  assign RetimeWrapper_77_io_in = x290_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@27960.4]
  assign x420_x13_1_clock = clock; // @[:@27967.4]
  assign x420_x13_1_reset = reset; // @[:@27968.4]
  assign x420_x13_1_io_a = RetimeWrapper_77_io_out; // @[Math.scala 151:17:@27969.4]
  assign x420_x13_1_io_b = _T_1268[31:0]; // @[Math.scala 152:17:@27970.4]
  assign x420_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27971.4]
  assign RetimeWrapper_78_clock = clock; // @[:@27977.4]
  assign RetimeWrapper_78_reset = reset; // @[:@27978.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27980.4]
  assign RetimeWrapper_78_io_in = x290_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@27979.4]
  assign x421_x14_1_clock = clock; // @[:@27986.4]
  assign x421_x14_1_reset = reset; // @[:@27987.4]
  assign x421_x14_1_io_a = RetimeWrapper_78_io_out; // @[Math.scala 151:17:@27988.4]
  assign x421_x14_1_io_b = _T_1273[31:0]; // @[Math.scala 152:17:@27989.4]
  assign x421_x14_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@27990.4]
  assign x422_x13_1_clock = clock; // @[:@27996.4]
  assign x422_x13_1_reset = reset; // @[:@27997.4]
  assign x422_x13_1_io_a = _T_1278[31:0]; // @[Math.scala 151:17:@27998.4]
  assign x422_x13_1_io_b = _T_1283[31:0]; // @[Math.scala 152:17:@27999.4]
  assign x422_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28000.4]
  assign RetimeWrapper_79_clock = clock; // @[:@28006.4]
  assign RetimeWrapper_79_reset = reset; // @[:@28007.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28009.4]
  assign RetimeWrapper_79_io_in = x290_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@28008.4]
  assign x423_x14_1_clock = clock; // @[:@28017.4]
  assign x423_x14_1_reset = reset; // @[:@28018.4]
  assign x423_x14_1_io_a = RetimeWrapper_79_io_out; // @[Math.scala 151:17:@28019.4]
  assign x423_x14_1_io_b = _T_1288[31:0]; // @[Math.scala 152:17:@28020.4]
  assign x423_x14_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28021.4]
  assign x424_x13_1_clock = clock; // @[:@28027.4]
  assign x424_x13_1_reset = reset; // @[:@28028.4]
  assign x424_x13_1_io_a = x420_x13_1_io_result; // @[Math.scala 151:17:@28029.4]
  assign x424_x13_1_io_b = x421_x14_1_io_result; // @[Math.scala 152:17:@28030.4]
  assign x424_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28031.4]
  assign x425_x14_1_clock = clock; // @[:@28037.4]
  assign x425_x14_1_reset = reset; // @[:@28038.4]
  assign x425_x14_1_io_a = x422_x13_1_io_result; // @[Math.scala 151:17:@28039.4]
  assign x425_x14_1_io_b = x423_x14_1_io_result; // @[Math.scala 152:17:@28040.4]
  assign x425_x14_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28041.4]
  assign x426_x13_1_clock = clock; // @[:@28047.4]
  assign x426_x13_1_reset = reset; // @[:@28048.4]
  assign x426_x13_1_io_a = x424_x13_1_io_result; // @[Math.scala 151:17:@28049.4]
  assign x426_x13_1_io_b = x425_x14_1_io_result; // @[Math.scala 152:17:@28050.4]
  assign x426_x13_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28051.4]
  assign RetimeWrapper_80_clock = clock; // @[:@28057.4]
  assign RetimeWrapper_80_reset = reset; // @[:@28058.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28060.4]
  assign RetimeWrapper_80_io_in = x290_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@28059.4]
  assign x427_sum_1_clock = clock; // @[:@28066.4]
  assign x427_sum_1_reset = reset; // @[:@28067.4]
  assign x427_sum_1_io_a = x426_x13_1_io_result; // @[Math.scala 151:17:@28068.4]
  assign x427_sum_1_io_b = RetimeWrapper_80_io_out; // @[Math.scala 152:17:@28069.4]
  assign x427_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28070.4]
  assign x428_1_io_b = x427_sum_1_io_result; // @[Math.scala 721:17:@28078.4]
  assign x429_mul_1_clock = clock; // @[:@28087.4]
  assign x429_mul_1_io_a = x428_1_io_result; // @[Math.scala 263:17:@28089.4]
  assign x429_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@28090.4]
  assign x429_mul_1_io_flow = io_in_x254_TREADY; // @[Math.scala 265:20:@28091.4]
  assign x430_1_io_b = x429_mul_1_io_result; // @[Math.scala 721:17:@28099.4]
  assign RetimeWrapper_81_clock = clock; // @[:@28106.4]
  assign RetimeWrapper_81_reset = reset; // @[:@28107.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28109.4]
  assign RetimeWrapper_81_io_in = x290_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@28108.4]
  assign x431_sub_1_clock = clock; // @[:@28115.4]
  assign x431_sub_1_reset = reset; // @[:@28116.4]
  assign x431_sub_1_io_a = RetimeWrapper_81_io_out; // @[Math.scala 192:17:@28117.4]
  assign x431_sub_1_io_b = x430_1_io_result; // @[Math.scala 193:17:@28118.4]
  assign x431_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@28119.4]
  assign x433_sub_1_clock = clock; // @[:@28130.4]
  assign x433_sub_1_reset = reset; // @[:@28131.4]
  assign x433_sub_1_io_a = x430_1_io_result; // @[Math.scala 192:17:@28132.4]
  assign x433_sub_1_io_b = RetimeWrapper_81_io_out; // @[Math.scala 193:17:@28133.4]
  assign x433_sub_1_io_flow = io_in_x254_TREADY; // @[Math.scala 194:20:@28134.4]
  assign RetimeWrapper_82_clock = clock; // @[:@28153.4]
  assign RetimeWrapper_82_reset = reset; // @[:@28154.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28156.4]
  assign RetimeWrapper_82_io_in = x435 ? x431_sub_number : 32'h0; // @[package.scala 94:16:@28155.4]
  assign x437_1_io_b = RetimeWrapper_82_io_out; // @[Math.scala 721:17:@28164.4]
  assign x438_mul_1_clock = clock; // @[:@28173.4]
  assign x438_mul_1_io_a = x437_1_io_result; // @[Math.scala 263:17:@28175.4]
  assign x438_mul_1_io_b = 32'h20; // @[Math.scala 264:17:@28176.4]
  assign x438_mul_1_io_flow = io_in_x254_TREADY; // @[Math.scala 265:20:@28177.4]
  assign x439_1_io_b = x438_mul_1_io_result; // @[Math.scala 721:17:@28185.4]
  assign RetimeWrapper_83_clock = clock; // @[:@28192.4]
  assign RetimeWrapper_83_reset = reset; // @[:@28193.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28195.4]
  assign RetimeWrapper_83_io_in = x290_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@28194.4]
  assign x440_sum_1_clock = clock; // @[:@28201.4]
  assign x440_sum_1_reset = reset; // @[:@28202.4]
  assign x440_sum_1_io_a = RetimeWrapper_83_io_out; // @[Math.scala 151:17:@28203.4]
  assign x440_sum_1_io_b = x439_1_io_result; // @[Math.scala 152:17:@28204.4]
  assign x440_sum_1_io_flow = io_in_x254_TREADY; // @[Math.scala 153:20:@28205.4]
  assign RetimeWrapper_84_clock = clock; // @[:@28217.4]
  assign RetimeWrapper_84_reset = reset; // @[:@28218.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28220.4]
  assign RetimeWrapper_84_io_in = {x414_sum_number,x440_sum_number}; // @[package.scala 94:16:@28219.4]
  assign RetimeWrapper_85_clock = clock; // @[:@28226.4]
  assign RetimeWrapper_85_reset = reset; // @[:@28227.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28229.4]
  assign RetimeWrapper_85_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@28228.4]
  assign RetimeWrapper_86_clock = clock; // @[:@28235.4]
  assign RetimeWrapper_86_reset = reset; // @[:@28236.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28238.4]
  assign RetimeWrapper_86_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@28237.4]
  assign RetimeWrapper_87_clock = clock; // @[:@28244.4]
  assign RetimeWrapper_87_reset = reset; // @[:@28245.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28247.4]
  assign RetimeWrapper_87_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28246.4]
endmodule
module x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1( // @[:@28265.2]
  input          clock, // @[:@28266.4]
  input          reset, // @[:@28267.4]
  input          io_in_x253_TVALID, // @[:@28268.4]
  output         io_in_x253_TREADY, // @[:@28268.4]
  input  [255:0] io_in_x253_TDATA, // @[:@28268.4]
  input  [7:0]   io_in_x253_TID, // @[:@28268.4]
  input  [7:0]   io_in_x253_TDEST, // @[:@28268.4]
  output         io_in_x254_TVALID, // @[:@28268.4]
  input          io_in_x254_TREADY, // @[:@28268.4]
  output [255:0] io_in_x254_TDATA, // @[:@28268.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@28268.4]
  input          io_sigsIn_smChildAcks_0, // @[:@28268.4]
  output         io_sigsOut_smDoneIn_0, // @[:@28268.4]
  input          io_rr // @[:@28268.4]
);
  wire  x283_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x283_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x283_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x283_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire [12:0] x283_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire [12:0] x283_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x283_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x283_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x283_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@28302.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@28390.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@28390.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@28390.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@28390.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@28390.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@28432.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@28432.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@28432.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@28432.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@28432.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@28440.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@28440.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@28440.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@28440.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@28440.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TREADY; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire [255:0] x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TDATA; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire [7:0] x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TID; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire [7:0] x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TDEST; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TVALID; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TREADY; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire [255:0] x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TDATA; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire [31:0] x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire [31:0] x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
  wire  _T_240; // @[package.scala 96:25:@28395.4 package.scala 96:25:@28396.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x446_outr_UnitPipe.scala 69:66:@28401.4]
  wire  _T_253; // @[package.scala 96:25:@28437.4 package.scala 96:25:@28438.4]
  wire  _T_259; // @[package.scala 96:25:@28445.4 package.scala 96:25:@28446.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@28448.4]
  wire  x445_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@28449.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@28457.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@28458.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@28470.4]
  x261_ctrchain x283_ctrchain ( // @[SpatialBlocks.scala 37:22:@28302.4]
    .clock(x283_ctrchain_clock),
    .reset(x283_ctrchain_reset),
    .io_input_reset(x283_ctrchain_io_input_reset),
    .io_input_enable(x283_ctrchain_io_input_enable),
    .io_output_counts_1(x283_ctrchain_io_output_counts_1),
    .io_output_counts_0(x283_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x283_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x283_ctrchain_io_output_oobs_1),
    .io_output_done(x283_ctrchain_io_output_done)
  );
  x445_inr_Foreach_SAMPLER_BOX_sm x445_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 32:18:@28362.4]
    .clock(x445_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x445_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x445_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x445_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x445_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x445_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x445_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x445_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x445_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@28390.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@28432.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@28440.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1 x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 602:24:@28474.4]
    .clock(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x253_TREADY(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TREADY),
    .io_in_x253_TDATA(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TDATA),
    .io_in_x253_TID(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TID),
    .io_in_x253_TDEST(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TDEST),
    .io_in_x254_TVALID(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TVALID),
    .io_in_x254_TREADY(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TREADY),
    .io_in_x254_TDATA(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TDATA),
    .io_sigsIn_backpressure(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@28395.4 package.scala 96:25:@28396.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x253_TVALID | x445_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x446_outr_UnitPipe.scala 69:66:@28401.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@28437.4 package.scala 96:25:@28438.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@28445.4 package.scala 96:25:@28446.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@28448.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@28449.4]
  assign _T_264 = x445_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@28457.4]
  assign _T_265 = ~ x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@28458.4]
  assign _T_272 = x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@28470.4]
  assign io_in_x253_TREADY = x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TREADY; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 48:23:@28532.4]
  assign io_in_x254_TVALID = x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TVALID; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 49:23:@28542.4]
  assign io_in_x254_TDATA = x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TDATA; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 49:23:@28540.4]
  assign io_sigsOut_smDoneIn_0 = x445_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@28455.4]
  assign x283_ctrchain_clock = clock; // @[:@28303.4]
  assign x283_ctrchain_reset = reset; // @[:@28304.4]
  assign x283_ctrchain_io_input_reset = x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@28473.4]
  assign x283_ctrchain_io_input_enable = _T_272 & x445_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@28425.4 SpatialBlocks.scala 159:42:@28472.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@28363.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@28364.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_io_enable = x445_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x445_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@28452.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x446_outr_UnitPipe.scala 67:50:@28398.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@28454.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x254_TREADY | x445_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@28426.4]
  assign x445_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x446_outr_UnitPipe.scala 71:48:@28404.4]
  assign RetimeWrapper_clock = clock; // @[:@28391.4]
  assign RetimeWrapper_reset = reset; // @[:@28392.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@28394.4]
  assign RetimeWrapper_io_in = x283_ctrchain_io_output_done; // @[package.scala 94:16:@28393.4]
  assign RetimeWrapper_1_clock = clock; // @[:@28433.4]
  assign RetimeWrapper_1_reset = reset; // @[:@28434.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@28436.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@28435.4]
  assign RetimeWrapper_2_clock = clock; // @[:@28441.4]
  assign RetimeWrapper_2_reset = reset; // @[:@28442.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@28444.4]
  assign RetimeWrapper_2_io_in = x445_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@28443.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@28475.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@28476.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TDATA = io_in_x253_TDATA; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 48:23:@28531.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TID = io_in_x253_TID; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 48:23:@28527.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x253_TDEST = io_in_x253_TDEST; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 48:23:@28526.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x254_TREADY = io_in_x254_TREADY; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 49:23:@28541.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x254_TREADY | x445_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28559.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28557.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x445_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28555.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x283_ctrchain_io_output_counts_1[12]}},x283_ctrchain_io_output_counts_1}; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28550.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x283_ctrchain_io_output_counts_0[12]}},x283_ctrchain_io_output_counts_0}; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28549.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x283_ctrchain_io_output_oobs_0; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28547.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x283_ctrchain_io_output_oobs_1; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 607:22:@28548.4]
  assign x445_inr_Foreach_SAMPLER_BOX_kernelx445_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x445_inr_Foreach_SAMPLER_BOX.scala 606:18:@28543.4]
endmodule
module x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1( // @[:@28573.2]
  input          clock, // @[:@28574.4]
  input          reset, // @[:@28575.4]
  input          io_in_x253_TVALID, // @[:@28576.4]
  output         io_in_x253_TREADY, // @[:@28576.4]
  input  [255:0] io_in_x253_TDATA, // @[:@28576.4]
  input  [7:0]   io_in_x253_TID, // @[:@28576.4]
  input  [7:0]   io_in_x253_TDEST, // @[:@28576.4]
  output         io_in_x254_TVALID, // @[:@28576.4]
  input          io_in_x254_TREADY, // @[:@28576.4]
  output [255:0] io_in_x254_TDATA, // @[:@28576.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@28576.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@28576.4]
  input          io_sigsIn_smChildAcks_0, // @[:@28576.4]
  input          io_sigsIn_smChildAcks_1, // @[:@28576.4]
  output         io_sigsOut_smDoneIn_0, // @[:@28576.4]
  output         io_sigsOut_smDoneIn_1, // @[:@28576.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@28576.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@28576.4]
  input          io_rr // @[:@28576.4]
);
  wire  x256_fifoinraw_0_clock; // @[m_x256_fifoinraw_0.scala 27:17:@28590.4]
  wire  x256_fifoinraw_0_reset; // @[m_x256_fifoinraw_0.scala 27:17:@28590.4]
  wire  x257_fifoinpacked_0_clock; // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
  wire  x257_fifoinpacked_0_reset; // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
  wire  x257_fifoinpacked_0_io_wPort_0_en_0; // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
  wire  x257_fifoinpacked_0_io_full; // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
  wire  x257_fifoinpacked_0_io_active_0_in; // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
  wire  x257_fifoinpacked_0_io_active_0_out; // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
  wire  x258_fifooutraw_0_clock; // @[m_x258_fifooutraw_0.scala 27:17:@28638.4]
  wire  x258_fifooutraw_0_reset; // @[m_x258_fifooutraw_0.scala 27:17:@28638.4]
  wire  x261_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x261_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x261_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x261_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire [12:0] x261_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire [12:0] x261_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x261_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x261_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x261_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@28662.4]
  wire  x279_inr_Foreach_sm_clock; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_reset; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_enable; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_done; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_doneLatch; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_ctrDone; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_datapathEn; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_ctrInc; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_ctrRst; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_parentAck; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_backpressure; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  x279_inr_Foreach_sm_io_break; // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@28750.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@28750.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@28750.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@28750.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@28750.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@28796.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@28796.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@28796.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@28796.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@28796.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@28804.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@28804.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@28804.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@28804.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@28804.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_clock; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_reset; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_wPort_0_en_0; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_full; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_active_0_in; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_active_0_out; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire [31:0] x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire [31:0] x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_rr; // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
  wire  x446_outr_UnitPipe_sm_clock; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_reset; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_enable; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_done; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_rst; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_ctrDone; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_ctrInc; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_parentAck; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  x446_outr_UnitPipe_sm_io_childAck_0; // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@29036.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@29036.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@29036.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@29036.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@29036.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_clock; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_reset; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TVALID; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TREADY; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire [255:0] x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TDATA; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire [7:0] x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TID; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire [7:0] x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TDEST; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TVALID; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TREADY; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire [255:0] x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TDATA; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_rr; // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
  wire  _T_254; // @[package.scala 96:25:@28755.4 package.scala 96:25:@28756.4]
  wire  _T_260; // @[implicits.scala 47:10:@28759.4]
  wire  _T_261; // @[sm_x447_outr_UnitPipe.scala 70:41:@28760.4]
  wire  _T_262; // @[sm_x447_outr_UnitPipe.scala 70:78:@28761.4]
  wire  _T_263; // @[sm_x447_outr_UnitPipe.scala 70:76:@28762.4]
  wire  _T_275; // @[package.scala 96:25:@28801.4 package.scala 96:25:@28802.4]
  wire  _T_281; // @[package.scala 96:25:@28809.4 package.scala 96:25:@28810.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@28812.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@28821.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@28822.4]
  wire  _T_354; // @[package.scala 100:49:@28999.4]
  reg  _T_357; // @[package.scala 48:56:@29000.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@29033.4 package.scala 96:25:@29034.4]
  wire  _T_377; // @[package.scala 96:25:@29041.4 package.scala 96:25:@29042.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@29044.4]
  x256_fifoinraw_0 x256_fifoinraw_0 ( // @[m_x256_fifoinraw_0.scala 27:17:@28590.4]
    .clock(x256_fifoinraw_0_clock),
    .reset(x256_fifoinraw_0_reset)
  );
  x257_fifoinpacked_0 x257_fifoinpacked_0 ( // @[m_x257_fifoinpacked_0.scala 27:17:@28614.4]
    .clock(x257_fifoinpacked_0_clock),
    .reset(x257_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x257_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x257_fifoinpacked_0_io_full),
    .io_active_0_in(x257_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x257_fifoinpacked_0_io_active_0_out)
  );
  x256_fifoinraw_0 x258_fifooutraw_0 ( // @[m_x258_fifooutraw_0.scala 27:17:@28638.4]
    .clock(x258_fifooutraw_0_clock),
    .reset(x258_fifooutraw_0_reset)
  );
  x261_ctrchain x261_ctrchain ( // @[SpatialBlocks.scala 37:22:@28662.4]
    .clock(x261_ctrchain_clock),
    .reset(x261_ctrchain_reset),
    .io_input_reset(x261_ctrchain_io_input_reset),
    .io_input_enable(x261_ctrchain_io_input_enable),
    .io_output_counts_1(x261_ctrchain_io_output_counts_1),
    .io_output_counts_0(x261_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x261_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x261_ctrchain_io_output_oobs_1),
    .io_output_done(x261_ctrchain_io_output_done)
  );
  x279_inr_Foreach_sm x279_inr_Foreach_sm ( // @[sm_x279_inr_Foreach.scala 32:18:@28722.4]
    .clock(x279_inr_Foreach_sm_clock),
    .reset(x279_inr_Foreach_sm_reset),
    .io_enable(x279_inr_Foreach_sm_io_enable),
    .io_done(x279_inr_Foreach_sm_io_done),
    .io_doneLatch(x279_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x279_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x279_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x279_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x279_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x279_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x279_inr_Foreach_sm_io_backpressure),
    .io_break(x279_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@28750.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@28796.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@28804.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x279_inr_Foreach_kernelx279_inr_Foreach_concrete1 x279_inr_Foreach_kernelx279_inr_Foreach_concrete1 ( // @[sm_x279_inr_Foreach.scala 106:24:@28839.4]
    .clock(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_clock),
    .reset(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_reset),
    .io_in_x257_fifoinpacked_0_wPort_0_en_0(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_wPort_0_en_0),
    .io_in_x257_fifoinpacked_0_full(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_full),
    .io_in_x257_fifoinpacked_0_active_0_in(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_active_0_in),
    .io_in_x257_fifoinpacked_0_active_0_out(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x446_outr_UnitPipe_sm ( // @[sm_x446_outr_UnitPipe.scala 32:18:@28971.4]
    .clock(x446_outr_UnitPipe_sm_clock),
    .reset(x446_outr_UnitPipe_sm_reset),
    .io_enable(x446_outr_UnitPipe_sm_io_enable),
    .io_done(x446_outr_UnitPipe_sm_io_done),
    .io_rst(x446_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x446_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x446_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x446_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x446_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x446_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x446_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@29028.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@29036.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1 x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1 ( // @[sm_x446_outr_UnitPipe.scala 76:24:@29066.4]
    .clock(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_clock),
    .reset(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_reset),
    .io_in_x253_TVALID(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TVALID),
    .io_in_x253_TREADY(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TREADY),
    .io_in_x253_TDATA(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TDATA),
    .io_in_x253_TID(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TID),
    .io_in_x253_TDEST(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TDEST),
    .io_in_x254_TVALID(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TVALID),
    .io_in_x254_TREADY(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TREADY),
    .io_in_x254_TDATA(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TDATA),
    .io_sigsIn_smEnableOuts_0(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@28755.4 package.scala 96:25:@28756.4]
  assign _T_260 = x257_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@28759.4]
  assign _T_261 = ~ _T_260; // @[sm_x447_outr_UnitPipe.scala 70:41:@28760.4]
  assign _T_262 = ~ x257_fifoinpacked_0_io_active_0_out; // @[sm_x447_outr_UnitPipe.scala 70:78:@28761.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x447_outr_UnitPipe.scala 70:76:@28762.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@28801.4 package.scala 96:25:@28802.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@28809.4 package.scala 96:25:@28810.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@28812.4]
  assign _T_286 = x279_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@28821.4]
  assign _T_287 = ~ x279_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@28822.4]
  assign _T_354 = x446_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@28999.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@29033.4 package.scala 96:25:@29034.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@29041.4 package.scala 96:25:@29042.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@29044.4]
  assign io_in_x253_TREADY = x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TREADY; // @[sm_x446_outr_UnitPipe.scala 48:23:@29122.4]
  assign io_in_x254_TVALID = x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TVALID; // @[sm_x446_outr_UnitPipe.scala 49:23:@29132.4]
  assign io_in_x254_TDATA = x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TDATA; // @[sm_x446_outr_UnitPipe.scala 49:23:@29130.4]
  assign io_sigsOut_smDoneIn_0 = x279_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@28819.4]
  assign io_sigsOut_smDoneIn_1 = x446_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@29051.4]
  assign io_sigsOut_smCtrCopyDone_0 = x279_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@28838.4]
  assign io_sigsOut_smCtrCopyDone_1 = x446_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@29065.4]
  assign x256_fifoinraw_0_clock = clock; // @[:@28591.4]
  assign x256_fifoinraw_0_reset = reset; // @[:@28592.4]
  assign x257_fifoinpacked_0_clock = clock; // @[:@28615.4]
  assign x257_fifoinpacked_0_reset = reset; // @[:@28616.4]
  assign x257_fifoinpacked_0_io_wPort_0_en_0 = x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@28899.4]
  assign x257_fifoinpacked_0_io_active_0_in = x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@28898.4]
  assign x258_fifooutraw_0_clock = clock; // @[:@28639.4]
  assign x258_fifooutraw_0_reset = reset; // @[:@28640.4]
  assign x261_ctrchain_clock = clock; // @[:@28663.4]
  assign x261_ctrchain_reset = reset; // @[:@28664.4]
  assign x261_ctrchain_io_input_reset = x279_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@28837.4]
  assign x261_ctrchain_io_input_enable = x279_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@28789.4 SpatialBlocks.scala 159:42:@28836.4]
  assign x279_inr_Foreach_sm_clock = clock; // @[:@28723.4]
  assign x279_inr_Foreach_sm_reset = reset; // @[:@28724.4]
  assign x279_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@28816.4]
  assign x279_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x447_outr_UnitPipe.scala 69:38:@28758.4]
  assign x279_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@28818.4]
  assign x279_inr_Foreach_sm_io_backpressure = _T_263 | x279_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@28790.4]
  assign x279_inr_Foreach_sm_io_break = 1'h0; // @[sm_x447_outr_UnitPipe.scala 73:36:@28768.4]
  assign RetimeWrapper_clock = clock; // @[:@28751.4]
  assign RetimeWrapper_reset = reset; // @[:@28752.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@28754.4]
  assign RetimeWrapper_io_in = x261_ctrchain_io_output_done; // @[package.scala 94:16:@28753.4]
  assign RetimeWrapper_1_clock = clock; // @[:@28797.4]
  assign RetimeWrapper_1_reset = reset; // @[:@28798.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@28800.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@28799.4]
  assign RetimeWrapper_2_clock = clock; // @[:@28805.4]
  assign RetimeWrapper_2_reset = reset; // @[:@28806.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@28808.4]
  assign RetimeWrapper_2_io_in = x279_inr_Foreach_sm_io_done; // @[package.scala 94:16:@28807.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_clock = clock; // @[:@28840.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_reset = reset; // @[:@28841.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_full = x257_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@28893.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_in_x257_fifoinpacked_0_active_0_out = x257_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@28892.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x279_inr_Foreach_sm_io_doneLatch; // @[sm_x279_inr_Foreach.scala 111:22:@28922.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x279_inr_Foreach.scala 111:22:@28920.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_break = x279_inr_Foreach_sm_io_break; // @[sm_x279_inr_Foreach.scala 111:22:@28918.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x261_ctrchain_io_output_counts_1[12]}},x261_ctrchain_io_output_counts_1}; // @[sm_x279_inr_Foreach.scala 111:22:@28913.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x261_ctrchain_io_output_counts_0[12]}},x261_ctrchain_io_output_counts_0}; // @[sm_x279_inr_Foreach.scala 111:22:@28912.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x261_ctrchain_io_output_oobs_0; // @[sm_x279_inr_Foreach.scala 111:22:@28910.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x261_ctrchain_io_output_oobs_1; // @[sm_x279_inr_Foreach.scala 111:22:@28911.4]
  assign x279_inr_Foreach_kernelx279_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x279_inr_Foreach.scala 110:18:@28906.4]
  assign x446_outr_UnitPipe_sm_clock = clock; // @[:@28972.4]
  assign x446_outr_UnitPipe_sm_reset = reset; // @[:@28973.4]
  assign x446_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@29048.4]
  assign x446_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@29023.4]
  assign x446_outr_UnitPipe_sm_io_ctrDone = x446_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x447_outr_UnitPipe.scala 78:40:@29003.4]
  assign x446_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@29050.4]
  assign x446_outr_UnitPipe_sm_io_doneIn_0 = x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@29020.4]
  assign RetimeWrapper_3_clock = clock; // @[:@29029.4]
  assign RetimeWrapper_3_reset = reset; // @[:@29030.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@29032.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@29031.4]
  assign RetimeWrapper_4_clock = clock; // @[:@29037.4]
  assign RetimeWrapper_4_reset = reset; // @[:@29038.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@29040.4]
  assign RetimeWrapper_4_io_in = x446_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@29039.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_clock = clock; // @[:@29067.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_reset = reset; // @[:@29068.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TVALID = io_in_x253_TVALID; // @[sm_x446_outr_UnitPipe.scala 48:23:@29123.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TDATA = io_in_x253_TDATA; // @[sm_x446_outr_UnitPipe.scala 48:23:@29121.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TID = io_in_x253_TID; // @[sm_x446_outr_UnitPipe.scala 48:23:@29117.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x253_TDEST = io_in_x253_TDEST; // @[sm_x446_outr_UnitPipe.scala 48:23:@29116.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_in_x254_TREADY = io_in_x254_TREADY; // @[sm_x446_outr_UnitPipe.scala 49:23:@29131.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x446_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x446_outr_UnitPipe.scala 81:22:@29141.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x446_outr_UnitPipe_sm_io_childAck_0; // @[sm_x446_outr_UnitPipe.scala 81:22:@29139.4]
  assign x446_outr_UnitPipe_kernelx446_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x446_outr_UnitPipe.scala 80:18:@29133.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x469_outr_UnitPipe_sm( // @[:@29630.2]
  input   clock, // @[:@29631.4]
  input   reset, // @[:@29632.4]
  input   io_enable, // @[:@29633.4]
  output  io_done, // @[:@29633.4]
  input   io_parentAck, // @[:@29633.4]
  input   io_doneIn_0, // @[:@29633.4]
  input   io_doneIn_1, // @[:@29633.4]
  input   io_doneIn_2, // @[:@29633.4]
  output  io_enableOut_0, // @[:@29633.4]
  output  io_enableOut_1, // @[:@29633.4]
  output  io_enableOut_2, // @[:@29633.4]
  output  io_childAck_0, // @[:@29633.4]
  output  io_childAck_1, // @[:@29633.4]
  output  io_childAck_2, // @[:@29633.4]
  input   io_ctrCopyDone_0, // @[:@29633.4]
  input   io_ctrCopyDone_1, // @[:@29633.4]
  input   io_ctrCopyDone_2 // @[:@29633.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@29636.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@29636.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@29636.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@29636.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@29636.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@29636.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@29639.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@29639.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@29639.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@29639.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@29639.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@29639.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@29642.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@29642.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@29642.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@29642.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@29642.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@29642.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@29645.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@29645.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@29645.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@29645.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@29645.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@29645.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@29648.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@29648.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@29648.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@29648.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@29648.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@29648.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@29651.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@29651.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@29651.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@29651.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@29651.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@29651.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@29692.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@29692.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@29692.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@29692.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@29692.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@29692.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@29695.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@29695.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@29695.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@29695.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@29695.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@29695.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@29698.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@29698.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@29698.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@29698.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@29698.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@29698.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29749.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29749.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29749.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29749.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29749.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29763.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29763.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29763.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29763.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29763.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29781.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29781.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29781.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29781.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29781.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@29818.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@29818.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@29818.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@29818.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@29818.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@29832.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@29832.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@29832.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@29832.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@29832.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@29850.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@29850.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@29850.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@29850.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@29850.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@29887.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@29887.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@29887.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@29887.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@29887.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@29901.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@29901.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@29901.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@29901.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@29901.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@29976.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@29976.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@29976.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@29976.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@29976.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@29993.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@29993.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@29993.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@29993.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@29993.4]
  wire  _T_77; // @[Controllers.scala 80:47:@29654.4]
  wire  allDone; // @[Controllers.scala 80:47:@29655.4]
  wire  _T_151; // @[Controllers.scala 165:35:@29733.4]
  wire  _T_153; // @[Controllers.scala 165:60:@29734.4]
  wire  _T_154; // @[Controllers.scala 165:58:@29735.4]
  wire  _T_156; // @[Controllers.scala 165:76:@29736.4]
  wire  _T_157; // @[Controllers.scala 165:74:@29737.4]
  wire  _T_161; // @[Controllers.scala 165:109:@29740.4]
  wire  _T_164; // @[Controllers.scala 165:141:@29742.4]
  wire  _T_172; // @[package.scala 96:25:@29754.4 package.scala 96:25:@29755.4]
  wire  _T_176; // @[Controllers.scala 167:54:@29757.4]
  wire  _T_177; // @[Controllers.scala 167:52:@29758.4]
  wire  _T_184; // @[package.scala 96:25:@29768.4 package.scala 96:25:@29769.4]
  wire  _T_202; // @[package.scala 96:25:@29786.4 package.scala 96:25:@29787.4]
  wire  _T_206; // @[Controllers.scala 169:67:@29789.4]
  wire  _T_207; // @[Controllers.scala 169:86:@29790.4]
  wire  _T_219; // @[Controllers.scala 165:35:@29802.4]
  wire  _T_221; // @[Controllers.scala 165:60:@29803.4]
  wire  _T_222; // @[Controllers.scala 165:58:@29804.4]
  wire  _T_224; // @[Controllers.scala 165:76:@29805.4]
  wire  _T_225; // @[Controllers.scala 165:74:@29806.4]
  wire  _T_229; // @[Controllers.scala 165:109:@29809.4]
  wire  _T_232; // @[Controllers.scala 165:141:@29811.4]
  wire  _T_240; // @[package.scala 96:25:@29823.4 package.scala 96:25:@29824.4]
  wire  _T_244; // @[Controllers.scala 167:54:@29826.4]
  wire  _T_245; // @[Controllers.scala 167:52:@29827.4]
  wire  _T_252; // @[package.scala 96:25:@29837.4 package.scala 96:25:@29838.4]
  wire  _T_270; // @[package.scala 96:25:@29855.4 package.scala 96:25:@29856.4]
  wire  _T_274; // @[Controllers.scala 169:67:@29858.4]
  wire  _T_275; // @[Controllers.scala 169:86:@29859.4]
  wire  _T_287; // @[Controllers.scala 165:35:@29871.4]
  wire  _T_289; // @[Controllers.scala 165:60:@29872.4]
  wire  _T_290; // @[Controllers.scala 165:58:@29873.4]
  wire  _T_292; // @[Controllers.scala 165:76:@29874.4]
  wire  _T_293; // @[Controllers.scala 165:74:@29875.4]
  wire  _T_297; // @[Controllers.scala 165:109:@29878.4]
  wire  _T_300; // @[Controllers.scala 165:141:@29880.4]
  wire  _T_308; // @[package.scala 96:25:@29892.4 package.scala 96:25:@29893.4]
  wire  _T_312; // @[Controllers.scala 167:54:@29895.4]
  wire  _T_313; // @[Controllers.scala 167:52:@29896.4]
  wire  _T_320; // @[package.scala 96:25:@29906.4 package.scala 96:25:@29907.4]
  wire  _T_338; // @[package.scala 96:25:@29924.4 package.scala 96:25:@29925.4]
  wire  _T_342; // @[Controllers.scala 169:67:@29927.4]
  wire  _T_343; // @[Controllers.scala 169:86:@29928.4]
  wire  _T_358; // @[Controllers.scala 213:68:@29946.4]
  wire  _T_360; // @[Controllers.scala 213:90:@29948.4]
  wire  _T_362; // @[Controllers.scala 213:132:@29950.4]
  wire  _T_366; // @[Controllers.scala 213:68:@29955.4]
  wire  _T_368; // @[Controllers.scala 213:90:@29957.4]
  wire  _T_374; // @[Controllers.scala 213:68:@29963.4]
  wire  _T_376; // @[Controllers.scala 213:90:@29965.4]
  wire  _T_383; // @[package.scala 100:49:@29971.4]
  reg  _T_386; // @[package.scala 48:56:@29972.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@29974.4]
  reg  _T_400; // @[package.scala 48:56:@29990.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@29636.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@29639.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@29642.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@29645.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@29648.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@29651.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@29692.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@29695.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@29698.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29749.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29763.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29781.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@29818.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@29832.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@29850.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@29887.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@29901.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@29919.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@29976.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@29993.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@29654.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@29655.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@29733.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@29734.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@29735.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@29736.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@29737.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@29740.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@29742.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@29754.4 package.scala 96:25:@29755.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@29757.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@29758.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29768.4 package.scala 96:25:@29769.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29786.4 package.scala 96:25:@29787.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@29789.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@29790.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@29802.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@29803.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@29804.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@29805.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@29806.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@29809.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@29811.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@29823.4 package.scala 96:25:@29824.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@29826.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@29827.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@29837.4 package.scala 96:25:@29838.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@29855.4 package.scala 96:25:@29856.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@29858.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@29859.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@29871.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@29872.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@29873.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@29874.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@29875.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@29878.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@29880.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@29892.4 package.scala 96:25:@29893.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@29895.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@29896.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@29906.4 package.scala 96:25:@29907.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@29924.4 package.scala 96:25:@29925.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@29927.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@29928.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@29946.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@29948.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@29950.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@29955.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@29957.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@29963.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@29965.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@29971.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@29974.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@30000.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@29954.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@29962.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@29970.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@29941.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@29943.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@29945.4]
  assign active_0_clock = clock; // @[:@29637.4]
  assign active_0_reset = reset; // @[:@29638.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@29744.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@29748.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@29658.4]
  assign active_1_clock = clock; // @[:@29640.4]
  assign active_1_reset = reset; // @[:@29641.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@29813.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@29817.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@29659.4]
  assign active_2_clock = clock; // @[:@29643.4]
  assign active_2_reset = reset; // @[:@29644.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@29882.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@29886.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@29660.4]
  assign done_0_clock = clock; // @[:@29646.4]
  assign done_0_reset = reset; // @[:@29647.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@29794.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@29672.4 Controllers.scala 170:32:@29801.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@29661.4]
  assign done_1_clock = clock; // @[:@29649.4]
  assign done_1_reset = reset; // @[:@29650.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@29863.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@29681.4 Controllers.scala 170:32:@29870.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@29662.4]
  assign done_2_clock = clock; // @[:@29652.4]
  assign done_2_reset = reset; // @[:@29653.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@29932.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@29690.4 Controllers.scala 170:32:@29939.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@29663.4]
  assign iterDone_0_clock = clock; // @[:@29693.4]
  assign iterDone_0_reset = reset; // @[:@29694.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@29762.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@29712.4 Controllers.scala 168:36:@29778.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@29701.4]
  assign iterDone_1_clock = clock; // @[:@29696.4]
  assign iterDone_1_reset = reset; // @[:@29697.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@29831.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@29721.4 Controllers.scala 168:36:@29847.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@29702.4]
  assign iterDone_2_clock = clock; // @[:@29699.4]
  assign iterDone_2_reset = reset; // @[:@29700.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@29900.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@29730.4 Controllers.scala 168:36:@29916.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@29703.4]
  assign RetimeWrapper_clock = clock; // @[:@29750.4]
  assign RetimeWrapper_reset = reset; // @[:@29751.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29753.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@29752.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29764.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29765.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29767.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@29766.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29782.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29783.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29785.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@29784.4]
  assign RetimeWrapper_3_clock = clock; // @[:@29819.4]
  assign RetimeWrapper_3_reset = reset; // @[:@29820.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@29822.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@29821.4]
  assign RetimeWrapper_4_clock = clock; // @[:@29833.4]
  assign RetimeWrapper_4_reset = reset; // @[:@29834.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@29836.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@29835.4]
  assign RetimeWrapper_5_clock = clock; // @[:@29851.4]
  assign RetimeWrapper_5_reset = reset; // @[:@29852.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@29854.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@29853.4]
  assign RetimeWrapper_6_clock = clock; // @[:@29888.4]
  assign RetimeWrapper_6_reset = reset; // @[:@29889.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@29891.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@29890.4]
  assign RetimeWrapper_7_clock = clock; // @[:@29902.4]
  assign RetimeWrapper_7_reset = reset; // @[:@29903.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@29905.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@29904.4]
  assign RetimeWrapper_8_clock = clock; // @[:@29920.4]
  assign RetimeWrapper_8_reset = reset; // @[:@29921.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@29923.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@29922.4]
  assign RetimeWrapper_9_clock = clock; // @[:@29977.4]
  assign RetimeWrapper_9_reset = reset; // @[:@29978.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@29980.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@29979.4]
  assign RetimeWrapper_10_clock = clock; // @[:@29994.4]
  assign RetimeWrapper_10_reset = reset; // @[:@29995.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@29997.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@29996.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x455_inr_UnitPipe_sm( // @[:@30173.2]
  input   clock, // @[:@30174.4]
  input   reset, // @[:@30175.4]
  input   io_enable, // @[:@30176.4]
  output  io_done, // @[:@30176.4]
  output  io_doneLatch, // @[:@30176.4]
  input   io_ctrDone, // @[:@30176.4]
  output  io_datapathEn, // @[:@30176.4]
  output  io_ctrInc, // @[:@30176.4]
  input   io_parentAck, // @[:@30176.4]
  input   io_backpressure // @[:@30176.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@30178.4]
  wire  active_reset; // @[Controllers.scala 261:22:@30178.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@30178.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@30178.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@30178.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@30178.4]
  wire  done_clock; // @[Controllers.scala 262:20:@30181.4]
  wire  done_reset; // @[Controllers.scala 262:20:@30181.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@30181.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@30181.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@30181.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@30181.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30235.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30235.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30235.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30235.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30235.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30243.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30243.4]
  wire  _T_80; // @[Controllers.scala 264:48:@30186.4]
  wire  _T_81; // @[Controllers.scala 264:46:@30187.4]
  wire  _T_82; // @[Controllers.scala 264:62:@30188.4]
  wire  _T_83; // @[Controllers.scala 264:60:@30189.4]
  wire  _T_100; // @[package.scala 100:49:@30206.4]
  reg  _T_103; // @[package.scala 48:56:@30207.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@30215.4]
  wire  _T_116; // @[Controllers.scala 283:41:@30223.4]
  wire  _T_117; // @[Controllers.scala 283:59:@30224.4]
  wire  _T_119; // @[Controllers.scala 284:37:@30227.4]
  reg  _T_125; // @[package.scala 48:56:@30231.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@30253.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@30256.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@30258.4]
  wire  _T_152; // @[Controllers.scala 292:61:@30259.4]
  wire  _T_153; // @[Controllers.scala 292:24:@30260.4]
  SRFF active ( // @[Controllers.scala 261:22:@30178.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@30181.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30235.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30243.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@30186.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@30187.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@30188.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@30189.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@30206.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@30215.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@30223.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@30224.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@30227.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@30258.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@30259.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@30260.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@30234.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@30262.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@30226.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@30229.4]
  assign active_clock = clock; // @[:@30179.4]
  assign active_reset = reset; // @[:@30180.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@30191.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@30195.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@30196.4]
  assign done_clock = clock; // @[:@30182.4]
  assign done_reset = reset; // @[:@30183.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@30211.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@30204.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@30205.4]
  assign RetimeWrapper_clock = clock; // @[:@30236.4]
  assign RetimeWrapper_reset = reset; // @[:@30237.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30239.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@30238.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30244.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30245.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30247.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@30246.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1( // @[:@30337.2]
  output        io_in_x448_valid, // @[:@30340.4]
  output [63:0] io_in_x448_bits_addr, // @[:@30340.4]
  output [31:0] io_in_x448_bits_size, // @[:@30340.4]
  input  [63:0] io_in_x251_outdram_number, // @[:@30340.4]
  input         io_sigsIn_backpressure, // @[:@30340.4]
  input         io_sigsIn_datapathEn, // @[:@30340.4]
  input         io_rr // @[:@30340.4]
);
  wire [96:0] x452_tuple; // @[Cat.scala 30:58:@30354.4]
  wire  _T_135; // @[implicits.scala 55:10:@30357.4]
  assign x452_tuple = {33'h7e9000,io_in_x251_outdram_number}; // @[Cat.scala 30:58:@30354.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@30357.4]
  assign io_in_x448_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x455_inr_UnitPipe.scala 65:18:@30360.4]
  assign io_in_x448_bits_addr = x452_tuple[63:0]; // @[sm_x455_inr_UnitPipe.scala 66:22:@30362.4]
  assign io_in_x448_bits_size = x452_tuple[95:64]; // @[sm_x455_inr_UnitPipe.scala 67:22:@30364.4]
endmodule
module FF_13( // @[:@30366.2]
  input         clock, // @[:@30367.4]
  input         reset, // @[:@30368.4]
  output [22:0] io_rPort_0_output_0, // @[:@30369.4]
  input  [22:0] io_wPort_0_data_0, // @[:@30369.4]
  input         io_wPort_0_reset, // @[:@30369.4]
  input         io_wPort_0_en_0 // @[:@30369.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@30384.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@30386.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@30387.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@30386.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@30387.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@30389.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@30404.2]
  input         clock, // @[:@30405.4]
  input         reset, // @[:@30406.4]
  input         io_input_reset, // @[:@30407.4]
  input         io_input_enable, // @[:@30407.4]
  output [22:0] io_output_count_0, // @[:@30407.4]
  output        io_output_oobs_0, // @[:@30407.4]
  output        io_output_done // @[:@30407.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@30420.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@30420.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@30420.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@30420.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@30420.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@30420.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@30436.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@30436.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@30436.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@30436.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@30436.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@30436.4]
  wire  _T_36; // @[Counter.scala 264:45:@30439.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@30464.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@30465.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@30466.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@30467.4]
  wire  _T_57; // @[Counter.scala 293:18:@30469.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@30477.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@30480.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@30481.4]
  wire  _T_75; // @[Counter.scala 322:102:@30485.4]
  wire  _T_77; // @[Counter.scala 322:130:@30486.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@30420.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@30436.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@30439.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@30464.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@30465.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@30466.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@30467.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@30469.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@30477.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@30480.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@30481.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@30485.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@30486.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@30484.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@30488.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@30490.4]
  assign bases_0_clock = clock; // @[:@30421.4]
  assign bases_0_reset = reset; // @[:@30422.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@30483.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@30462.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@30463.4]
  assign SRFF_clock = clock; // @[:@30437.4]
  assign SRFF_reset = reset; // @[:@30438.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@30441.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@30443.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@30444.4]
endmodule
module x457_ctrchain( // @[:@30495.2]
  input         clock, // @[:@30496.4]
  input         reset, // @[:@30497.4]
  input         io_input_reset, // @[:@30498.4]
  input         io_input_enable, // @[:@30498.4]
  output [22:0] io_output_counts_0, // @[:@30498.4]
  output        io_output_oobs_0, // @[:@30498.4]
  output        io_output_done // @[:@30498.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@30500.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@30500.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@30500.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@30500.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@30500.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@30500.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@30500.4]
  reg  wasDone; // @[Counter.scala 542:24:@30509.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@30515.4]
  wire  _T_47; // @[Counter.scala 546:80:@30516.4]
  reg  doneLatch; // @[Counter.scala 550:26:@30521.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@30522.4]
  wire  _T_55; // @[Counter.scala 551:19:@30523.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@30500.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@30515.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@30516.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@30522.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@30523.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@30525.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@30527.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@30518.4]
  assign ctrs_0_clock = clock; // @[:@30501.4]
  assign ctrs_0_reset = reset; // @[:@30502.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@30506.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@30507.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x464_inr_Foreach_sm( // @[:@30715.2]
  input   clock, // @[:@30716.4]
  input   reset, // @[:@30717.4]
  input   io_enable, // @[:@30718.4]
  output  io_done, // @[:@30718.4]
  output  io_doneLatch, // @[:@30718.4]
  input   io_ctrDone, // @[:@30718.4]
  output  io_datapathEn, // @[:@30718.4]
  output  io_ctrInc, // @[:@30718.4]
  output  io_ctrRst, // @[:@30718.4]
  input   io_parentAck, // @[:@30718.4]
  input   io_backpressure, // @[:@30718.4]
  input   io_break // @[:@30718.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@30720.4]
  wire  active_reset; // @[Controllers.scala 261:22:@30720.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@30720.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@30720.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@30720.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@30720.4]
  wire  done_clock; // @[Controllers.scala 262:20:@30723.4]
  wire  done_reset; // @[Controllers.scala 262:20:@30723.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@30723.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@30723.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@30723.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@30723.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30757.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30757.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30757.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30757.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30757.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30779.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30779.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30779.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30779.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30779.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30791.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30791.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30791.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30791.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30791.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30799.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30815.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30815.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30815.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30815.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30815.4]
  wire  _T_80; // @[Controllers.scala 264:48:@30728.4]
  wire  _T_81; // @[Controllers.scala 264:46:@30729.4]
  wire  _T_82; // @[Controllers.scala 264:62:@30730.4]
  wire  _T_83; // @[Controllers.scala 264:60:@30731.4]
  wire  _T_100; // @[package.scala 100:49:@30748.4]
  reg  _T_103; // @[package.scala 48:56:@30749.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@30762.4 package.scala 96:25:@30763.4]
  wire  _T_110; // @[package.scala 100:49:@30764.4]
  reg  _T_113; // @[package.scala 48:56:@30765.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@30767.4]
  wire  _T_118; // @[Controllers.scala 283:41:@30772.4]
  wire  _T_119; // @[Controllers.scala 283:59:@30773.4]
  wire  _T_121; // @[Controllers.scala 284:37:@30776.4]
  wire  _T_124; // @[package.scala 96:25:@30784.4 package.scala 96:25:@30785.4]
  wire  _T_126; // @[package.scala 100:49:@30786.4]
  reg  _T_129; // @[package.scala 48:56:@30787.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@30809.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@30811.4]
  reg  _T_153; // @[package.scala 48:56:@30812.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@30820.4 package.scala 96:25:@30821.4]
  wire  _T_158; // @[Controllers.scala 292:61:@30822.4]
  wire  _T_159; // @[Controllers.scala 292:24:@30823.4]
  SRFF active ( // @[Controllers.scala 261:22:@30720.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@30723.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@30757.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@30779.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30791.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30799.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30815.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@30728.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@30729.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@30730.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@30731.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@30748.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@30762.4 package.scala 96:25:@30763.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@30764.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@30767.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@30772.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@30773.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@30776.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30784.4 package.scala 96:25:@30785.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@30786.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@30811.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30820.4 package.scala 96:25:@30821.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@30822.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@30823.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@30790.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@30825.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@30775.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@30778.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@30770.4]
  assign active_clock = clock; // @[:@30721.4]
  assign active_reset = reset; // @[:@30722.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@30733.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@30737.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@30738.4]
  assign done_clock = clock; // @[:@30724.4]
  assign done_reset = reset; // @[:@30725.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@30753.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@30746.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@30747.4]
  assign RetimeWrapper_clock = clock; // @[:@30758.4]
  assign RetimeWrapper_reset = reset; // @[:@30759.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@30761.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@30760.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30780.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30781.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@30783.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@30782.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30792.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30793.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30795.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@30794.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30800.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30801.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30803.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@30802.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30816.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30817.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@30819.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@30818.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x464_inr_Foreach_kernelx464_inr_Foreach_concrete1( // @[:@31032.2]
  input         clock, // @[:@31033.4]
  input         reset, // @[:@31034.4]
  output        io_in_x449_valid, // @[:@31035.4]
  output [31:0] io_in_x449_bits_wdata_0, // @[:@31035.4]
  output        io_in_x449_bits_wstrb, // @[:@31035.4]
  output [20:0] io_in_x255_outbuf_0_rPort_0_ofs_0, // @[:@31035.4]
  output        io_in_x255_outbuf_0_rPort_0_en_0, // @[:@31035.4]
  output        io_in_x255_outbuf_0_rPort_0_backpressure, // @[:@31035.4]
  input  [31:0] io_in_x255_outbuf_0_rPort_0_output_0, // @[:@31035.4]
  input         io_sigsIn_backpressure, // @[:@31035.4]
  input         io_sigsIn_datapathEn, // @[:@31035.4]
  input         io_sigsIn_break, // @[:@31035.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@31035.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@31035.4]
  input         io_rr // @[:@31035.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@31062.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@31062.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31091.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31091.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31091.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31091.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31091.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31100.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31100.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31100.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31100.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31100.4]
  wire  b459; // @[sm_x464_inr_Foreach.scala 62:18:@31070.4]
  wire  _T_274; // @[sm_x464_inr_Foreach.scala 67:129:@31074.4]
  wire  _T_278; // @[implicits.scala 55:10:@31077.4]
  wire  _T_279; // @[sm_x464_inr_Foreach.scala 67:146:@31078.4]
  wire [32:0] x462_tuple; // @[Cat.scala 30:58:@31088.4]
  wire  _T_290; // @[package.scala 96:25:@31105.4 package.scala 96:25:@31106.4]
  wire  _T_292; // @[implicits.scala 55:10:@31107.4]
  wire  x589_b459_D2; // @[package.scala 96:25:@31096.4 package.scala 96:25:@31097.4]
  wire  _T_293; // @[sm_x464_inr_Foreach.scala 74:112:@31108.4]
  wire [31:0] b458_number; // @[Math.scala 723:22:@31067.4 Math.scala 724:14:@31068.4]
  _ _ ( // @[Math.scala 720:24:@31062.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@31091.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@31100.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b459 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x464_inr_Foreach.scala 62:18:@31070.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x464_inr_Foreach.scala 67:129:@31074.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@31077.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x464_inr_Foreach.scala 67:146:@31078.4]
  assign x462_tuple = {1'h1,io_in_x255_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@31088.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31105.4 package.scala 96:25:@31106.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@31107.4]
  assign x589_b459_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@31096.4 package.scala 96:25:@31097.4]
  assign _T_293 = _T_292 & x589_b459_D2; // @[sm_x464_inr_Foreach.scala 74:112:@31108.4]
  assign b458_number = __io_result; // @[Math.scala 723:22:@31067.4 Math.scala 724:14:@31068.4]
  assign io_in_x449_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x464_inr_Foreach.scala 74:18:@31110.4]
  assign io_in_x449_bits_wdata_0 = x462_tuple[31:0]; // @[sm_x464_inr_Foreach.scala 75:26:@31112.4]
  assign io_in_x449_bits_wstrb = x462_tuple[32]; // @[sm_x464_inr_Foreach.scala 76:23:@31114.4]
  assign io_in_x255_outbuf_0_rPort_0_ofs_0 = b458_number[20:0]; // @[MemInterfaceType.scala 107:54:@31081.4]
  assign io_in_x255_outbuf_0_rPort_0_en_0 = _T_279 & b459; // @[MemInterfaceType.scala 110:79:@31083.4]
  assign io_in_x255_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31082.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@31065.4]
  assign RetimeWrapper_clock = clock; // @[:@31092.4]
  assign RetimeWrapper_reset = reset; // @[:@31093.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31095.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@31094.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31101.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31102.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31104.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31103.4]
endmodule
module x468_inr_UnitPipe_sm( // @[:@31270.2]
  input   clock, // @[:@31271.4]
  input   reset, // @[:@31272.4]
  input   io_enable, // @[:@31273.4]
  output  io_done, // @[:@31273.4]
  output  io_doneLatch, // @[:@31273.4]
  input   io_ctrDone, // @[:@31273.4]
  output  io_datapathEn, // @[:@31273.4]
  output  io_ctrInc, // @[:@31273.4]
  input   io_parentAck // @[:@31273.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31275.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31275.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31275.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31275.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31275.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31275.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31278.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31278.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31278.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31278.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31278.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31278.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31312.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31312.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31312.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31312.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31312.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31334.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31334.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31334.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31334.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31334.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31346.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31346.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31346.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31346.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31346.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31354.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31354.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31354.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31354.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31354.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31283.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31284.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31285.4]
  wire  _T_100; // @[package.scala 100:49:@31303.4]
  reg  _T_103; // @[package.scala 48:56:@31304.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@31327.4]
  wire  _T_124; // @[package.scala 96:25:@31339.4 package.scala 96:25:@31340.4]
  wire  _T_126; // @[package.scala 100:49:@31341.4]
  reg  _T_129; // @[package.scala 48:56:@31342.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@31364.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@31366.4]
  reg  _T_153; // @[package.scala 48:56:@31367.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@31369.4]
  wire  _T_156; // @[Controllers.scala 292:61:@31370.4]
  wire  _T_157; // @[Controllers.scala 292:24:@31371.4]
  SRFF active ( // @[Controllers.scala 261:22:@31275.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31278.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31312.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31334.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31346.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31354.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31283.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31284.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31285.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31303.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31327.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31339.4 package.scala 96:25:@31340.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@31341.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@31366.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@31369.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@31370.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@31371.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@31345.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@31373.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@31330.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@31333.4]
  assign active_clock = clock; // @[:@31276.4]
  assign active_reset = reset; // @[:@31277.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@31288.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31292.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31293.4]
  assign done_clock = clock; // @[:@31279.4]
  assign done_reset = reset; // @[:@31280.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31308.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31301.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31302.4]
  assign RetimeWrapper_clock = clock; // @[:@31313.4]
  assign RetimeWrapper_reset = reset; // @[:@31314.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31316.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@31315.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31335.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31336.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31338.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@31337.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31347.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31348.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31350.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@31349.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31355.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31356.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31358.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@31357.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1( // @[:@31448.2]
  output  io_in_x450_ready, // @[:@31451.4]
  input   io_sigsIn_datapathEn // @[:@31451.4]
);
  assign io_in_x450_ready = io_sigsIn_datapathEn; // @[sm_x468_inr_UnitPipe.scala 57:18:@31463.4]
endmodule
module x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1( // @[:@31466.2]
  input         clock, // @[:@31467.4]
  input         reset, // @[:@31468.4]
  input         io_in_x449_ready, // @[:@31469.4]
  output        io_in_x449_valid, // @[:@31469.4]
  output [31:0] io_in_x449_bits_wdata_0, // @[:@31469.4]
  output        io_in_x449_bits_wstrb, // @[:@31469.4]
  input         io_in_x448_ready, // @[:@31469.4]
  output        io_in_x448_valid, // @[:@31469.4]
  output [63:0] io_in_x448_bits_addr, // @[:@31469.4]
  output [31:0] io_in_x448_bits_size, // @[:@31469.4]
  input  [63:0] io_in_x251_outdram_number, // @[:@31469.4]
  output [20:0] io_in_x255_outbuf_0_rPort_0_ofs_0, // @[:@31469.4]
  output        io_in_x255_outbuf_0_rPort_0_en_0, // @[:@31469.4]
  output        io_in_x255_outbuf_0_rPort_0_backpressure, // @[:@31469.4]
  input  [31:0] io_in_x255_outbuf_0_rPort_0_output_0, // @[:@31469.4]
  output        io_in_x450_ready, // @[:@31469.4]
  input         io_in_x450_valid, // @[:@31469.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@31469.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@31469.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@31469.4]
  input         io_sigsIn_smChildAcks_0, // @[:@31469.4]
  input         io_sigsIn_smChildAcks_1, // @[:@31469.4]
  input         io_sigsIn_smChildAcks_2, // @[:@31469.4]
  output        io_sigsOut_smDoneIn_0, // @[:@31469.4]
  output        io_sigsOut_smDoneIn_1, // @[:@31469.4]
  output        io_sigsOut_smDoneIn_2, // @[:@31469.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@31469.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@31469.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@31469.4]
  input         io_rr // @[:@31469.4]
);
  wire  x455_inr_UnitPipe_sm_clock; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_reset; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_enable; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_done; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_doneLatch; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_ctrDone; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_datapathEn; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_ctrInc; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_parentAck; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  x455_inr_UnitPipe_sm_io_backpressure; // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31601.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31601.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31601.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31601.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31601.4]
  wire  x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_valid; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire [63:0] x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_bits_addr; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire [31:0] x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_bits_size; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire [63:0] x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x251_outdram_number; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire  x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire  x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire  x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_rr; // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
  wire  x457_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire  x457_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire  x457_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire  x457_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire [22:0] x457_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire  x457_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire  x457_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@31699.4]
  wire  x464_inr_Foreach_sm_clock; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_reset; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_enable; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_done; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_doneLatch; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_ctrDone; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_datapathEn; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_ctrInc; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_ctrRst; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_parentAck; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_backpressure; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  x464_inr_Foreach_sm_io_break; // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31780.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31780.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31780.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31780.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31780.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31820.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31820.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31820.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31820.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31820.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31828.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31828.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31828.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@31828.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@31828.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_clock; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_reset; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_valid; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire [31:0] x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_bits_wdata_0; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_bits_wstrb; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire [20:0] x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_en_0; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire [31:0] x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_output_0; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire [31:0] x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_rr; // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
  wire  x468_inr_UnitPipe_sm_clock; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_reset; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_enable; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_done; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_doneLatch; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_ctrDone; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_datapathEn; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_ctrInc; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  x468_inr_UnitPipe_sm_io_parentAck; // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@32040.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@32040.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@32040.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@32040.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@32040.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@32048.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@32048.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@32048.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@32048.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@32048.4]
  wire  x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1_io_in_x450_ready; // @[sm_x468_inr_UnitPipe.scala 60:24:@32078.4]
  wire  x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x468_inr_UnitPipe.scala 60:24:@32078.4]
  wire  _T_359; // @[package.scala 100:49:@31564.4]
  reg  _T_362; // @[package.scala 48:56:@31565.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@31598.4 package.scala 96:25:@31599.4]
  wire  _T_381; // @[package.scala 96:25:@31606.4 package.scala 96:25:@31607.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@31609.4]
  wire  _T_454; // @[package.scala 96:25:@31785.4 package.scala 96:25:@31786.4]
  wire  _T_468; // @[package.scala 96:25:@31825.4 package.scala 96:25:@31826.4]
  wire  _T_474; // @[package.scala 96:25:@31833.4 package.scala 96:25:@31834.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@31836.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@31845.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@31846.4]
  wire  _T_547; // @[package.scala 100:49:@32011.4]
  reg  _T_550; // @[package.scala 48:56:@32012.4]
  reg [31:0] _RAND_1;
  wire  x468_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x469_outr_UnitPipe.scala 101:55:@32018.4]
  wire  _T_563; // @[package.scala 96:25:@32045.4 package.scala 96:25:@32046.4]
  wire  _T_569; // @[package.scala 96:25:@32053.4 package.scala 96:25:@32054.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@32056.4]
  wire  x468_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@32057.4]
  x455_inr_UnitPipe_sm x455_inr_UnitPipe_sm ( // @[sm_x455_inr_UnitPipe.scala 33:18:@31536.4]
    .clock(x455_inr_UnitPipe_sm_clock),
    .reset(x455_inr_UnitPipe_sm_reset),
    .io_enable(x455_inr_UnitPipe_sm_io_enable),
    .io_done(x455_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x455_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x455_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x455_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x455_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x455_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x455_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31593.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31601.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1 x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1 ( // @[sm_x455_inr_UnitPipe.scala 69:24:@31631.4]
    .io_in_x448_valid(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_valid),
    .io_in_x448_bits_addr(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_bits_addr),
    .io_in_x448_bits_size(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_bits_size),
    .io_in_x251_outdram_number(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x251_outdram_number),
    .io_sigsIn_backpressure(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_rr)
  );
  x457_ctrchain x457_ctrchain ( // @[SpatialBlocks.scala 37:22:@31699.4]
    .clock(x457_ctrchain_clock),
    .reset(x457_ctrchain_reset),
    .io_input_reset(x457_ctrchain_io_input_reset),
    .io_input_enable(x457_ctrchain_io_input_enable),
    .io_output_counts_0(x457_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x457_ctrchain_io_output_oobs_0),
    .io_output_done(x457_ctrchain_io_output_done)
  );
  x464_inr_Foreach_sm x464_inr_Foreach_sm ( // @[sm_x464_inr_Foreach.scala 33:18:@31752.4]
    .clock(x464_inr_Foreach_sm_clock),
    .reset(x464_inr_Foreach_sm_reset),
    .io_enable(x464_inr_Foreach_sm_io_enable),
    .io_done(x464_inr_Foreach_sm_io_done),
    .io_doneLatch(x464_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x464_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x464_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x464_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x464_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x464_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x464_inr_Foreach_sm_io_backpressure),
    .io_break(x464_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31780.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31820.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@31828.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x464_inr_Foreach_kernelx464_inr_Foreach_concrete1 x464_inr_Foreach_kernelx464_inr_Foreach_concrete1 ( // @[sm_x464_inr_Foreach.scala 78:24:@31863.4]
    .clock(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_clock),
    .reset(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_reset),
    .io_in_x449_valid(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_valid),
    .io_in_x449_bits_wdata_0(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_bits_wdata_0),
    .io_in_x449_bits_wstrb(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_bits_wstrb),
    .io_in_x255_outbuf_0_rPort_0_ofs_0(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0),
    .io_in_x255_outbuf_0_rPort_0_en_0(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_en_0),
    .io_in_x255_outbuf_0_rPort_0_backpressure(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure),
    .io_in_x255_outbuf_0_rPort_0_output_0(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_output_0),
    .io_sigsIn_backpressure(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_rr)
  );
  x468_inr_UnitPipe_sm x468_inr_UnitPipe_sm ( // @[sm_x468_inr_UnitPipe.scala 32:18:@31983.4]
    .clock(x468_inr_UnitPipe_sm_clock),
    .reset(x468_inr_UnitPipe_sm_reset),
    .io_enable(x468_inr_UnitPipe_sm_io_enable),
    .io_done(x468_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x468_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x468_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x468_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x468_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x468_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@32040.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@32048.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1 x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1 ( // @[sm_x468_inr_UnitPipe.scala 60:24:@32078.4]
    .io_in_x450_ready(x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1_io_in_x450_ready),
    .io_sigsIn_datapathEn(x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x455_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@31564.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@31598.4 package.scala 96:25:@31599.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31606.4 package.scala 96:25:@31607.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@31609.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@31785.4 package.scala 96:25:@31786.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@31825.4 package.scala 96:25:@31826.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31833.4 package.scala 96:25:@31834.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@31836.4]
  assign _T_479 = x464_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@31845.4]
  assign _T_480 = ~ x464_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@31846.4]
  assign _T_547 = x468_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32011.4]
  assign x468_inr_UnitPipe_sigsIn_forwardpressure = io_in_x450_valid | x468_inr_UnitPipe_sm_io_doneLatch; // @[sm_x469_outr_UnitPipe.scala 101:55:@32018.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@32045.4 package.scala 96:25:@32046.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@32053.4 package.scala 96:25:@32054.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@32056.4]
  assign x468_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@32057.4]
  assign io_in_x449_valid = x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_valid; // @[sm_x464_inr_Foreach.scala 49:23:@31913.4]
  assign io_in_x449_bits_wdata_0 = x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_bits_wdata_0; // @[sm_x464_inr_Foreach.scala 49:23:@31912.4]
  assign io_in_x449_bits_wstrb = x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x449_bits_wstrb; // @[sm_x464_inr_Foreach.scala 49:23:@31911.4]
  assign io_in_x448_valid = x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_valid; // @[sm_x455_inr_UnitPipe.scala 49:23:@31669.4]
  assign io_in_x448_bits_addr = x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_bits_addr; // @[sm_x455_inr_UnitPipe.scala 49:23:@31668.4]
  assign io_in_x448_bits_size = x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x448_bits_size; // @[sm_x455_inr_UnitPipe.scala 49:23:@31667.4]
  assign io_in_x255_outbuf_0_rPort_0_ofs_0 = x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@31918.4]
  assign io_in_x255_outbuf_0_rPort_0_en_0 = x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@31917.4]
  assign io_in_x255_outbuf_0_rPort_0_backpressure = x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@31916.4]
  assign io_in_x450_ready = x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1_io_in_x450_ready; // @[sm_x468_inr_UnitPipe.scala 46:23:@32114.4]
  assign io_sigsOut_smDoneIn_0 = x455_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31616.4]
  assign io_sigsOut_smDoneIn_1 = x464_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@31843.4]
  assign io_sigsOut_smDoneIn_2 = x468_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@32063.4]
  assign io_sigsOut_smCtrCopyDone_0 = x455_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@31630.4]
  assign io_sigsOut_smCtrCopyDone_1 = x464_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@31862.4]
  assign io_sigsOut_smCtrCopyDone_2 = x468_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@32077.4]
  assign x455_inr_UnitPipe_sm_clock = clock; // @[:@31537.4]
  assign x455_inr_UnitPipe_sm_reset = reset; // @[:@31538.4]
  assign x455_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@31613.4]
  assign x455_inr_UnitPipe_sm_io_ctrDone = x455_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x469_outr_UnitPipe.scala 77:39:@31568.4]
  assign x455_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@31615.4]
  assign x455_inr_UnitPipe_sm_io_backpressure = io_in_x448_ready | x455_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@31587.4]
  assign RetimeWrapper_clock = clock; // @[:@31594.4]
  assign RetimeWrapper_reset = reset; // @[:@31595.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31597.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@31596.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31602.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31603.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31605.4]
  assign RetimeWrapper_1_io_in = x455_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31604.4]
  assign x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_in_x251_outdram_number = io_in_x251_outdram_number; // @[sm_x455_inr_UnitPipe.scala 50:31:@31671.4]
  assign x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x448_ready | x455_inr_UnitPipe_sm_io_doneLatch; // @[sm_x455_inr_UnitPipe.scala 74:22:@31686.4]
  assign x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x455_inr_UnitPipe_sm_io_datapathEn; // @[sm_x455_inr_UnitPipe.scala 74:22:@31684.4]
  assign x455_inr_UnitPipe_kernelx455_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x455_inr_UnitPipe.scala 73:18:@31672.4]
  assign x457_ctrchain_clock = clock; // @[:@31700.4]
  assign x457_ctrchain_reset = reset; // @[:@31701.4]
  assign x457_ctrchain_io_input_reset = x464_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@31861.4]
  assign x457_ctrchain_io_input_enable = x464_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@31813.4 SpatialBlocks.scala 159:42:@31860.4]
  assign x464_inr_Foreach_sm_clock = clock; // @[:@31753.4]
  assign x464_inr_Foreach_sm_reset = reset; // @[:@31754.4]
  assign x464_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@31840.4]
  assign x464_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x469_outr_UnitPipe.scala 90:38:@31788.4]
  assign x464_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@31842.4]
  assign x464_inr_Foreach_sm_io_backpressure = io_in_x449_ready | x464_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@31814.4]
  assign x464_inr_Foreach_sm_io_break = 1'h0; // @[sm_x469_outr_UnitPipe.scala 94:36:@31794.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31781.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31782.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31784.4]
  assign RetimeWrapper_2_io_in = x457_ctrchain_io_output_done; // @[package.scala 94:16:@31783.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31821.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31822.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31824.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@31823.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31829.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31830.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@31832.4]
  assign RetimeWrapper_4_io_in = x464_inr_Foreach_sm_io_done; // @[package.scala 94:16:@31831.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_clock = clock; // @[:@31864.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_reset = reset; // @[:@31865.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_in_x255_outbuf_0_rPort_0_output_0 = io_in_x255_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@31915.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x449_ready | x464_inr_Foreach_sm_io_doneLatch; // @[sm_x464_inr_Foreach.scala 83:22:@31934.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x464_inr_Foreach.scala 83:22:@31932.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_break = x464_inr_Foreach_sm_io_break; // @[sm_x464_inr_Foreach.scala 83:22:@31930.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x457_ctrchain_io_output_counts_0[22]}},x457_ctrchain_io_output_counts_0}; // @[sm_x464_inr_Foreach.scala 83:22:@31925.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x457_ctrchain_io_output_oobs_0; // @[sm_x464_inr_Foreach.scala 83:22:@31924.4]
  assign x464_inr_Foreach_kernelx464_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x464_inr_Foreach.scala 82:18:@31920.4]
  assign x468_inr_UnitPipe_sm_clock = clock; // @[:@31984.4]
  assign x468_inr_UnitPipe_sm_reset = reset; // @[:@31985.4]
  assign x468_inr_UnitPipe_sm_io_enable = x468_inr_UnitPipe_sigsIn_baseEn & x468_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@32060.4]
  assign x468_inr_UnitPipe_sm_io_ctrDone = x468_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x469_outr_UnitPipe.scala 99:39:@32015.4]
  assign x468_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@32062.4]
  assign RetimeWrapper_5_clock = clock; // @[:@32041.4]
  assign RetimeWrapper_5_reset = reset; // @[:@32042.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@32044.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@32043.4]
  assign RetimeWrapper_6_clock = clock; // @[:@32049.4]
  assign RetimeWrapper_6_reset = reset; // @[:@32050.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@32052.4]
  assign RetimeWrapper_6_io_in = x468_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@32051.4]
  assign x468_inr_UnitPipe_kernelx468_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x468_inr_UnitPipe_sm_io_datapathEn; // @[sm_x468_inr_UnitPipe.scala 65:22:@32127.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x522_kernelx522_concrete1( // @[:@32143.2]
  input          clock, // @[:@32144.4]
  input          reset, // @[:@32145.4]
  input          io_in_x449_ready, // @[:@32146.4]
  output         io_in_x449_valid, // @[:@32146.4]
  output [31:0]  io_in_x449_bits_wdata_0, // @[:@32146.4]
  output         io_in_x449_bits_wstrb, // @[:@32146.4]
  input          io_in_x448_ready, // @[:@32146.4]
  output         io_in_x448_valid, // @[:@32146.4]
  output [63:0]  io_in_x448_bits_addr, // @[:@32146.4]
  output [31:0]  io_in_x448_bits_size, // @[:@32146.4]
  input          io_in_x253_TVALID, // @[:@32146.4]
  output         io_in_x253_TREADY, // @[:@32146.4]
  input  [255:0] io_in_x253_TDATA, // @[:@32146.4]
  input  [7:0]   io_in_x253_TID, // @[:@32146.4]
  input  [7:0]   io_in_x253_TDEST, // @[:@32146.4]
  input  [63:0]  io_in_x251_outdram_number, // @[:@32146.4]
  output [20:0]  io_in_x255_outbuf_0_rPort_0_ofs_0, // @[:@32146.4]
  output         io_in_x255_outbuf_0_rPort_0_en_0, // @[:@32146.4]
  output         io_in_x255_outbuf_0_rPort_0_backpressure, // @[:@32146.4]
  input  [31:0]  io_in_x255_outbuf_0_rPort_0_output_0, // @[:@32146.4]
  output         io_in_x450_ready, // @[:@32146.4]
  input          io_in_x450_valid, // @[:@32146.4]
  output         io_in_x254_TVALID, // @[:@32146.4]
  input          io_in_x254_TREADY, // @[:@32146.4]
  output [255:0] io_in_x254_TDATA, // @[:@32146.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@32146.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@32146.4]
  input          io_sigsIn_smChildAcks_0, // @[:@32146.4]
  input          io_sigsIn_smChildAcks_1, // @[:@32146.4]
  output         io_sigsOut_smDoneIn_0, // @[:@32146.4]
  output         io_sigsOut_smDoneIn_1, // @[:@32146.4]
  input          io_rr // @[:@32146.4]
);
  wire  x447_outr_UnitPipe_sm_clock; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_reset; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_enable; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_done; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_parentAck; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_childAck_0; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_childAck_1; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  x447_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32281.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32281.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32281.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32281.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32281.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32289.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32289.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_clock; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_reset; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TVALID; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TREADY; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire [255:0] x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TDATA; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire [7:0] x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TID; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire [7:0] x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TDEST; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TVALID; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TREADY; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire [255:0] x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TDATA; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_rr; // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
  wire  x469_outr_UnitPipe_sm_clock; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_reset; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_enable; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_done; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_parentAck; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_childAck_0; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_childAck_1; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_childAck_2; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  x469_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32570.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32570.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32570.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32570.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32570.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32578.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32578.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32578.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32578.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32578.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_clock; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_reset; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_ready; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_valid; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire [31:0] x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_bits_wdata_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_bits_wstrb; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_ready; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_valid; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire [63:0] x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_bits_addr; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire [31:0] x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_bits_size; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire [63:0] x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x251_outdram_number; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire [20:0] x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_en_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire [31:0] x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_output_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x450_ready; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x450_valid; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_rr; // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
  wire  _T_408; // @[package.scala 96:25:@32286.4 package.scala 96:25:@32287.4]
  wire  _T_414; // @[package.scala 96:25:@32294.4 package.scala 96:25:@32295.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@32297.4]
  wire  _T_508; // @[package.scala 96:25:@32575.4 package.scala 96:25:@32576.4]
  wire  _T_514; // @[package.scala 96:25:@32583.4 package.scala 96:25:@32584.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@32586.4]
  x447_outr_UnitPipe_sm x447_outr_UnitPipe_sm ( // @[sm_x447_outr_UnitPipe.scala 32:18:@32219.4]
    .clock(x447_outr_UnitPipe_sm_clock),
    .reset(x447_outr_UnitPipe_sm_reset),
    .io_enable(x447_outr_UnitPipe_sm_io_enable),
    .io_done(x447_outr_UnitPipe_sm_io_done),
    .io_parentAck(x447_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x447_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x447_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x447_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x447_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x447_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x447_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x447_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x447_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32281.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32289.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1 x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1 ( // @[sm_x447_outr_UnitPipe.scala 87:24:@32320.4]
    .clock(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_clock),
    .reset(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_reset),
    .io_in_x253_TVALID(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TVALID),
    .io_in_x253_TREADY(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TREADY),
    .io_in_x253_TDATA(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TDATA),
    .io_in_x253_TID(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TID),
    .io_in_x253_TDEST(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TDEST),
    .io_in_x254_TVALID(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TVALID),
    .io_in_x254_TREADY(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TREADY),
    .io_in_x254_TDATA(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TDATA),
    .io_sigsIn_smEnableOuts_0(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_rr)
  );
  x469_outr_UnitPipe_sm x469_outr_UnitPipe_sm ( // @[sm_x469_outr_UnitPipe.scala 36:18:@32498.4]
    .clock(x469_outr_UnitPipe_sm_clock),
    .reset(x469_outr_UnitPipe_sm_reset),
    .io_enable(x469_outr_UnitPipe_sm_io_enable),
    .io_done(x469_outr_UnitPipe_sm_io_done),
    .io_parentAck(x469_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x469_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x469_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x469_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x469_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x469_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x469_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x469_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x469_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x469_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x469_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x469_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x469_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32570.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32578.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1 x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1 ( // @[sm_x469_outr_UnitPipe.scala 108:24:@32610.4]
    .clock(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_clock),
    .reset(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_reset),
    .io_in_x449_ready(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_ready),
    .io_in_x449_valid(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_valid),
    .io_in_x449_bits_wdata_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_bits_wdata_0),
    .io_in_x449_bits_wstrb(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_bits_wstrb),
    .io_in_x448_ready(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_ready),
    .io_in_x448_valid(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_valid),
    .io_in_x448_bits_addr(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_bits_addr),
    .io_in_x448_bits_size(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_bits_size),
    .io_in_x251_outdram_number(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x251_outdram_number),
    .io_in_x255_outbuf_0_rPort_0_ofs_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0),
    .io_in_x255_outbuf_0_rPort_0_en_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_en_0),
    .io_in_x255_outbuf_0_rPort_0_backpressure(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure),
    .io_in_x255_outbuf_0_rPort_0_output_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_output_0),
    .io_in_x450_ready(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x450_ready),
    .io_in_x450_valid(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x450_valid),
    .io_sigsIn_smEnableOuts_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@32286.4 package.scala 96:25:@32287.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32294.4 package.scala 96:25:@32295.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@32297.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@32575.4 package.scala 96:25:@32576.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32583.4 package.scala 96:25:@32584.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@32586.4]
  assign io_in_x449_valid = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_valid; // @[sm_x469_outr_UnitPipe.scala 58:23:@32692.4]
  assign io_in_x449_bits_wdata_0 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_bits_wdata_0; // @[sm_x469_outr_UnitPipe.scala 58:23:@32691.4]
  assign io_in_x449_bits_wstrb = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_bits_wstrb; // @[sm_x469_outr_UnitPipe.scala 58:23:@32690.4]
  assign io_in_x448_valid = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_valid; // @[sm_x469_outr_UnitPipe.scala 59:23:@32696.4]
  assign io_in_x448_bits_addr = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_bits_addr; // @[sm_x469_outr_UnitPipe.scala 59:23:@32695.4]
  assign io_in_x448_bits_size = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_bits_size; // @[sm_x469_outr_UnitPipe.scala 59:23:@32694.4]
  assign io_in_x253_TREADY = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TREADY; // @[sm_x447_outr_UnitPipe.scala 48:23:@32388.4]
  assign io_in_x255_outbuf_0_rPort_0_ofs_0 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@32702.4]
  assign io_in_x255_outbuf_0_rPort_0_en_0 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@32701.4]
  assign io_in_x255_outbuf_0_rPort_0_backpressure = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@32700.4]
  assign io_in_x450_ready = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x450_ready; // @[sm_x469_outr_UnitPipe.scala 62:23:@32706.4]
  assign io_in_x254_TVALID = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TVALID; // @[sm_x447_outr_UnitPipe.scala 49:23:@32398.4]
  assign io_in_x254_TDATA = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TDATA; // @[sm_x447_outr_UnitPipe.scala 49:23:@32396.4]
  assign io_sigsOut_smDoneIn_0 = x447_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@32304.4]
  assign io_sigsOut_smDoneIn_1 = x469_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@32593.4]
  assign x447_outr_UnitPipe_sm_clock = clock; // @[:@32220.4]
  assign x447_outr_UnitPipe_sm_reset = reset; // @[:@32221.4]
  assign x447_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@32301.4]
  assign x447_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@32303.4]
  assign x447_outr_UnitPipe_sm_io_doneIn_0 = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@32271.4]
  assign x447_outr_UnitPipe_sm_io_doneIn_1 = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@32272.4]
  assign x447_outr_UnitPipe_sm_io_ctrCopyDone_0 = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@32318.4]
  assign x447_outr_UnitPipe_sm_io_ctrCopyDone_1 = x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@32319.4]
  assign RetimeWrapper_clock = clock; // @[:@32282.4]
  assign RetimeWrapper_reset = reset; // @[:@32283.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32285.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@32284.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32290.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32291.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32293.4]
  assign RetimeWrapper_1_io_in = x447_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@32292.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_clock = clock; // @[:@32321.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_reset = reset; // @[:@32322.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TVALID = io_in_x253_TVALID; // @[sm_x447_outr_UnitPipe.scala 48:23:@32389.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TDATA = io_in_x253_TDATA; // @[sm_x447_outr_UnitPipe.scala 48:23:@32387.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TID = io_in_x253_TID; // @[sm_x447_outr_UnitPipe.scala 48:23:@32383.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x253_TDEST = io_in_x253_TDEST; // @[sm_x447_outr_UnitPipe.scala 48:23:@32382.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_in_x254_TREADY = io_in_x254_TREADY; // @[sm_x447_outr_UnitPipe.scala 49:23:@32397.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x447_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x447_outr_UnitPipe.scala 92:22:@32414.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x447_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x447_outr_UnitPipe.scala 92:22:@32415.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x447_outr_UnitPipe_sm_io_childAck_0; // @[sm_x447_outr_UnitPipe.scala 92:22:@32410.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x447_outr_UnitPipe_sm_io_childAck_1; // @[sm_x447_outr_UnitPipe.scala 92:22:@32411.4]
  assign x447_outr_UnitPipe_kernelx447_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x447_outr_UnitPipe.scala 91:18:@32399.4]
  assign x469_outr_UnitPipe_sm_clock = clock; // @[:@32499.4]
  assign x469_outr_UnitPipe_sm_reset = reset; // @[:@32500.4]
  assign x469_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@32590.4]
  assign x469_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@32592.4]
  assign x469_outr_UnitPipe_sm_io_doneIn_0 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@32558.4]
  assign x469_outr_UnitPipe_sm_io_doneIn_1 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@32559.4]
  assign x469_outr_UnitPipe_sm_io_doneIn_2 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@32560.4]
  assign x469_outr_UnitPipe_sm_io_ctrCopyDone_0 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@32607.4]
  assign x469_outr_UnitPipe_sm_io_ctrCopyDone_1 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@32608.4]
  assign x469_outr_UnitPipe_sm_io_ctrCopyDone_2 = x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@32609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32571.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32572.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32574.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@32573.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32579.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32580.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32582.4]
  assign RetimeWrapper_3_io_in = x469_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@32581.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_clock = clock; // @[:@32611.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_reset = reset; // @[:@32612.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x449_ready = io_in_x449_ready; // @[sm_x469_outr_UnitPipe.scala 58:23:@32693.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x448_ready = io_in_x448_ready; // @[sm_x469_outr_UnitPipe.scala 59:23:@32697.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x251_outdram_number = io_in_x251_outdram_number; // @[sm_x469_outr_UnitPipe.scala 60:31:@32698.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x255_outbuf_0_rPort_0_output_0 = io_in_x255_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@32699.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_in_x450_valid = io_in_x450_valid; // @[sm_x469_outr_UnitPipe.scala 62:23:@32705.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x469_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x469_outr_UnitPipe.scala 113:22:@32729.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x469_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x469_outr_UnitPipe.scala 113:22:@32730.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x469_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x469_outr_UnitPipe.scala 113:22:@32731.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x469_outr_UnitPipe_sm_io_childAck_0; // @[sm_x469_outr_UnitPipe.scala 113:22:@32723.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x469_outr_UnitPipe_sm_io_childAck_1; // @[sm_x469_outr_UnitPipe.scala 113:22:@32724.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x469_outr_UnitPipe_sm_io_childAck_2; // @[sm_x469_outr_UnitPipe.scala 113:22:@32725.4]
  assign x469_outr_UnitPipe_kernelx469_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x469_outr_UnitPipe.scala 112:18:@32707.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@32759.2]
  input          clock, // @[:@32760.4]
  input          reset, // @[:@32761.4]
  input          io_in_x449_ready, // @[:@32762.4]
  output         io_in_x449_valid, // @[:@32762.4]
  output [31:0]  io_in_x449_bits_wdata_0, // @[:@32762.4]
  output         io_in_x449_bits_wstrb, // @[:@32762.4]
  input          io_in_x448_ready, // @[:@32762.4]
  output         io_in_x448_valid, // @[:@32762.4]
  output [63:0]  io_in_x448_bits_addr, // @[:@32762.4]
  output [31:0]  io_in_x448_bits_size, // @[:@32762.4]
  input          io_in_x253_TVALID, // @[:@32762.4]
  output         io_in_x253_TREADY, // @[:@32762.4]
  input  [255:0] io_in_x253_TDATA, // @[:@32762.4]
  input  [7:0]   io_in_x253_TID, // @[:@32762.4]
  input  [7:0]   io_in_x253_TDEST, // @[:@32762.4]
  input  [63:0]  io_in_x251_outdram_number, // @[:@32762.4]
  output         io_in_x450_ready, // @[:@32762.4]
  input          io_in_x450_valid, // @[:@32762.4]
  output         io_in_x254_TVALID, // @[:@32762.4]
  input          io_in_x254_TREADY, // @[:@32762.4]
  output [255:0] io_in_x254_TDATA, // @[:@32762.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@32762.4]
  input          io_sigsIn_smChildAcks_0, // @[:@32762.4]
  output         io_sigsOut_smDoneIn_0, // @[:@32762.4]
  input          io_rr // @[:@32762.4]
);
  wire  x255_outbuf_0_clock; // @[m_x255_outbuf_0.scala 27:17:@32772.4]
  wire  x255_outbuf_0_reset; // @[m_x255_outbuf_0.scala 27:17:@32772.4]
  wire [20:0] x255_outbuf_0_io_rPort_0_ofs_0; // @[m_x255_outbuf_0.scala 27:17:@32772.4]
  wire  x255_outbuf_0_io_rPort_0_en_0; // @[m_x255_outbuf_0.scala 27:17:@32772.4]
  wire  x255_outbuf_0_io_rPort_0_backpressure; // @[m_x255_outbuf_0.scala 27:17:@32772.4]
  wire [31:0] x255_outbuf_0_io_rPort_0_output_0; // @[m_x255_outbuf_0.scala 27:17:@32772.4]
  wire  x522_sm_clock; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_reset; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_enable; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_done; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_ctrDone; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_ctrInc; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_parentAck; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_doneIn_0; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_doneIn_1; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_enableOut_0; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_enableOut_1; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_childAck_0; // @[sm_x522.scala 37:18:@32830.4]
  wire  x522_sm_io_childAck_1; // @[sm_x522.scala 37:18:@32830.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32897.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32905.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32905.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32905.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32905.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32905.4]
  wire  x522_kernelx522_concrete1_clock; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_reset; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x449_ready; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x449_valid; // @[sm_x522.scala 102:24:@32934.4]
  wire [31:0] x522_kernelx522_concrete1_io_in_x449_bits_wdata_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x449_bits_wstrb; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x448_ready; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x448_valid; // @[sm_x522.scala 102:24:@32934.4]
  wire [63:0] x522_kernelx522_concrete1_io_in_x448_bits_addr; // @[sm_x522.scala 102:24:@32934.4]
  wire [31:0] x522_kernelx522_concrete1_io_in_x448_bits_size; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x253_TVALID; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x253_TREADY; // @[sm_x522.scala 102:24:@32934.4]
  wire [255:0] x522_kernelx522_concrete1_io_in_x253_TDATA; // @[sm_x522.scala 102:24:@32934.4]
  wire [7:0] x522_kernelx522_concrete1_io_in_x253_TID; // @[sm_x522.scala 102:24:@32934.4]
  wire [7:0] x522_kernelx522_concrete1_io_in_x253_TDEST; // @[sm_x522.scala 102:24:@32934.4]
  wire [63:0] x522_kernelx522_concrete1_io_in_x251_outdram_number; // @[sm_x522.scala 102:24:@32934.4]
  wire [20:0] x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_en_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure; // @[sm_x522.scala 102:24:@32934.4]
  wire [31:0] x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_output_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x450_ready; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x450_valid; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x254_TVALID; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_in_x254_TREADY; // @[sm_x522.scala 102:24:@32934.4]
  wire [255:0] x522_kernelx522_concrete1_io_in_x254_TDATA; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x522.scala 102:24:@32934.4]
  wire  x522_kernelx522_concrete1_io_rr; // @[sm_x522.scala 102:24:@32934.4]
  wire  _T_266; // @[package.scala 100:49:@32863.4]
  reg  _T_269; // @[package.scala 48:56:@32864.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@32902.4 package.scala 96:25:@32903.4]
  wire  _T_289; // @[package.scala 96:25:@32910.4 package.scala 96:25:@32911.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@32913.4]
  x255_outbuf_0 x255_outbuf_0 ( // @[m_x255_outbuf_0.scala 27:17:@32772.4]
    .clock(x255_outbuf_0_clock),
    .reset(x255_outbuf_0_reset),
    .io_rPort_0_ofs_0(x255_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x255_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x255_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x255_outbuf_0_io_rPort_0_output_0)
  );
  x522_sm x522_sm ( // @[sm_x522.scala 37:18:@32830.4]
    .clock(x522_sm_clock),
    .reset(x522_sm_reset),
    .io_enable(x522_sm_io_enable),
    .io_done(x522_sm_io_done),
    .io_ctrDone(x522_sm_io_ctrDone),
    .io_ctrInc(x522_sm_io_ctrInc),
    .io_parentAck(x522_sm_io_parentAck),
    .io_doneIn_0(x522_sm_io_doneIn_0),
    .io_doneIn_1(x522_sm_io_doneIn_1),
    .io_enableOut_0(x522_sm_io_enableOut_0),
    .io_enableOut_1(x522_sm_io_enableOut_1),
    .io_childAck_0(x522_sm_io_childAck_0),
    .io_childAck_1(x522_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32897.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32905.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x522_kernelx522_concrete1 x522_kernelx522_concrete1 ( // @[sm_x522.scala 102:24:@32934.4]
    .clock(x522_kernelx522_concrete1_clock),
    .reset(x522_kernelx522_concrete1_reset),
    .io_in_x449_ready(x522_kernelx522_concrete1_io_in_x449_ready),
    .io_in_x449_valid(x522_kernelx522_concrete1_io_in_x449_valid),
    .io_in_x449_bits_wdata_0(x522_kernelx522_concrete1_io_in_x449_bits_wdata_0),
    .io_in_x449_bits_wstrb(x522_kernelx522_concrete1_io_in_x449_bits_wstrb),
    .io_in_x448_ready(x522_kernelx522_concrete1_io_in_x448_ready),
    .io_in_x448_valid(x522_kernelx522_concrete1_io_in_x448_valid),
    .io_in_x448_bits_addr(x522_kernelx522_concrete1_io_in_x448_bits_addr),
    .io_in_x448_bits_size(x522_kernelx522_concrete1_io_in_x448_bits_size),
    .io_in_x253_TVALID(x522_kernelx522_concrete1_io_in_x253_TVALID),
    .io_in_x253_TREADY(x522_kernelx522_concrete1_io_in_x253_TREADY),
    .io_in_x253_TDATA(x522_kernelx522_concrete1_io_in_x253_TDATA),
    .io_in_x253_TID(x522_kernelx522_concrete1_io_in_x253_TID),
    .io_in_x253_TDEST(x522_kernelx522_concrete1_io_in_x253_TDEST),
    .io_in_x251_outdram_number(x522_kernelx522_concrete1_io_in_x251_outdram_number),
    .io_in_x255_outbuf_0_rPort_0_ofs_0(x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0),
    .io_in_x255_outbuf_0_rPort_0_en_0(x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_en_0),
    .io_in_x255_outbuf_0_rPort_0_backpressure(x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure),
    .io_in_x255_outbuf_0_rPort_0_output_0(x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_output_0),
    .io_in_x450_ready(x522_kernelx522_concrete1_io_in_x450_ready),
    .io_in_x450_valid(x522_kernelx522_concrete1_io_in_x450_valid),
    .io_in_x254_TVALID(x522_kernelx522_concrete1_io_in_x254_TVALID),
    .io_in_x254_TREADY(x522_kernelx522_concrete1_io_in_x254_TREADY),
    .io_in_x254_TDATA(x522_kernelx522_concrete1_io_in_x254_TDATA),
    .io_sigsIn_smEnableOuts_0(x522_kernelx522_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x522_kernelx522_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x522_kernelx522_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x522_kernelx522_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x522_kernelx522_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x522_kernelx522_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x522_kernelx522_concrete1_io_rr)
  );
  assign _T_266 = x522_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32863.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@32902.4 package.scala 96:25:@32903.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32910.4 package.scala 96:25:@32911.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@32913.4]
  assign io_in_x449_valid = x522_kernelx522_concrete1_io_in_x449_valid; // @[sm_x522.scala 63:23:@33015.4]
  assign io_in_x449_bits_wdata_0 = x522_kernelx522_concrete1_io_in_x449_bits_wdata_0; // @[sm_x522.scala 63:23:@33014.4]
  assign io_in_x449_bits_wstrb = x522_kernelx522_concrete1_io_in_x449_bits_wstrb; // @[sm_x522.scala 63:23:@33013.4]
  assign io_in_x448_valid = x522_kernelx522_concrete1_io_in_x448_valid; // @[sm_x522.scala 64:23:@33019.4]
  assign io_in_x448_bits_addr = x522_kernelx522_concrete1_io_in_x448_bits_addr; // @[sm_x522.scala 64:23:@33018.4]
  assign io_in_x448_bits_size = x522_kernelx522_concrete1_io_in_x448_bits_size; // @[sm_x522.scala 64:23:@33017.4]
  assign io_in_x253_TREADY = x522_kernelx522_concrete1_io_in_x253_TREADY; // @[sm_x522.scala 65:23:@33028.4]
  assign io_in_x450_ready = x522_kernelx522_concrete1_io_in_x450_ready; // @[sm_x522.scala 68:23:@33038.4]
  assign io_in_x254_TVALID = x522_kernelx522_concrete1_io_in_x254_TVALID; // @[sm_x522.scala 69:23:@33047.4]
  assign io_in_x254_TDATA = x522_kernelx522_concrete1_io_in_x254_TDATA; // @[sm_x522.scala 69:23:@33045.4]
  assign io_sigsOut_smDoneIn_0 = x522_sm_io_done; // @[SpatialBlocks.scala 156:53:@32920.4]
  assign x255_outbuf_0_clock = clock; // @[:@32773.4]
  assign x255_outbuf_0_reset = reset; // @[:@32774.4]
  assign x255_outbuf_0_io_rPort_0_ofs_0 = x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@33034.4]
  assign x255_outbuf_0_io_rPort_0_en_0 = x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@33033.4]
  assign x255_outbuf_0_io_rPort_0_backpressure = x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@33032.4]
  assign x522_sm_clock = clock; // @[:@32831.4]
  assign x522_sm_reset = reset; // @[:@32832.4]
  assign x522_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@32917.4]
  assign x522_sm_io_ctrDone = x522_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@32867.4]
  assign x522_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@32919.4]
  assign x522_sm_io_doneIn_0 = x522_kernelx522_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@32887.4]
  assign x522_sm_io_doneIn_1 = x522_kernelx522_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@32888.4]
  assign RetimeWrapper_clock = clock; // @[:@32898.4]
  assign RetimeWrapper_reset = reset; // @[:@32899.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32901.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@32900.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32906.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32907.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32909.4]
  assign RetimeWrapper_1_io_in = x522_sm_io_done; // @[package.scala 94:16:@32908.4]
  assign x522_kernelx522_concrete1_clock = clock; // @[:@32935.4]
  assign x522_kernelx522_concrete1_reset = reset; // @[:@32936.4]
  assign x522_kernelx522_concrete1_io_in_x449_ready = io_in_x449_ready; // @[sm_x522.scala 63:23:@33016.4]
  assign x522_kernelx522_concrete1_io_in_x448_ready = io_in_x448_ready; // @[sm_x522.scala 64:23:@33020.4]
  assign x522_kernelx522_concrete1_io_in_x253_TVALID = io_in_x253_TVALID; // @[sm_x522.scala 65:23:@33029.4]
  assign x522_kernelx522_concrete1_io_in_x253_TDATA = io_in_x253_TDATA; // @[sm_x522.scala 65:23:@33027.4]
  assign x522_kernelx522_concrete1_io_in_x253_TID = io_in_x253_TID; // @[sm_x522.scala 65:23:@33023.4]
  assign x522_kernelx522_concrete1_io_in_x253_TDEST = io_in_x253_TDEST; // @[sm_x522.scala 65:23:@33022.4]
  assign x522_kernelx522_concrete1_io_in_x251_outdram_number = io_in_x251_outdram_number; // @[sm_x522.scala 66:31:@33030.4]
  assign x522_kernelx522_concrete1_io_in_x255_outbuf_0_rPort_0_output_0 = x255_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@33031.4]
  assign x522_kernelx522_concrete1_io_in_x450_valid = io_in_x450_valid; // @[sm_x522.scala 68:23:@33037.4]
  assign x522_kernelx522_concrete1_io_in_x254_TREADY = io_in_x254_TREADY; // @[sm_x522.scala 69:23:@33046.4]
  assign x522_kernelx522_concrete1_io_sigsIn_smEnableOuts_0 = x522_sm_io_enableOut_0; // @[sm_x522.scala 107:22:@33058.4]
  assign x522_kernelx522_concrete1_io_sigsIn_smEnableOuts_1 = x522_sm_io_enableOut_1; // @[sm_x522.scala 107:22:@33059.4]
  assign x522_kernelx522_concrete1_io_sigsIn_smChildAcks_0 = x522_sm_io_childAck_0; // @[sm_x522.scala 107:22:@33054.4]
  assign x522_kernelx522_concrete1_io_sigsIn_smChildAcks_1 = x522_sm_io_childAck_1; // @[sm_x522.scala 107:22:@33055.4]
  assign x522_kernelx522_concrete1_io_rr = io_rr; // @[sm_x522.scala 106:18:@33048.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@33081.2]
  input          clock, // @[:@33082.4]
  input          reset, // @[:@33083.4]
  input          io_enable, // @[:@33084.4]
  output         io_done, // @[:@33084.4]
  input          io_reset, // @[:@33084.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@33084.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@33084.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@33084.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@33084.4]
  output         io_memStreams_loads_0_data_ready, // @[:@33084.4]
  input          io_memStreams_loads_0_data_valid, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@33084.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@33084.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@33084.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@33084.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@33084.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@33084.4]
  input          io_memStreams_stores_0_data_ready, // @[:@33084.4]
  output         io_memStreams_stores_0_data_valid, // @[:@33084.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@33084.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@33084.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@33084.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@33084.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@33084.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@33084.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@33084.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@33084.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@33084.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@33084.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@33084.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@33084.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@33084.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@33084.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@33084.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@33084.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@33084.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@33084.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@33084.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@33084.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@33084.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@33084.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@33084.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@33084.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@33084.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@33084.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@33084.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@33084.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@33084.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@33084.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@33084.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@33084.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@33084.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@33084.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@33084.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@33084.4]
  output         io_heap_0_req_valid, // @[:@33084.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@33084.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@33084.4]
  input          io_heap_0_resp_valid, // @[:@33084.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@33084.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@33084.4]
  input  [63:0]  io_argIns_0, // @[:@33084.4]
  input  [63:0]  io_argIns_1, // @[:@33084.4]
  input          io_argOuts_0_port_ready, // @[:@33084.4]
  output         io_argOuts_0_port_valid, // @[:@33084.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@33084.4]
  input  [63:0]  io_argOuts_0_echo // @[:@33084.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@33232.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@33232.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@33232.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@33232.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33250.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33250.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33250.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33250.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33250.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@33259.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@33259.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@33259.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@33259.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@33259.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@33259.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@33298.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33330.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33330.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33330.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33330.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33330.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x449_ready; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x449_valid; // @[sm_RootController.scala 91:24:@33392.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x449_bits_wdata_0; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x449_bits_wstrb; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x448_ready; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x448_valid; // @[sm_RootController.scala 91:24:@33392.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x448_bits_addr; // @[sm_RootController.scala 91:24:@33392.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x448_bits_size; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x253_TVALID; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x253_TREADY; // @[sm_RootController.scala 91:24:@33392.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x253_TDATA; // @[sm_RootController.scala 91:24:@33392.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x253_TID; // @[sm_RootController.scala 91:24:@33392.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x253_TDEST; // @[sm_RootController.scala 91:24:@33392.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x251_outdram_number; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x450_ready; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x450_valid; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x254_TVALID; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_in_x254_TREADY; // @[sm_RootController.scala 91:24:@33392.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x254_TDATA; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@33392.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@33392.4]
  wire  _T_599; // @[package.scala 96:25:@33255.4 package.scala 96:25:@33256.4]
  wire  _T_664; // @[Main.scala 46:50:@33326.4]
  wire  _T_665; // @[Main.scala 46:59:@33327.4]
  wire  _T_677; // @[package.scala 100:49:@33347.4]
  reg  _T_680; // @[package.scala 48:56:@33348.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@33232.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33250.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@33259.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@33298.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33330.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@33392.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x449_ready(RootController_kernelRootController_concrete1_io_in_x449_ready),
    .io_in_x449_valid(RootController_kernelRootController_concrete1_io_in_x449_valid),
    .io_in_x449_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x449_bits_wdata_0),
    .io_in_x449_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x449_bits_wstrb),
    .io_in_x448_ready(RootController_kernelRootController_concrete1_io_in_x448_ready),
    .io_in_x448_valid(RootController_kernelRootController_concrete1_io_in_x448_valid),
    .io_in_x448_bits_addr(RootController_kernelRootController_concrete1_io_in_x448_bits_addr),
    .io_in_x448_bits_size(RootController_kernelRootController_concrete1_io_in_x448_bits_size),
    .io_in_x253_TVALID(RootController_kernelRootController_concrete1_io_in_x253_TVALID),
    .io_in_x253_TREADY(RootController_kernelRootController_concrete1_io_in_x253_TREADY),
    .io_in_x253_TDATA(RootController_kernelRootController_concrete1_io_in_x253_TDATA),
    .io_in_x253_TID(RootController_kernelRootController_concrete1_io_in_x253_TID),
    .io_in_x253_TDEST(RootController_kernelRootController_concrete1_io_in_x253_TDEST),
    .io_in_x251_outdram_number(RootController_kernelRootController_concrete1_io_in_x251_outdram_number),
    .io_in_x450_ready(RootController_kernelRootController_concrete1_io_in_x450_ready),
    .io_in_x450_valid(RootController_kernelRootController_concrete1_io_in_x450_valid),
    .io_in_x254_TVALID(RootController_kernelRootController_concrete1_io_in_x254_TVALID),
    .io_in_x254_TREADY(RootController_kernelRootController_concrete1_io_in_x254_TREADY),
    .io_in_x254_TDATA(RootController_kernelRootController_concrete1_io_in_x254_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@33255.4 package.scala 96:25:@33256.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@33326.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@33327.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33347.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@33346.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x448_valid; // @[sm_RootController.scala 61:23:@33459.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x448_bits_addr; // @[sm_RootController.scala 61:23:@33458.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x448_bits_size; // @[sm_RootController.scala 61:23:@33457.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x449_valid; // @[sm_RootController.scala 60:23:@33455.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x449_bits_wdata_0; // @[sm_RootController.scala 60:23:@33454.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x449_bits_wstrb; // @[sm_RootController.scala 60:23:@33453.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x450_ready; // @[sm_RootController.scala 64:23:@33473.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x253_TREADY; // @[sm_RootController.scala 62:23:@33468.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x254_TVALID; // @[sm_RootController.scala 65:23:@33482.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x254_TDATA; // @[sm_RootController.scala 65:23:@33480.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 65:23:@33479.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 65:23:@33478.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 65:23:@33477.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 65:23:@33476.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 65:23:@33475.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 65:23:@33474.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@33233.4]
  assign SingleCounter_reset = reset; // @[:@33234.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@33248.4]
  assign RetimeWrapper_clock = clock; // @[:@33251.4]
  assign RetimeWrapper_reset = reset; // @[:@33252.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33254.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@33253.4]
  assign SRFF_clock = clock; // @[:@33260.4]
  assign SRFF_reset = reset; // @[:@33261.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@33510.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@33344.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@33345.4]
  assign RootController_sm_clock = clock; // @[:@33299.4]
  assign RootController_sm_reset = reset; // @[:@33300.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@33343.4 SpatialBlocks.scala 140:18:@33377.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@33371.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@33351.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@33339.4 SpatialBlocks.scala 142:21:@33379.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33368.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33331.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33332.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33334.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@33333.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@33393.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@33394.4]
  assign RootController_kernelRootController_concrete1_io_in_x449_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 60:23:@33456.4]
  assign RootController_kernelRootController_concrete1_io_in_x448_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 61:23:@33460.4]
  assign RootController_kernelRootController_concrete1_io_in_x253_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 62:23:@33469.4]
  assign RootController_kernelRootController_concrete1_io_in_x253_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 62:23:@33467.4]
  assign RootController_kernelRootController_concrete1_io_in_x253_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 62:23:@33463.4]
  assign RootController_kernelRootController_concrete1_io_in_x253_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 62:23:@33462.4]
  assign RootController_kernelRootController_concrete1_io_in_x251_outdram_number = io_argIns_1; // @[sm_RootController.scala 63:31:@33470.4]
  assign RootController_kernelRootController_concrete1_io_in_x450_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 64:23:@33472.4]
  assign RootController_kernelRootController_concrete1_io_in_x254_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 65:23:@33481.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@33491.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@33489.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@33483.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@33512.2]
  input        clock, // @[:@33513.4]
  input        reset, // @[:@33514.4]
  input        io_enable, // @[:@33515.4]
  output [5:0] io_out, // @[:@33515.4]
  output [5:0] io_next // @[:@33515.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@33517.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@33518.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@33519.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@33524.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@33518.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@33519.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@33524.6]
  assign io_out = count; // @[Counter.scala 25:10:@33527.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@33528.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_17( // @[:@33564.2]
  input         clock, // @[:@33565.4]
  input         reset, // @[:@33566.4]
  input  [5:0]  io_raddr, // @[:@33567.4]
  input         io_wen, // @[:@33567.4]
  input  [5:0]  io_waddr, // @[:@33567.4]
  input  [63:0] io_wdata_addr, // @[:@33567.4]
  input  [31:0] io_wdata_size, // @[:@33567.4]
  output [63:0] io_rdata_addr, // @[:@33567.4]
  output [31:0] io_rdata_size // @[:@33567.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@33569.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@33569.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@33569.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@33569.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@33569.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@33569.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@33569.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@33569.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@33569.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@33583.4]
  wire  _T_20; // @[SRAM.scala 182:49:@33588.4]
  wire  _T_21; // @[SRAM.scala 182:37:@33589.4]
  reg  _T_24; // @[SRAM.scala 182:29:@33590.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@33593.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@33595.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@33569.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@33583.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@33588.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@33589.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@33595.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@33604.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@33603.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@33584.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@33585.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@33581.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@33587.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@33586.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@33582.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@33580.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@33579.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@33606.2]
  input         clock, // @[:@33607.4]
  input         reset, // @[:@33608.4]
  output        io_in_ready, // @[:@33609.4]
  input         io_in_valid, // @[:@33609.4]
  input  [63:0] io_in_bits_addr, // @[:@33609.4]
  input  [31:0] io_in_bits_size, // @[:@33609.4]
  input         io_out_ready, // @[:@33609.4]
  output        io_out_valid, // @[:@33609.4]
  output [63:0] io_out_bits_addr, // @[:@33609.4]
  output [31:0] io_out_bits_size // @[:@33609.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@34005.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@34005.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@34005.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@34005.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@34005.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@34015.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@34015.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@34015.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@34015.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@34015.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@34030.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@34030.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@34030.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@34030.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@34030.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@34030.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@34030.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@34030.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@34030.4]
  wire  writeEn; // @[FIFO.scala 30:29:@34003.4]
  wire  readEn; // @[FIFO.scala 31:29:@34004.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@34025.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@34026.4]
  wire  _T_824; // @[FIFO.scala 45:27:@34027.4]
  wire  empty; // @[FIFO.scala 45:24:@34028.4]
  wire  full; // @[FIFO.scala 46:23:@34029.4]
  wire  _T_827; // @[FIFO.scala 83:17:@34042.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@34043.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@34005.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@34015.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_17 SRAM ( // @[FIFO.scala 73:19:@34030.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@34003.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@34004.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@34026.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@34027.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@34028.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@34029.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@34042.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@34043.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@34049.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@34047.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@34040.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@34039.4]
  assign enqCounter_clock = clock; // @[:@34006.4]
  assign enqCounter_reset = reset; // @[:@34007.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@34013.4]
  assign deqCounter_clock = clock; // @[:@34016.4]
  assign deqCounter_reset = reset; // @[:@34017.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@34023.4]
  assign SRAM_clock = clock; // @[:@34031.4]
  assign SRAM_reset = reset; // @[:@34032.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@34034.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@34035.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@34036.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@34038.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@34037.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@34051.2]
  input        clock, // @[:@34052.4]
  input        reset, // @[:@34053.4]
  input        io_enable, // @[:@34054.4]
  output [3:0] io_out // @[:@34054.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@34056.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@34057.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@34058.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@34063.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@34057.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@34058.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@34063.6]
  assign io_out = count; // @[Counter.scala 25:10:@34066.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@34087.2]
  input        clock, // @[:@34088.4]
  input        reset, // @[:@34089.4]
  input        io_reset, // @[:@34090.4]
  input        io_enable, // @[:@34090.4]
  input  [1:0] io_stride, // @[:@34090.4]
  output [1:0] io_out, // @[:@34090.4]
  output [1:0] io_next // @[:@34090.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@34092.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@34093.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@34094.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@34099.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@34095.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@34093.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@34094.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@34099.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@34095.4]
  assign io_out = count; // @[Counter.scala 25:10:@34102.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@34103.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_18( // @[:@34139.2]
  input         clock, // @[:@34140.4]
  input         reset, // @[:@34141.4]
  input  [1:0]  io_raddr, // @[:@34142.4]
  input         io_wen, // @[:@34142.4]
  input  [1:0]  io_waddr, // @[:@34142.4]
  input  [31:0] io_wdata, // @[:@34142.4]
  output [31:0] io_rdata, // @[:@34142.4]
  input         io_backpressure // @[:@34142.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@34144.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@34144.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@34144.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@34144.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@34144.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@34144.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@34144.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@34144.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@34144.4]
  wire  _T_19; // @[SRAM.scala 182:49:@34162.4]
  wire  _T_20; // @[SRAM.scala 182:37:@34163.4]
  reg  _T_23; // @[SRAM.scala 182:29:@34164.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@34166.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@34144.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@34162.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@34163.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@34171.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@34158.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@34159.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@34156.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@34161.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@34160.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@34157.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@34155.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@34154.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@34173.2]
  input         clock, // @[:@34174.4]
  input         reset, // @[:@34175.4]
  output        io_in_ready, // @[:@34176.4]
  input         io_in_valid, // @[:@34176.4]
  input  [31:0] io_in_bits, // @[:@34176.4]
  input         io_out_ready, // @[:@34176.4]
  output        io_out_valid, // @[:@34176.4]
  output [31:0] io_out_bits // @[:@34176.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@34202.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@34202.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@34202.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@34202.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@34202.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@34202.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@34202.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@34212.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@34212.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@34212.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@34212.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@34212.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@34212.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@34212.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@34227.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@34227.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@34227.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@34227.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@34227.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@34227.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@34227.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@34227.4]
  wire  writeEn; // @[FIFO.scala 30:29:@34200.4]
  wire  readEn; // @[FIFO.scala 31:29:@34201.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@34222.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@34223.4]
  wire  _T_104; // @[FIFO.scala 45:27:@34224.4]
  wire  empty; // @[FIFO.scala 45:24:@34225.4]
  wire  full; // @[FIFO.scala 46:23:@34226.4]
  wire  _T_107; // @[FIFO.scala 83:17:@34237.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@34238.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@34202.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@34212.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_18 SRAM ( // @[FIFO.scala 73:19:@34227.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@34200.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@34201.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@34223.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@34224.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@34225.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@34226.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@34237.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@34238.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@34244.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@34242.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@34235.4]
  assign enqCounter_clock = clock; // @[:@34203.4]
  assign enqCounter_reset = reset; // @[:@34204.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@34210.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@34211.4]
  assign deqCounter_clock = clock; // @[:@34213.4]
  assign deqCounter_reset = reset; // @[:@34214.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@34220.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@34221.4]
  assign SRAM_clock = clock; // @[:@34228.4]
  assign SRAM_reset = reset; // @[:@34229.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@34231.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@34232.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@34233.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@34234.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@34236.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@36631.2]
  input         clock, // @[:@36632.4]
  input         reset, // @[:@36633.4]
  output        io_in_ready, // @[:@36634.4]
  input         io_in_valid, // @[:@36634.4]
  input  [31:0] io_in_bits_0, // @[:@36634.4]
  input         io_out_ready, // @[:@36634.4]
  output        io_out_valid, // @[:@36634.4]
  output [31:0] io_out_bits_0, // @[:@36634.4]
  output [31:0] io_out_bits_1, // @[:@36634.4]
  output [31:0] io_out_bits_2, // @[:@36634.4]
  output [31:0] io_out_bits_3, // @[:@36634.4]
  output [31:0] io_out_bits_4, // @[:@36634.4]
  output [31:0] io_out_bits_5, // @[:@36634.4]
  output [31:0] io_out_bits_6, // @[:@36634.4]
  output [31:0] io_out_bits_7, // @[:@36634.4]
  output [31:0] io_out_bits_8, // @[:@36634.4]
  output [31:0] io_out_bits_9, // @[:@36634.4]
  output [31:0] io_out_bits_10, // @[:@36634.4]
  output [31:0] io_out_bits_11, // @[:@36634.4]
  output [31:0] io_out_bits_12, // @[:@36634.4]
  output [31:0] io_out_bits_13, // @[:@36634.4]
  output [31:0] io_out_bits_14, // @[:@36634.4]
  output [31:0] io_out_bits_15 // @[:@36634.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@36638.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@36638.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@36638.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@36638.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@36649.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@36649.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@36649.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@36649.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@36662.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@36662.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@36662.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@36662.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@36662.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@36662.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@36662.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@36662.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@36697.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@36697.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@36697.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@36697.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@36697.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@36697.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@36697.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@36697.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@36732.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@36732.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@36732.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@36732.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@36732.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@36732.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@36732.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@36732.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@36767.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@36767.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@36767.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@36767.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@36767.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@36767.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@36767.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@36767.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@36802.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@36802.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@36802.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@36802.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@36802.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@36802.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@36802.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@36802.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@36837.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@36837.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@36837.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@36837.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@36837.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@36837.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@36837.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@36837.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@36872.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@36872.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@36872.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@36872.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@36872.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@36872.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@36872.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@36872.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@36907.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@36907.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@36907.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@36907.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@36907.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@36907.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@36907.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@36907.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@36942.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@36942.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@36942.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@36942.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@36942.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@36942.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@36942.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@36942.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@36977.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@36977.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@36977.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@36977.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@36977.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@36977.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@36977.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@36977.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@37012.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@37012.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@37012.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@37012.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@37012.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@37012.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@37012.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@37012.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@37047.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@37047.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@37047.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@37047.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@37047.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@37047.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@37047.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@37047.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@37082.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@37082.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@37082.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@37082.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@37082.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@37082.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@37082.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@37082.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@37117.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@37117.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@37117.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@37117.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@37117.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@37117.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@37117.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@37117.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@37152.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@37152.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@37152.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@37152.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@37152.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@37152.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@37152.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@37152.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@37187.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@37187.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@37187.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@37187.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@37187.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@37187.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@37187.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@37187.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@36637.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@36660.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@36687.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@36722.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@36757.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@36792.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@36827.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@36862.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@36897.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@36932.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@36967.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@37002.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@37037.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@37072.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@37107.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@37142.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@37177.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@37212.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37223.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37224.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37225.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37226.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37227.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37228.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37229.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37230.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37231.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37232.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37233.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37234.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37235.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37236.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37237.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@37254.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37238.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@37273.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@37274.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@37275.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@37276.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@37277.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@37278.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@37279.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@37280.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@37281.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@37282.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@37283.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@37284.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@37285.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@37286.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@36638.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@36649.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@36662.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@36697.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@36732.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@36767.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@36802.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@36837.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@36872.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@36907.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@36942.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@36977.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@37012.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@37047.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@37082.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@37117.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@37152.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@37187.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@36637.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@36660.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@36687.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@36722.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@36757.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@36792.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@36827.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@36862.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@36897.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@36932.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@36967.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@37002.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@37037.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@37072.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@37107.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@37142.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@37177.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@37212.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37223.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37224.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37225.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37226.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37227.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37228.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37229.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37230.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37231.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37232.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37233.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37234.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37235.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37236.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37237.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@37254.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@37222.4 FIFOVec.scala 49:42:@37238.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@37273.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@37274.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@37275.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@37276.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@37277.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@37278.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@37279.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@37280.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@37281.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@37282.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@37283.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@37284.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@37285.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@37286.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@37255.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@37289.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@37597.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@37598.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@37599.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@37600.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@37601.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@37602.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@37603.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@37604.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@37605.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@37606.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@37607.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@37608.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@37609.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@37610.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@37611.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@37612.4]
  assign enqCounter_clock = clock; // @[:@36639.4]
  assign enqCounter_reset = reset; // @[:@36640.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@36647.4]
  assign deqCounter_clock = clock; // @[:@36650.4]
  assign deqCounter_reset = reset; // @[:@36651.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@36658.4]
  assign fifos_0_clock = clock; // @[:@36663.4]
  assign fifos_0_reset = reset; // @[:@36664.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@36690.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36692.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36696.4]
  assign fifos_1_clock = clock; // @[:@36698.4]
  assign fifos_1_reset = reset; // @[:@36699.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@36725.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36727.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36731.4]
  assign fifos_2_clock = clock; // @[:@36733.4]
  assign fifos_2_reset = reset; // @[:@36734.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@36760.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36762.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36766.4]
  assign fifos_3_clock = clock; // @[:@36768.4]
  assign fifos_3_reset = reset; // @[:@36769.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@36795.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36797.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36801.4]
  assign fifos_4_clock = clock; // @[:@36803.4]
  assign fifos_4_reset = reset; // @[:@36804.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@36830.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36832.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36836.4]
  assign fifos_5_clock = clock; // @[:@36838.4]
  assign fifos_5_reset = reset; // @[:@36839.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@36865.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36867.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36871.4]
  assign fifos_6_clock = clock; // @[:@36873.4]
  assign fifos_6_reset = reset; // @[:@36874.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@36900.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36902.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36906.4]
  assign fifos_7_clock = clock; // @[:@36908.4]
  assign fifos_7_reset = reset; // @[:@36909.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@36935.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36937.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36941.4]
  assign fifos_8_clock = clock; // @[:@36943.4]
  assign fifos_8_reset = reset; // @[:@36944.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@36970.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36972.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36976.4]
  assign fifos_9_clock = clock; // @[:@36978.4]
  assign fifos_9_reset = reset; // @[:@36979.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@37005.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37007.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37011.4]
  assign fifos_10_clock = clock; // @[:@37013.4]
  assign fifos_10_reset = reset; // @[:@37014.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@37040.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37042.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37046.4]
  assign fifos_11_clock = clock; // @[:@37048.4]
  assign fifos_11_reset = reset; // @[:@37049.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@37075.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37077.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37081.4]
  assign fifos_12_clock = clock; // @[:@37083.4]
  assign fifos_12_reset = reset; // @[:@37084.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@37110.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37112.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37116.4]
  assign fifos_13_clock = clock; // @[:@37118.4]
  assign fifos_13_reset = reset; // @[:@37119.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@37145.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37147.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37151.4]
  assign fifos_14_clock = clock; // @[:@37153.4]
  assign fifos_14_reset = reset; // @[:@37154.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@37180.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37182.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37186.4]
  assign fifos_15_clock = clock; // @[:@37188.4]
  assign fifos_15_reset = reset; // @[:@37189.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@37215.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37217.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37221.4]
endmodule
module FFRAM( // @[:@37686.2]
  input        clock, // @[:@37687.4]
  input        reset, // @[:@37688.4]
  input  [1:0] io_raddr, // @[:@37689.4]
  input        io_wen, // @[:@37689.4]
  input  [1:0] io_waddr, // @[:@37689.4]
  input        io_wdata, // @[:@37689.4]
  output       io_rdata, // @[:@37689.4]
  input        io_banks_0_wdata_valid, // @[:@37689.4]
  input        io_banks_0_wdata_bits, // @[:@37689.4]
  input        io_banks_1_wdata_valid, // @[:@37689.4]
  input        io_banks_1_wdata_bits, // @[:@37689.4]
  input        io_banks_2_wdata_valid, // @[:@37689.4]
  input        io_banks_2_wdata_bits, // @[:@37689.4]
  input        io_banks_3_wdata_valid, // @[:@37689.4]
  input        io_banks_3_wdata_bits // @[:@37689.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@37693.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@37694.4]
  wire  _T_89; // @[SRAM.scala 148:25:@37695.4]
  wire  _T_90; // @[SRAM.scala 148:15:@37696.4]
  wire  _T_91; // @[SRAM.scala 149:15:@37698.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@37697.4]
  reg  regs_1; // @[SRAM.scala 145:20:@37704.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@37705.4]
  wire  _T_98; // @[SRAM.scala 148:25:@37706.4]
  wire  _T_99; // @[SRAM.scala 148:15:@37707.4]
  wire  _T_100; // @[SRAM.scala 149:15:@37709.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@37708.4]
  reg  regs_2; // @[SRAM.scala 145:20:@37715.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@37716.4]
  wire  _T_107; // @[SRAM.scala 148:25:@37717.4]
  wire  _T_108; // @[SRAM.scala 148:15:@37718.4]
  wire  _T_109; // @[SRAM.scala 149:15:@37720.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@37719.4]
  reg  regs_3; // @[SRAM.scala 145:20:@37726.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@37727.4]
  wire  _T_116; // @[SRAM.scala 148:25:@37728.4]
  wire  _T_117; // @[SRAM.scala 148:15:@37729.4]
  wire  _T_118; // @[SRAM.scala 149:15:@37731.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@37730.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@37740.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@37740.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@37694.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@37695.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@37696.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@37698.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@37697.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@37705.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@37706.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@37707.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@37709.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@37708.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@37716.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@37717.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@37718.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@37720.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@37719.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@37727.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@37728.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@37729.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@37731.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@37730.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@37740.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@37740.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@37740.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@37742.2]
  input   clock, // @[:@37743.4]
  input   reset, // @[:@37744.4]
  output  io_in_ready, // @[:@37745.4]
  input   io_in_valid, // @[:@37745.4]
  input   io_in_bits, // @[:@37745.4]
  input   io_out_ready, // @[:@37745.4]
  output  io_out_valid, // @[:@37745.4]
  output  io_out_bits // @[:@37745.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@37771.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@37771.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@37771.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@37771.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@37771.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@37771.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@37771.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@37781.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@37781.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@37781.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@37781.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@37781.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@37781.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@37781.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@37796.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@37796.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@37796.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@37796.4]
  wire  writeEn; // @[FIFO.scala 30:29:@37769.4]
  wire  readEn; // @[FIFO.scala 31:29:@37770.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@37791.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@37792.4]
  wire  _T_104; // @[FIFO.scala 45:27:@37793.4]
  wire  empty; // @[FIFO.scala 45:24:@37794.4]
  wire  full; // @[FIFO.scala 46:23:@37795.4]
  wire  _T_157; // @[FIFO.scala 83:17:@37882.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@37883.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@37771.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@37781.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@37796.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@37769.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@37770.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@37792.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@37793.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@37794.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@37795.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@37882.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@37883.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@37889.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@37887.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@37821.4]
  assign enqCounter_clock = clock; // @[:@37772.4]
  assign enqCounter_reset = reset; // @[:@37773.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@37779.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@37780.4]
  assign deqCounter_clock = clock; // @[:@37782.4]
  assign deqCounter_reset = reset; // @[:@37783.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@37789.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@37790.4]
  assign FFRAM_clock = clock; // @[:@37797.4]
  assign FFRAM_reset = reset; // @[:@37798.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@37817.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@37818.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@37819.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@37820.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@37823.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@37822.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@37826.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@37825.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@37829.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@37828.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@37832.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@37831.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@41506.2]
  input   clock, // @[:@41507.4]
  input   reset, // @[:@41508.4]
  output  io_in_ready, // @[:@41509.4]
  input   io_in_valid, // @[:@41509.4]
  input   io_in_bits_0, // @[:@41509.4]
  input   io_out_ready, // @[:@41509.4]
  output  io_out_valid, // @[:@41509.4]
  output  io_out_bits_0, // @[:@41509.4]
  output  io_out_bits_1, // @[:@41509.4]
  output  io_out_bits_2, // @[:@41509.4]
  output  io_out_bits_3, // @[:@41509.4]
  output  io_out_bits_4, // @[:@41509.4]
  output  io_out_bits_5, // @[:@41509.4]
  output  io_out_bits_6, // @[:@41509.4]
  output  io_out_bits_7, // @[:@41509.4]
  output  io_out_bits_8, // @[:@41509.4]
  output  io_out_bits_9, // @[:@41509.4]
  output  io_out_bits_10, // @[:@41509.4]
  output  io_out_bits_11, // @[:@41509.4]
  output  io_out_bits_12, // @[:@41509.4]
  output  io_out_bits_13, // @[:@41509.4]
  output  io_out_bits_14, // @[:@41509.4]
  output  io_out_bits_15 // @[:@41509.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@41513.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@41513.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@41513.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@41513.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@41524.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@41524.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@41524.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@41524.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@41537.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@41572.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@41607.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@41642.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@41677.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@41712.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@41747.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@41782.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@41817.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@41852.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@41887.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@41922.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@41957.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@41992.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@42027.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@42062.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@42062.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@41512.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@41535.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@41562.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@41597.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@41632.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@41667.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@41702.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@41737.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@41772.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@41807.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@41842.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@41877.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@41912.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@41947.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@41982.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@42017.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@42052.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@42087.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42098.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42099.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42100.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42101.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42102.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42103.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42104.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42105.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42106.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42107.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42108.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42109.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42110.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42111.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42112.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@42129.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42113.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@42148.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@42149.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@42150.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@42151.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@42152.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@42153.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@42154.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@42155.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@42156.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@42157.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@42158.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@42159.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@42160.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@42161.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@41513.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@41524.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@41537.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@41572.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@41607.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@41642.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@41677.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@41712.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@41747.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@41782.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@41817.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@41852.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@41887.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@41922.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@41957.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@41992.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@42027.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@42062.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@41512.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@41535.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@41562.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@41597.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@41632.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@41667.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@41702.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@41737.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@41772.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@41807.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@41842.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@41877.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@41912.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@41947.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@41982.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@42017.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@42052.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@42087.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42098.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42099.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42100.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42101.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42102.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42103.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42104.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42105.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42106.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42107.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42108.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42109.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42110.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42111.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42112.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@42129.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@42097.4 FIFOVec.scala 49:42:@42113.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@42148.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@42149.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@42150.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@42151.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@42152.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@42153.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@42154.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@42155.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@42156.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@42157.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@42158.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@42159.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@42160.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@42161.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@42130.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@42164.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@42472.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@42473.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@42474.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@42475.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@42476.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@42477.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@42478.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@42479.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@42480.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@42481.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@42482.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@42483.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@42484.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@42485.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@42486.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@42487.4]
  assign enqCounter_clock = clock; // @[:@41514.4]
  assign enqCounter_reset = reset; // @[:@41515.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@41522.4]
  assign deqCounter_clock = clock; // @[:@41525.4]
  assign deqCounter_reset = reset; // @[:@41526.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@41533.4]
  assign fifos_0_clock = clock; // @[:@41538.4]
  assign fifos_0_reset = reset; // @[:@41539.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@41565.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41567.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41571.4]
  assign fifos_1_clock = clock; // @[:@41573.4]
  assign fifos_1_reset = reset; // @[:@41574.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@41600.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41602.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41606.4]
  assign fifos_2_clock = clock; // @[:@41608.4]
  assign fifos_2_reset = reset; // @[:@41609.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@41635.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41637.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41641.4]
  assign fifos_3_clock = clock; // @[:@41643.4]
  assign fifos_3_reset = reset; // @[:@41644.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@41670.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41672.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41676.4]
  assign fifos_4_clock = clock; // @[:@41678.4]
  assign fifos_4_reset = reset; // @[:@41679.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@41705.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41707.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41711.4]
  assign fifos_5_clock = clock; // @[:@41713.4]
  assign fifos_5_reset = reset; // @[:@41714.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@41740.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41742.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41746.4]
  assign fifos_6_clock = clock; // @[:@41748.4]
  assign fifos_6_reset = reset; // @[:@41749.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@41775.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41777.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41781.4]
  assign fifos_7_clock = clock; // @[:@41783.4]
  assign fifos_7_reset = reset; // @[:@41784.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@41810.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41812.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41816.4]
  assign fifos_8_clock = clock; // @[:@41818.4]
  assign fifos_8_reset = reset; // @[:@41819.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@41845.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41847.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41851.4]
  assign fifos_9_clock = clock; // @[:@41853.4]
  assign fifos_9_reset = reset; // @[:@41854.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@41880.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41882.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41886.4]
  assign fifos_10_clock = clock; // @[:@41888.4]
  assign fifos_10_reset = reset; // @[:@41889.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@41915.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41917.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41921.4]
  assign fifos_11_clock = clock; // @[:@41923.4]
  assign fifos_11_reset = reset; // @[:@41924.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@41950.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41952.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41956.4]
  assign fifos_12_clock = clock; // @[:@41958.4]
  assign fifos_12_reset = reset; // @[:@41959.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@41985.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41987.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41991.4]
  assign fifos_13_clock = clock; // @[:@41993.4]
  assign fifos_13_reset = reset; // @[:@41994.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@42020.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42022.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42026.4]
  assign fifos_14_clock = clock; // @[:@42028.4]
  assign fifos_14_reset = reset; // @[:@42029.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@42055.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42057.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42061.4]
  assign fifos_15_clock = clock; // @[:@42063.4]
  assign fifos_15_reset = reset; // @[:@42064.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@42090.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42092.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42096.4]
endmodule
module FIFOWidthConvert( // @[:@42489.2]
  input         clock, // @[:@42490.4]
  input         reset, // @[:@42491.4]
  output        io_in_ready, // @[:@42492.4]
  input         io_in_valid, // @[:@42492.4]
  input  [31:0] io_in_bits_data_0, // @[:@42492.4]
  input         io_in_bits_strobe, // @[:@42492.4]
  input         io_out_ready, // @[:@42492.4]
  output        io_out_valid, // @[:@42492.4]
  output [31:0] io_out_bits_data_0, // @[:@42492.4]
  output [31:0] io_out_bits_data_1, // @[:@42492.4]
  output [31:0] io_out_bits_data_2, // @[:@42492.4]
  output [31:0] io_out_bits_data_3, // @[:@42492.4]
  output [31:0] io_out_bits_data_4, // @[:@42492.4]
  output [31:0] io_out_bits_data_5, // @[:@42492.4]
  output [31:0] io_out_bits_data_6, // @[:@42492.4]
  output [31:0] io_out_bits_data_7, // @[:@42492.4]
  output [31:0] io_out_bits_data_8, // @[:@42492.4]
  output [31:0] io_out_bits_data_9, // @[:@42492.4]
  output [31:0] io_out_bits_data_10, // @[:@42492.4]
  output [31:0] io_out_bits_data_11, // @[:@42492.4]
  output [31:0] io_out_bits_data_12, // @[:@42492.4]
  output [31:0] io_out_bits_data_13, // @[:@42492.4]
  output [31:0] io_out_bits_data_14, // @[:@42492.4]
  output [31:0] io_out_bits_data_15, // @[:@42492.4]
  output [63:0] io_out_bits_strobe // @[:@42492.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@42494.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@42535.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@42594.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@42600.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@42658.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@42664.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@42665.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@42669.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@42673.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@42677.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@42681.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@42685.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@42689.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@42693.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@42697.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@42701.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@42705.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@42709.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@42713.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@42717.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@42721.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@42725.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@42802.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@42811.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@42820.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@42829.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@42838.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@42847.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@42855.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@42494.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@42535.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@42594.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@42600.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@42658.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@42664.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@42665.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@42669.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@42673.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@42677.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@42681.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@42685.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@42689.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@42693.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@42697.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@42701.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@42705.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@42709.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@42713.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@42717.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@42721.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@42725.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@42802.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@42811.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@42820.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@42829.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@42838.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@42847.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@42855.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@42584.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@42585.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@42634.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@42635.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@42636.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@42637.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@42638.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@42639.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@42640.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@42641.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@42642.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@42643.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@42644.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@42645.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@42646.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@42647.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@42648.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@42649.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@42857.4]
  assign FIFOVec_clock = clock; // @[:@42495.4]
  assign FIFOVec_reset = reset; // @[:@42496.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@42581.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@42580.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@42858.4]
  assign FIFOVec_1_clock = clock; // @[:@42536.4]
  assign FIFOVec_1_reset = reset; // @[:@42537.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@42583.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@42582.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@42859.4]
endmodule
module FFRAM_16( // @[:@42897.2]
  input        clock, // @[:@42898.4]
  input        reset, // @[:@42899.4]
  input  [5:0] io_raddr, // @[:@42900.4]
  input        io_wen, // @[:@42900.4]
  input  [5:0] io_waddr, // @[:@42900.4]
  input        io_wdata, // @[:@42900.4]
  output       io_rdata, // @[:@42900.4]
  input        io_banks_0_wdata_valid, // @[:@42900.4]
  input        io_banks_0_wdata_bits, // @[:@42900.4]
  input        io_banks_1_wdata_valid, // @[:@42900.4]
  input        io_banks_1_wdata_bits, // @[:@42900.4]
  input        io_banks_2_wdata_valid, // @[:@42900.4]
  input        io_banks_2_wdata_bits, // @[:@42900.4]
  input        io_banks_3_wdata_valid, // @[:@42900.4]
  input        io_banks_3_wdata_bits, // @[:@42900.4]
  input        io_banks_4_wdata_valid, // @[:@42900.4]
  input        io_banks_4_wdata_bits, // @[:@42900.4]
  input        io_banks_5_wdata_valid, // @[:@42900.4]
  input        io_banks_5_wdata_bits, // @[:@42900.4]
  input        io_banks_6_wdata_valid, // @[:@42900.4]
  input        io_banks_6_wdata_bits, // @[:@42900.4]
  input        io_banks_7_wdata_valid, // @[:@42900.4]
  input        io_banks_7_wdata_bits, // @[:@42900.4]
  input        io_banks_8_wdata_valid, // @[:@42900.4]
  input        io_banks_8_wdata_bits, // @[:@42900.4]
  input        io_banks_9_wdata_valid, // @[:@42900.4]
  input        io_banks_9_wdata_bits, // @[:@42900.4]
  input        io_banks_10_wdata_valid, // @[:@42900.4]
  input        io_banks_10_wdata_bits, // @[:@42900.4]
  input        io_banks_11_wdata_valid, // @[:@42900.4]
  input        io_banks_11_wdata_bits, // @[:@42900.4]
  input        io_banks_12_wdata_valid, // @[:@42900.4]
  input        io_banks_12_wdata_bits, // @[:@42900.4]
  input        io_banks_13_wdata_valid, // @[:@42900.4]
  input        io_banks_13_wdata_bits, // @[:@42900.4]
  input        io_banks_14_wdata_valid, // @[:@42900.4]
  input        io_banks_14_wdata_bits, // @[:@42900.4]
  input        io_banks_15_wdata_valid, // @[:@42900.4]
  input        io_banks_15_wdata_bits, // @[:@42900.4]
  input        io_banks_16_wdata_valid, // @[:@42900.4]
  input        io_banks_16_wdata_bits, // @[:@42900.4]
  input        io_banks_17_wdata_valid, // @[:@42900.4]
  input        io_banks_17_wdata_bits, // @[:@42900.4]
  input        io_banks_18_wdata_valid, // @[:@42900.4]
  input        io_banks_18_wdata_bits, // @[:@42900.4]
  input        io_banks_19_wdata_valid, // @[:@42900.4]
  input        io_banks_19_wdata_bits, // @[:@42900.4]
  input        io_banks_20_wdata_valid, // @[:@42900.4]
  input        io_banks_20_wdata_bits, // @[:@42900.4]
  input        io_banks_21_wdata_valid, // @[:@42900.4]
  input        io_banks_21_wdata_bits, // @[:@42900.4]
  input        io_banks_22_wdata_valid, // @[:@42900.4]
  input        io_banks_22_wdata_bits, // @[:@42900.4]
  input        io_banks_23_wdata_valid, // @[:@42900.4]
  input        io_banks_23_wdata_bits, // @[:@42900.4]
  input        io_banks_24_wdata_valid, // @[:@42900.4]
  input        io_banks_24_wdata_bits, // @[:@42900.4]
  input        io_banks_25_wdata_valid, // @[:@42900.4]
  input        io_banks_25_wdata_bits, // @[:@42900.4]
  input        io_banks_26_wdata_valid, // @[:@42900.4]
  input        io_banks_26_wdata_bits, // @[:@42900.4]
  input        io_banks_27_wdata_valid, // @[:@42900.4]
  input        io_banks_27_wdata_bits, // @[:@42900.4]
  input        io_banks_28_wdata_valid, // @[:@42900.4]
  input        io_banks_28_wdata_bits, // @[:@42900.4]
  input        io_banks_29_wdata_valid, // @[:@42900.4]
  input        io_banks_29_wdata_bits, // @[:@42900.4]
  input        io_banks_30_wdata_valid, // @[:@42900.4]
  input        io_banks_30_wdata_bits, // @[:@42900.4]
  input        io_banks_31_wdata_valid, // @[:@42900.4]
  input        io_banks_31_wdata_bits, // @[:@42900.4]
  input        io_banks_32_wdata_valid, // @[:@42900.4]
  input        io_banks_32_wdata_bits, // @[:@42900.4]
  input        io_banks_33_wdata_valid, // @[:@42900.4]
  input        io_banks_33_wdata_bits, // @[:@42900.4]
  input        io_banks_34_wdata_valid, // @[:@42900.4]
  input        io_banks_34_wdata_bits, // @[:@42900.4]
  input        io_banks_35_wdata_valid, // @[:@42900.4]
  input        io_banks_35_wdata_bits, // @[:@42900.4]
  input        io_banks_36_wdata_valid, // @[:@42900.4]
  input        io_banks_36_wdata_bits, // @[:@42900.4]
  input        io_banks_37_wdata_valid, // @[:@42900.4]
  input        io_banks_37_wdata_bits, // @[:@42900.4]
  input        io_banks_38_wdata_valid, // @[:@42900.4]
  input        io_banks_38_wdata_bits, // @[:@42900.4]
  input        io_banks_39_wdata_valid, // @[:@42900.4]
  input        io_banks_39_wdata_bits, // @[:@42900.4]
  input        io_banks_40_wdata_valid, // @[:@42900.4]
  input        io_banks_40_wdata_bits, // @[:@42900.4]
  input        io_banks_41_wdata_valid, // @[:@42900.4]
  input        io_banks_41_wdata_bits, // @[:@42900.4]
  input        io_banks_42_wdata_valid, // @[:@42900.4]
  input        io_banks_42_wdata_bits, // @[:@42900.4]
  input        io_banks_43_wdata_valid, // @[:@42900.4]
  input        io_banks_43_wdata_bits, // @[:@42900.4]
  input        io_banks_44_wdata_valid, // @[:@42900.4]
  input        io_banks_44_wdata_bits, // @[:@42900.4]
  input        io_banks_45_wdata_valid, // @[:@42900.4]
  input        io_banks_45_wdata_bits, // @[:@42900.4]
  input        io_banks_46_wdata_valid, // @[:@42900.4]
  input        io_banks_46_wdata_bits, // @[:@42900.4]
  input        io_banks_47_wdata_valid, // @[:@42900.4]
  input        io_banks_47_wdata_bits, // @[:@42900.4]
  input        io_banks_48_wdata_valid, // @[:@42900.4]
  input        io_banks_48_wdata_bits, // @[:@42900.4]
  input        io_banks_49_wdata_valid, // @[:@42900.4]
  input        io_banks_49_wdata_bits, // @[:@42900.4]
  input        io_banks_50_wdata_valid, // @[:@42900.4]
  input        io_banks_50_wdata_bits, // @[:@42900.4]
  input        io_banks_51_wdata_valid, // @[:@42900.4]
  input        io_banks_51_wdata_bits, // @[:@42900.4]
  input        io_banks_52_wdata_valid, // @[:@42900.4]
  input        io_banks_52_wdata_bits, // @[:@42900.4]
  input        io_banks_53_wdata_valid, // @[:@42900.4]
  input        io_banks_53_wdata_bits, // @[:@42900.4]
  input        io_banks_54_wdata_valid, // @[:@42900.4]
  input        io_banks_54_wdata_bits, // @[:@42900.4]
  input        io_banks_55_wdata_valid, // @[:@42900.4]
  input        io_banks_55_wdata_bits, // @[:@42900.4]
  input        io_banks_56_wdata_valid, // @[:@42900.4]
  input        io_banks_56_wdata_bits, // @[:@42900.4]
  input        io_banks_57_wdata_valid, // @[:@42900.4]
  input        io_banks_57_wdata_bits, // @[:@42900.4]
  input        io_banks_58_wdata_valid, // @[:@42900.4]
  input        io_banks_58_wdata_bits, // @[:@42900.4]
  input        io_banks_59_wdata_valid, // @[:@42900.4]
  input        io_banks_59_wdata_bits, // @[:@42900.4]
  input        io_banks_60_wdata_valid, // @[:@42900.4]
  input        io_banks_60_wdata_bits, // @[:@42900.4]
  input        io_banks_61_wdata_valid, // @[:@42900.4]
  input        io_banks_61_wdata_bits, // @[:@42900.4]
  input        io_banks_62_wdata_valid, // @[:@42900.4]
  input        io_banks_62_wdata_bits, // @[:@42900.4]
  input        io_banks_63_wdata_valid, // @[:@42900.4]
  input        io_banks_63_wdata_bits // @[:@42900.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@42904.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@42905.4]
  wire  _T_689; // @[SRAM.scala 148:25:@42906.4]
  wire  _T_690; // @[SRAM.scala 148:15:@42907.4]
  wire  _T_691; // @[SRAM.scala 149:15:@42909.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@42908.4]
  reg  regs_1; // @[SRAM.scala 145:20:@42915.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@42916.4]
  wire  _T_698; // @[SRAM.scala 148:25:@42917.4]
  wire  _T_699; // @[SRAM.scala 148:15:@42918.4]
  wire  _T_700; // @[SRAM.scala 149:15:@42920.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@42919.4]
  reg  regs_2; // @[SRAM.scala 145:20:@42926.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@42927.4]
  wire  _T_707; // @[SRAM.scala 148:25:@42928.4]
  wire  _T_708; // @[SRAM.scala 148:15:@42929.4]
  wire  _T_709; // @[SRAM.scala 149:15:@42931.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@42930.4]
  reg  regs_3; // @[SRAM.scala 145:20:@42937.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@42938.4]
  wire  _T_716; // @[SRAM.scala 148:25:@42939.4]
  wire  _T_717; // @[SRAM.scala 148:15:@42940.4]
  wire  _T_718; // @[SRAM.scala 149:15:@42942.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@42941.4]
  reg  regs_4; // @[SRAM.scala 145:20:@42948.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@42949.4]
  wire  _T_725; // @[SRAM.scala 148:25:@42950.4]
  wire  _T_726; // @[SRAM.scala 148:15:@42951.4]
  wire  _T_727; // @[SRAM.scala 149:15:@42953.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@42952.4]
  reg  regs_5; // @[SRAM.scala 145:20:@42959.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@42960.4]
  wire  _T_734; // @[SRAM.scala 148:25:@42961.4]
  wire  _T_735; // @[SRAM.scala 148:15:@42962.4]
  wire  _T_736; // @[SRAM.scala 149:15:@42964.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@42963.4]
  reg  regs_6; // @[SRAM.scala 145:20:@42970.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@42971.4]
  wire  _T_743; // @[SRAM.scala 148:25:@42972.4]
  wire  _T_744; // @[SRAM.scala 148:15:@42973.4]
  wire  _T_745; // @[SRAM.scala 149:15:@42975.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@42974.4]
  reg  regs_7; // @[SRAM.scala 145:20:@42981.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@42982.4]
  wire  _T_752; // @[SRAM.scala 148:25:@42983.4]
  wire  _T_753; // @[SRAM.scala 148:15:@42984.4]
  wire  _T_754; // @[SRAM.scala 149:15:@42986.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@42985.4]
  reg  regs_8; // @[SRAM.scala 145:20:@42992.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@42993.4]
  wire  _T_761; // @[SRAM.scala 148:25:@42994.4]
  wire  _T_762; // @[SRAM.scala 148:15:@42995.4]
  wire  _T_763; // @[SRAM.scala 149:15:@42997.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@42996.4]
  reg  regs_9; // @[SRAM.scala 145:20:@43003.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@43004.4]
  wire  _T_770; // @[SRAM.scala 148:25:@43005.4]
  wire  _T_771; // @[SRAM.scala 148:15:@43006.4]
  wire  _T_772; // @[SRAM.scala 149:15:@43008.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@43007.4]
  reg  regs_10; // @[SRAM.scala 145:20:@43014.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@43015.4]
  wire  _T_779; // @[SRAM.scala 148:25:@43016.4]
  wire  _T_780; // @[SRAM.scala 148:15:@43017.4]
  wire  _T_781; // @[SRAM.scala 149:15:@43019.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@43018.4]
  reg  regs_11; // @[SRAM.scala 145:20:@43025.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@43026.4]
  wire  _T_788; // @[SRAM.scala 148:25:@43027.4]
  wire  _T_789; // @[SRAM.scala 148:15:@43028.4]
  wire  _T_790; // @[SRAM.scala 149:15:@43030.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@43029.4]
  reg  regs_12; // @[SRAM.scala 145:20:@43036.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@43037.4]
  wire  _T_797; // @[SRAM.scala 148:25:@43038.4]
  wire  _T_798; // @[SRAM.scala 148:15:@43039.4]
  wire  _T_799; // @[SRAM.scala 149:15:@43041.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@43040.4]
  reg  regs_13; // @[SRAM.scala 145:20:@43047.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@43048.4]
  wire  _T_806; // @[SRAM.scala 148:25:@43049.4]
  wire  _T_807; // @[SRAM.scala 148:15:@43050.4]
  wire  _T_808; // @[SRAM.scala 149:15:@43052.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@43051.4]
  reg  regs_14; // @[SRAM.scala 145:20:@43058.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@43059.4]
  wire  _T_815; // @[SRAM.scala 148:25:@43060.4]
  wire  _T_816; // @[SRAM.scala 148:15:@43061.4]
  wire  _T_817; // @[SRAM.scala 149:15:@43063.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@43062.4]
  reg  regs_15; // @[SRAM.scala 145:20:@43069.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@43070.4]
  wire  _T_824; // @[SRAM.scala 148:25:@43071.4]
  wire  _T_825; // @[SRAM.scala 148:15:@43072.4]
  wire  _T_826; // @[SRAM.scala 149:15:@43074.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@43073.4]
  reg  regs_16; // @[SRAM.scala 145:20:@43080.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@43081.4]
  wire  _T_833; // @[SRAM.scala 148:25:@43082.4]
  wire  _T_834; // @[SRAM.scala 148:15:@43083.4]
  wire  _T_835; // @[SRAM.scala 149:15:@43085.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@43084.4]
  reg  regs_17; // @[SRAM.scala 145:20:@43091.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@43092.4]
  wire  _T_842; // @[SRAM.scala 148:25:@43093.4]
  wire  _T_843; // @[SRAM.scala 148:15:@43094.4]
  wire  _T_844; // @[SRAM.scala 149:15:@43096.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@43095.4]
  reg  regs_18; // @[SRAM.scala 145:20:@43102.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@43103.4]
  wire  _T_851; // @[SRAM.scala 148:25:@43104.4]
  wire  _T_852; // @[SRAM.scala 148:15:@43105.4]
  wire  _T_853; // @[SRAM.scala 149:15:@43107.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@43106.4]
  reg  regs_19; // @[SRAM.scala 145:20:@43113.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@43114.4]
  wire  _T_860; // @[SRAM.scala 148:25:@43115.4]
  wire  _T_861; // @[SRAM.scala 148:15:@43116.4]
  wire  _T_862; // @[SRAM.scala 149:15:@43118.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@43117.4]
  reg  regs_20; // @[SRAM.scala 145:20:@43124.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@43125.4]
  wire  _T_869; // @[SRAM.scala 148:25:@43126.4]
  wire  _T_870; // @[SRAM.scala 148:15:@43127.4]
  wire  _T_871; // @[SRAM.scala 149:15:@43129.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@43128.4]
  reg  regs_21; // @[SRAM.scala 145:20:@43135.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@43136.4]
  wire  _T_878; // @[SRAM.scala 148:25:@43137.4]
  wire  _T_879; // @[SRAM.scala 148:15:@43138.4]
  wire  _T_880; // @[SRAM.scala 149:15:@43140.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@43139.4]
  reg  regs_22; // @[SRAM.scala 145:20:@43146.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@43147.4]
  wire  _T_887; // @[SRAM.scala 148:25:@43148.4]
  wire  _T_888; // @[SRAM.scala 148:15:@43149.4]
  wire  _T_889; // @[SRAM.scala 149:15:@43151.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@43150.4]
  reg  regs_23; // @[SRAM.scala 145:20:@43157.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@43158.4]
  wire  _T_896; // @[SRAM.scala 148:25:@43159.4]
  wire  _T_897; // @[SRAM.scala 148:15:@43160.4]
  wire  _T_898; // @[SRAM.scala 149:15:@43162.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@43161.4]
  reg  regs_24; // @[SRAM.scala 145:20:@43168.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@43169.4]
  wire  _T_905; // @[SRAM.scala 148:25:@43170.4]
  wire  _T_906; // @[SRAM.scala 148:15:@43171.4]
  wire  _T_907; // @[SRAM.scala 149:15:@43173.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@43172.4]
  reg  regs_25; // @[SRAM.scala 145:20:@43179.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@43180.4]
  wire  _T_914; // @[SRAM.scala 148:25:@43181.4]
  wire  _T_915; // @[SRAM.scala 148:15:@43182.4]
  wire  _T_916; // @[SRAM.scala 149:15:@43184.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@43183.4]
  reg  regs_26; // @[SRAM.scala 145:20:@43190.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@43191.4]
  wire  _T_923; // @[SRAM.scala 148:25:@43192.4]
  wire  _T_924; // @[SRAM.scala 148:15:@43193.4]
  wire  _T_925; // @[SRAM.scala 149:15:@43195.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@43194.4]
  reg  regs_27; // @[SRAM.scala 145:20:@43201.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@43202.4]
  wire  _T_932; // @[SRAM.scala 148:25:@43203.4]
  wire  _T_933; // @[SRAM.scala 148:15:@43204.4]
  wire  _T_934; // @[SRAM.scala 149:15:@43206.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@43205.4]
  reg  regs_28; // @[SRAM.scala 145:20:@43212.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@43213.4]
  wire  _T_941; // @[SRAM.scala 148:25:@43214.4]
  wire  _T_942; // @[SRAM.scala 148:15:@43215.4]
  wire  _T_943; // @[SRAM.scala 149:15:@43217.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@43216.4]
  reg  regs_29; // @[SRAM.scala 145:20:@43223.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@43224.4]
  wire  _T_950; // @[SRAM.scala 148:25:@43225.4]
  wire  _T_951; // @[SRAM.scala 148:15:@43226.4]
  wire  _T_952; // @[SRAM.scala 149:15:@43228.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@43227.4]
  reg  regs_30; // @[SRAM.scala 145:20:@43234.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@43235.4]
  wire  _T_959; // @[SRAM.scala 148:25:@43236.4]
  wire  _T_960; // @[SRAM.scala 148:15:@43237.4]
  wire  _T_961; // @[SRAM.scala 149:15:@43239.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@43238.4]
  reg  regs_31; // @[SRAM.scala 145:20:@43245.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@43246.4]
  wire  _T_968; // @[SRAM.scala 148:25:@43247.4]
  wire  _T_969; // @[SRAM.scala 148:15:@43248.4]
  wire  _T_970; // @[SRAM.scala 149:15:@43250.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@43249.4]
  reg  regs_32; // @[SRAM.scala 145:20:@43256.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@43257.4]
  wire  _T_977; // @[SRAM.scala 148:25:@43258.4]
  wire  _T_978; // @[SRAM.scala 148:15:@43259.4]
  wire  _T_979; // @[SRAM.scala 149:15:@43261.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@43260.4]
  reg  regs_33; // @[SRAM.scala 145:20:@43267.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@43268.4]
  wire  _T_986; // @[SRAM.scala 148:25:@43269.4]
  wire  _T_987; // @[SRAM.scala 148:15:@43270.4]
  wire  _T_988; // @[SRAM.scala 149:15:@43272.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@43271.4]
  reg  regs_34; // @[SRAM.scala 145:20:@43278.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@43279.4]
  wire  _T_995; // @[SRAM.scala 148:25:@43280.4]
  wire  _T_996; // @[SRAM.scala 148:15:@43281.4]
  wire  _T_997; // @[SRAM.scala 149:15:@43283.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@43282.4]
  reg  regs_35; // @[SRAM.scala 145:20:@43289.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@43290.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@43291.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@43292.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@43294.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@43293.4]
  reg  regs_36; // @[SRAM.scala 145:20:@43300.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@43301.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@43302.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@43303.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@43305.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@43304.4]
  reg  regs_37; // @[SRAM.scala 145:20:@43311.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@43312.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@43313.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@43314.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@43316.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@43315.4]
  reg  regs_38; // @[SRAM.scala 145:20:@43322.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@43323.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@43324.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@43325.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@43327.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@43326.4]
  reg  regs_39; // @[SRAM.scala 145:20:@43333.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@43334.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@43335.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@43336.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@43338.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@43337.4]
  reg  regs_40; // @[SRAM.scala 145:20:@43344.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@43345.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@43346.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@43347.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@43349.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@43348.4]
  reg  regs_41; // @[SRAM.scala 145:20:@43355.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@43356.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@43357.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@43358.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@43360.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@43359.4]
  reg  regs_42; // @[SRAM.scala 145:20:@43366.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@43367.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@43368.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@43369.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@43371.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@43370.4]
  reg  regs_43; // @[SRAM.scala 145:20:@43377.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@43378.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@43379.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@43380.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@43382.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@43381.4]
  reg  regs_44; // @[SRAM.scala 145:20:@43388.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@43389.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@43390.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@43391.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@43393.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@43392.4]
  reg  regs_45; // @[SRAM.scala 145:20:@43399.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@43400.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@43401.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@43402.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@43404.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@43403.4]
  reg  regs_46; // @[SRAM.scala 145:20:@43410.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@43411.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@43412.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@43413.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@43415.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@43414.4]
  reg  regs_47; // @[SRAM.scala 145:20:@43421.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@43422.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@43423.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@43424.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@43426.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@43425.4]
  reg  regs_48; // @[SRAM.scala 145:20:@43432.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@43433.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@43434.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@43435.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@43437.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@43436.4]
  reg  regs_49; // @[SRAM.scala 145:20:@43443.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@43444.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@43445.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@43446.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@43448.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@43447.4]
  reg  regs_50; // @[SRAM.scala 145:20:@43454.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@43455.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@43456.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@43457.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@43459.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@43458.4]
  reg  regs_51; // @[SRAM.scala 145:20:@43465.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@43466.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@43467.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@43468.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@43470.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@43469.4]
  reg  regs_52; // @[SRAM.scala 145:20:@43476.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@43477.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@43478.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@43479.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@43481.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@43480.4]
  reg  regs_53; // @[SRAM.scala 145:20:@43487.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@43488.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@43489.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@43490.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@43492.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@43491.4]
  reg  regs_54; // @[SRAM.scala 145:20:@43498.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@43499.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@43500.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@43501.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@43503.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@43502.4]
  reg  regs_55; // @[SRAM.scala 145:20:@43509.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@43510.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@43511.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@43512.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@43514.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@43513.4]
  reg  regs_56; // @[SRAM.scala 145:20:@43520.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@43521.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@43522.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@43523.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@43525.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@43524.4]
  reg  regs_57; // @[SRAM.scala 145:20:@43531.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@43532.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@43533.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@43534.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@43536.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@43535.4]
  reg  regs_58; // @[SRAM.scala 145:20:@43542.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@43543.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@43544.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@43545.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@43547.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@43546.4]
  reg  regs_59; // @[SRAM.scala 145:20:@43553.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@43554.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@43555.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@43556.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@43558.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@43557.4]
  reg  regs_60; // @[SRAM.scala 145:20:@43564.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@43565.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@43566.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@43567.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@43569.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@43568.4]
  reg  regs_61; // @[SRAM.scala 145:20:@43575.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@43576.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@43577.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@43578.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@43580.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@43579.4]
  reg  regs_62; // @[SRAM.scala 145:20:@43586.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@43587.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@43588.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@43589.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@43591.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@43590.4]
  reg  regs_63; // @[SRAM.scala 145:20:@43597.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@43598.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@43599.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@43600.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@43602.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@43601.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@43671.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@43671.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@42905.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@42906.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@42907.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42909.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@42908.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@42916.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@42917.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@42918.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42920.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@42919.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@42927.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@42928.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@42929.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42931.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@42930.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@42938.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@42939.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@42940.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42942.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@42941.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@42949.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@42950.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@42951.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42953.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@42952.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@42960.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@42961.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@42962.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42964.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@42963.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@42971.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@42972.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@42973.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42975.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@42974.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@42982.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@42983.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@42984.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42986.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@42985.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@42993.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@42994.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@42995.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42997.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@42996.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@43004.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@43005.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@43006.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43008.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@43007.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@43015.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@43016.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@43017.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43019.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@43018.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@43026.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@43027.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@43028.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43030.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@43029.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@43037.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@43038.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@43039.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43041.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@43040.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@43048.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@43049.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@43050.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43052.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@43051.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@43059.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@43060.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@43061.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43063.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@43062.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@43070.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@43071.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@43072.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43074.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@43073.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@43081.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@43082.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@43083.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43085.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@43084.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@43092.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@43093.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@43094.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43096.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@43095.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@43103.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@43104.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@43105.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43107.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@43106.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@43114.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@43115.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@43116.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43118.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@43117.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@43125.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@43126.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@43127.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43129.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@43128.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@43136.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@43137.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@43138.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43140.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@43139.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@43147.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@43148.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@43149.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43151.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@43150.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@43158.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@43159.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@43160.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43162.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@43161.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@43169.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@43170.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@43171.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43173.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@43172.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@43180.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@43181.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@43182.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43184.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@43183.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@43191.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@43192.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@43193.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43195.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@43194.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@43202.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@43203.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@43204.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43206.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@43205.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@43213.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@43214.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@43215.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43217.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@43216.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@43224.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@43225.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@43226.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43228.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@43227.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@43235.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@43236.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@43237.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43239.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@43238.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@43246.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@43247.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@43248.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43250.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@43249.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@43257.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@43258.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@43259.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43261.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@43260.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@43268.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@43269.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@43270.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43272.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@43271.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@43279.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@43280.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@43281.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43283.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@43282.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@43290.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@43291.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@43292.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43294.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@43293.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@43301.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@43302.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@43303.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43305.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@43304.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@43312.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@43313.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@43314.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43316.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@43315.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@43323.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@43324.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@43325.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43327.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@43326.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@43334.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@43335.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@43336.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43338.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@43337.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@43345.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@43346.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@43347.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43349.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@43348.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@43356.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@43357.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@43358.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43360.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@43359.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@43367.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@43368.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@43369.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43371.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@43370.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@43378.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@43379.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@43380.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43382.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@43381.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@43389.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@43390.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@43391.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43393.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@43392.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@43400.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@43401.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@43402.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43404.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@43403.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@43411.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@43412.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@43413.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43415.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@43414.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@43422.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@43423.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@43424.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43426.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@43425.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@43433.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@43434.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@43435.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43437.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@43436.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@43444.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@43445.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@43446.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43448.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@43447.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@43455.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@43456.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@43457.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43459.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@43458.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@43466.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@43467.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@43468.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43470.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@43469.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@43477.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@43478.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@43479.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43481.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@43480.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@43488.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@43489.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@43490.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43492.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@43491.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@43499.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@43500.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@43501.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43503.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@43502.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@43510.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@43511.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@43512.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43514.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@43513.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@43521.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@43522.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@43523.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43525.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@43524.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@43532.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@43533.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@43534.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43536.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@43535.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@43543.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@43544.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@43545.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43547.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@43546.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@43554.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@43555.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@43556.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43558.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@43557.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@43565.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@43566.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@43567.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43569.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@43568.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@43576.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@43577.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@43578.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43580.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@43579.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@43587.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@43588.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@43589.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43591.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@43590.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@43598.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@43599.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@43600.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43602.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@43601.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@43671.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@43671.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@43671.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@43673.2]
  input   clock, // @[:@43674.4]
  input   reset, // @[:@43675.4]
  output  io_in_ready, // @[:@43676.4]
  input   io_in_valid, // @[:@43676.4]
  input   io_in_bits, // @[:@43676.4]
  input   io_out_ready, // @[:@43676.4]
  output  io_out_valid, // @[:@43676.4]
  output  io_out_bits, // @[:@43676.4]
  input   io_banks_0_wdata_valid, // @[:@43676.4]
  input   io_banks_0_wdata_bits, // @[:@43676.4]
  input   io_banks_1_wdata_valid, // @[:@43676.4]
  input   io_banks_1_wdata_bits, // @[:@43676.4]
  input   io_banks_2_wdata_valid, // @[:@43676.4]
  input   io_banks_2_wdata_bits, // @[:@43676.4]
  input   io_banks_3_wdata_valid, // @[:@43676.4]
  input   io_banks_3_wdata_bits, // @[:@43676.4]
  input   io_banks_4_wdata_valid, // @[:@43676.4]
  input   io_banks_4_wdata_bits, // @[:@43676.4]
  input   io_banks_5_wdata_valid, // @[:@43676.4]
  input   io_banks_5_wdata_bits, // @[:@43676.4]
  input   io_banks_6_wdata_valid, // @[:@43676.4]
  input   io_banks_6_wdata_bits, // @[:@43676.4]
  input   io_banks_7_wdata_valid, // @[:@43676.4]
  input   io_banks_7_wdata_bits, // @[:@43676.4]
  input   io_banks_8_wdata_valid, // @[:@43676.4]
  input   io_banks_8_wdata_bits, // @[:@43676.4]
  input   io_banks_9_wdata_valid, // @[:@43676.4]
  input   io_banks_9_wdata_bits, // @[:@43676.4]
  input   io_banks_10_wdata_valid, // @[:@43676.4]
  input   io_banks_10_wdata_bits, // @[:@43676.4]
  input   io_banks_11_wdata_valid, // @[:@43676.4]
  input   io_banks_11_wdata_bits, // @[:@43676.4]
  input   io_banks_12_wdata_valid, // @[:@43676.4]
  input   io_banks_12_wdata_bits, // @[:@43676.4]
  input   io_banks_13_wdata_valid, // @[:@43676.4]
  input   io_banks_13_wdata_bits, // @[:@43676.4]
  input   io_banks_14_wdata_valid, // @[:@43676.4]
  input   io_banks_14_wdata_bits, // @[:@43676.4]
  input   io_banks_15_wdata_valid, // @[:@43676.4]
  input   io_banks_15_wdata_bits, // @[:@43676.4]
  input   io_banks_16_wdata_valid, // @[:@43676.4]
  input   io_banks_16_wdata_bits, // @[:@43676.4]
  input   io_banks_17_wdata_valid, // @[:@43676.4]
  input   io_banks_17_wdata_bits, // @[:@43676.4]
  input   io_banks_18_wdata_valid, // @[:@43676.4]
  input   io_banks_18_wdata_bits, // @[:@43676.4]
  input   io_banks_19_wdata_valid, // @[:@43676.4]
  input   io_banks_19_wdata_bits, // @[:@43676.4]
  input   io_banks_20_wdata_valid, // @[:@43676.4]
  input   io_banks_20_wdata_bits, // @[:@43676.4]
  input   io_banks_21_wdata_valid, // @[:@43676.4]
  input   io_banks_21_wdata_bits, // @[:@43676.4]
  input   io_banks_22_wdata_valid, // @[:@43676.4]
  input   io_banks_22_wdata_bits, // @[:@43676.4]
  input   io_banks_23_wdata_valid, // @[:@43676.4]
  input   io_banks_23_wdata_bits, // @[:@43676.4]
  input   io_banks_24_wdata_valid, // @[:@43676.4]
  input   io_banks_24_wdata_bits, // @[:@43676.4]
  input   io_banks_25_wdata_valid, // @[:@43676.4]
  input   io_banks_25_wdata_bits, // @[:@43676.4]
  input   io_banks_26_wdata_valid, // @[:@43676.4]
  input   io_banks_26_wdata_bits, // @[:@43676.4]
  input   io_banks_27_wdata_valid, // @[:@43676.4]
  input   io_banks_27_wdata_bits, // @[:@43676.4]
  input   io_banks_28_wdata_valid, // @[:@43676.4]
  input   io_banks_28_wdata_bits, // @[:@43676.4]
  input   io_banks_29_wdata_valid, // @[:@43676.4]
  input   io_banks_29_wdata_bits, // @[:@43676.4]
  input   io_banks_30_wdata_valid, // @[:@43676.4]
  input   io_banks_30_wdata_bits, // @[:@43676.4]
  input   io_banks_31_wdata_valid, // @[:@43676.4]
  input   io_banks_31_wdata_bits, // @[:@43676.4]
  input   io_banks_32_wdata_valid, // @[:@43676.4]
  input   io_banks_32_wdata_bits, // @[:@43676.4]
  input   io_banks_33_wdata_valid, // @[:@43676.4]
  input   io_banks_33_wdata_bits, // @[:@43676.4]
  input   io_banks_34_wdata_valid, // @[:@43676.4]
  input   io_banks_34_wdata_bits, // @[:@43676.4]
  input   io_banks_35_wdata_valid, // @[:@43676.4]
  input   io_banks_35_wdata_bits, // @[:@43676.4]
  input   io_banks_36_wdata_valid, // @[:@43676.4]
  input   io_banks_36_wdata_bits, // @[:@43676.4]
  input   io_banks_37_wdata_valid, // @[:@43676.4]
  input   io_banks_37_wdata_bits, // @[:@43676.4]
  input   io_banks_38_wdata_valid, // @[:@43676.4]
  input   io_banks_38_wdata_bits, // @[:@43676.4]
  input   io_banks_39_wdata_valid, // @[:@43676.4]
  input   io_banks_39_wdata_bits, // @[:@43676.4]
  input   io_banks_40_wdata_valid, // @[:@43676.4]
  input   io_banks_40_wdata_bits, // @[:@43676.4]
  input   io_banks_41_wdata_valid, // @[:@43676.4]
  input   io_banks_41_wdata_bits, // @[:@43676.4]
  input   io_banks_42_wdata_valid, // @[:@43676.4]
  input   io_banks_42_wdata_bits, // @[:@43676.4]
  input   io_banks_43_wdata_valid, // @[:@43676.4]
  input   io_banks_43_wdata_bits, // @[:@43676.4]
  input   io_banks_44_wdata_valid, // @[:@43676.4]
  input   io_banks_44_wdata_bits, // @[:@43676.4]
  input   io_banks_45_wdata_valid, // @[:@43676.4]
  input   io_banks_45_wdata_bits, // @[:@43676.4]
  input   io_banks_46_wdata_valid, // @[:@43676.4]
  input   io_banks_46_wdata_bits, // @[:@43676.4]
  input   io_banks_47_wdata_valid, // @[:@43676.4]
  input   io_banks_47_wdata_bits, // @[:@43676.4]
  input   io_banks_48_wdata_valid, // @[:@43676.4]
  input   io_banks_48_wdata_bits, // @[:@43676.4]
  input   io_banks_49_wdata_valid, // @[:@43676.4]
  input   io_banks_49_wdata_bits, // @[:@43676.4]
  input   io_banks_50_wdata_valid, // @[:@43676.4]
  input   io_banks_50_wdata_bits, // @[:@43676.4]
  input   io_banks_51_wdata_valid, // @[:@43676.4]
  input   io_banks_51_wdata_bits, // @[:@43676.4]
  input   io_banks_52_wdata_valid, // @[:@43676.4]
  input   io_banks_52_wdata_bits, // @[:@43676.4]
  input   io_banks_53_wdata_valid, // @[:@43676.4]
  input   io_banks_53_wdata_bits, // @[:@43676.4]
  input   io_banks_54_wdata_valid, // @[:@43676.4]
  input   io_banks_54_wdata_bits, // @[:@43676.4]
  input   io_banks_55_wdata_valid, // @[:@43676.4]
  input   io_banks_55_wdata_bits, // @[:@43676.4]
  input   io_banks_56_wdata_valid, // @[:@43676.4]
  input   io_banks_56_wdata_bits, // @[:@43676.4]
  input   io_banks_57_wdata_valid, // @[:@43676.4]
  input   io_banks_57_wdata_bits, // @[:@43676.4]
  input   io_banks_58_wdata_valid, // @[:@43676.4]
  input   io_banks_58_wdata_bits, // @[:@43676.4]
  input   io_banks_59_wdata_valid, // @[:@43676.4]
  input   io_banks_59_wdata_bits, // @[:@43676.4]
  input   io_banks_60_wdata_valid, // @[:@43676.4]
  input   io_banks_60_wdata_bits, // @[:@43676.4]
  input   io_banks_61_wdata_valid, // @[:@43676.4]
  input   io_banks_61_wdata_bits, // @[:@43676.4]
  input   io_banks_62_wdata_valid, // @[:@43676.4]
  input   io_banks_62_wdata_bits, // @[:@43676.4]
  input   io_banks_63_wdata_valid, // @[:@43676.4]
  input   io_banks_63_wdata_bits // @[:@43676.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@43942.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@43942.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@43942.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@43942.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@43942.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@43952.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@43952.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@43952.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@43952.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@43952.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@43967.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@43967.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@43967.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@43967.4]
  wire  writeEn; // @[FIFO.scala 30:29:@43940.4]
  wire  readEn; // @[FIFO.scala 31:29:@43941.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@43962.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@43963.4]
  wire  _T_824; // @[FIFO.scala 45:27:@43964.4]
  wire  empty; // @[FIFO.scala 45:24:@43965.4]
  wire  full; // @[FIFO.scala 46:23:@43966.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@45133.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@45134.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@43942.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@43952.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@43967.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@43940.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@43941.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@43963.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@43964.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@43965.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@43966.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@45133.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@45134.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@45140.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@45138.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@44172.4]
  assign enqCounter_clock = clock; // @[:@43943.4]
  assign enqCounter_reset = reset; // @[:@43944.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@43950.4]
  assign deqCounter_clock = clock; // @[:@43953.4]
  assign deqCounter_reset = reset; // @[:@43954.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@43960.4]
  assign FFRAM_clock = clock; // @[:@43968.4]
  assign FFRAM_reset = reset; // @[:@43969.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@44168.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@44169.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@44170.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@44171.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@44174.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@44173.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@44177.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@44176.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@44180.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@44179.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@44183.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@44182.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@44186.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@44185.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@44189.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@44188.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@44192.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@44191.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@44195.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@44194.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@44198.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@44197.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@44201.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@44200.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@44204.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@44203.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@44207.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@44206.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@44210.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@44209.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@44213.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@44212.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@44216.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@44215.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@44219.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@44218.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@44222.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@44221.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@44225.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@44224.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@44228.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@44227.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@44231.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@44230.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@44234.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@44233.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@44237.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@44236.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@44240.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@44239.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@44243.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@44242.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@44246.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@44245.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@44249.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@44248.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@44252.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@44251.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@44255.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@44254.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@44258.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@44257.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@44261.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@44260.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@44264.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@44263.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@44267.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@44266.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@44270.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@44269.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@44273.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@44272.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@44276.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@44275.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@44279.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@44278.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@44282.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@44281.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@44285.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@44284.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@44288.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@44287.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@44291.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@44290.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@44294.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@44293.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@44297.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@44296.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@44300.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@44299.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@44303.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@44302.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@44306.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@44305.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@44309.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@44308.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@44312.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@44311.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@44315.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@44314.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@44318.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@44317.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@44321.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@44320.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@44324.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@44323.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@44327.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@44326.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@44330.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@44329.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@44333.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@44332.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@44336.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@44335.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@44339.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@44338.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@44342.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@44341.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@44345.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@44344.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@44348.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@44347.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@44351.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@44350.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@44354.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@44353.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@44357.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@44356.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@44360.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@44359.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@44363.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@44362.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@45142.2]
  input         clock, // @[:@45143.4]
  input         reset, // @[:@45144.4]
  input         io_dram_cmd_ready, // @[:@45145.4]
  output        io_dram_cmd_valid, // @[:@45145.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@45145.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@45145.4]
  input         io_dram_wdata_ready, // @[:@45145.4]
  output        io_dram_wdata_valid, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@45145.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@45145.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@45145.4]
  output        io_dram_wresp_ready, // @[:@45145.4]
  input         io_dram_wresp_valid, // @[:@45145.4]
  output        io_store_cmd_ready, // @[:@45145.4]
  input         io_store_cmd_valid, // @[:@45145.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@45145.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@45145.4]
  output        io_store_data_ready, // @[:@45145.4]
  input         io_store_data_valid, // @[:@45145.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@45145.4]
  input         io_store_data_bits_wstrb, // @[:@45145.4]
  input         io_store_wresp_ready, // @[:@45145.4]
  output        io_store_wresp_valid, // @[:@45145.4]
  output        io_store_wresp_bits // @[:@45145.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@45270.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@45270.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@45270.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@45270.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@45270.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@45270.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@45270.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@45270.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@45270.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@45270.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@45676.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@45676.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@45676.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@45676.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@45676.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@45676.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@45676.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@45676.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@45676.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@45917.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@45917.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@45673.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@45270.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@45676.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@45917.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@45673.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@45670.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@45671.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@45674.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@45706.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@45707.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@45708.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@45709.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@45710.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@45711.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@45712.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@45713.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@45714.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@45715.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@45716.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@45717.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@45718.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@45719.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@45720.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@45721.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@45722.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@45852.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@45853.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@45854.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@45855.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@45856.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@45857.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@45858.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@45859.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@45860.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@45861.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@45862.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@45863.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@45864.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@45865.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@45866.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@45867.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@45868.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@45869.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@45870.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@45871.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@45872.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@45873.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@45874.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@45875.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@45876.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@45877.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@45878.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@45879.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@45880.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@45881.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@45882.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@45883.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@45884.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@45885.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@45886.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@45887.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@45888.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@45889.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@45890.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@45891.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@45892.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@45893.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@45894.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@45895.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@45896.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@45897.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@45898.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@45899.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@45900.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@45901.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@45902.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@45903.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@45904.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@45905.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@45906.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@45907.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@45908.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@45909.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@45910.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@45911.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@45912.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@45913.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@45914.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@45915.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@46184.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@45668.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@45705.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@46185.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@46186.4]
  assign cmd_clock = clock; // @[:@45271.4]
  assign cmd_reset = reset; // @[:@45272.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@45665.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@45667.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@45666.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@45669.4]
  assign wdata_clock = clock; // @[:@45677.4]
  assign wdata_reset = reset; // @[:@45678.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@45702.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@45703.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@45704.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@45916.4]
  assign wresp_clock = clock; // @[:@45918.4]
  assign wresp_reset = reset; // @[:@45919.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@46182.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@46183.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@46187.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@46253.2]
  output        io_in_ready, // @[:@46256.4]
  input         io_in_valid, // @[:@46256.4]
  input  [63:0] io_in_bits_0_addr, // @[:@46256.4]
  input  [31:0] io_in_bits_0_size, // @[:@46256.4]
  input         io_in_bits_0_isWr, // @[:@46256.4]
  input  [31:0] io_in_bits_0_tag, // @[:@46256.4]
  input         io_out_ready, // @[:@46256.4]
  output        io_out_valid, // @[:@46256.4]
  output [63:0] io_out_bits_addr, // @[:@46256.4]
  output [31:0] io_out_bits_size, // @[:@46256.4]
  output        io_out_bits_isWr, // @[:@46256.4]
  output [31:0] io_out_bits_tag // @[:@46256.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@46258.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@46258.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@46267.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@46266.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@46272.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@46271.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@46269.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@46268.4]
endmodule
module MuxPipe_1( // @[:@46274.2]
  output        io_in_ready, // @[:@46277.4]
  input         io_in_valid, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@46277.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@46277.4]
  input         io_in_bits_0_wstrb_0, // @[:@46277.4]
  input         io_in_bits_0_wstrb_1, // @[:@46277.4]
  input         io_in_bits_0_wstrb_2, // @[:@46277.4]
  input         io_in_bits_0_wstrb_3, // @[:@46277.4]
  input         io_in_bits_0_wstrb_4, // @[:@46277.4]
  input         io_in_bits_0_wstrb_5, // @[:@46277.4]
  input         io_in_bits_0_wstrb_6, // @[:@46277.4]
  input         io_in_bits_0_wstrb_7, // @[:@46277.4]
  input         io_in_bits_0_wstrb_8, // @[:@46277.4]
  input         io_in_bits_0_wstrb_9, // @[:@46277.4]
  input         io_in_bits_0_wstrb_10, // @[:@46277.4]
  input         io_in_bits_0_wstrb_11, // @[:@46277.4]
  input         io_in_bits_0_wstrb_12, // @[:@46277.4]
  input         io_in_bits_0_wstrb_13, // @[:@46277.4]
  input         io_in_bits_0_wstrb_14, // @[:@46277.4]
  input         io_in_bits_0_wstrb_15, // @[:@46277.4]
  input         io_in_bits_0_wstrb_16, // @[:@46277.4]
  input         io_in_bits_0_wstrb_17, // @[:@46277.4]
  input         io_in_bits_0_wstrb_18, // @[:@46277.4]
  input         io_in_bits_0_wstrb_19, // @[:@46277.4]
  input         io_in_bits_0_wstrb_20, // @[:@46277.4]
  input         io_in_bits_0_wstrb_21, // @[:@46277.4]
  input         io_in_bits_0_wstrb_22, // @[:@46277.4]
  input         io_in_bits_0_wstrb_23, // @[:@46277.4]
  input         io_in_bits_0_wstrb_24, // @[:@46277.4]
  input         io_in_bits_0_wstrb_25, // @[:@46277.4]
  input         io_in_bits_0_wstrb_26, // @[:@46277.4]
  input         io_in_bits_0_wstrb_27, // @[:@46277.4]
  input         io_in_bits_0_wstrb_28, // @[:@46277.4]
  input         io_in_bits_0_wstrb_29, // @[:@46277.4]
  input         io_in_bits_0_wstrb_30, // @[:@46277.4]
  input         io_in_bits_0_wstrb_31, // @[:@46277.4]
  input         io_in_bits_0_wstrb_32, // @[:@46277.4]
  input         io_in_bits_0_wstrb_33, // @[:@46277.4]
  input         io_in_bits_0_wstrb_34, // @[:@46277.4]
  input         io_in_bits_0_wstrb_35, // @[:@46277.4]
  input         io_in_bits_0_wstrb_36, // @[:@46277.4]
  input         io_in_bits_0_wstrb_37, // @[:@46277.4]
  input         io_in_bits_0_wstrb_38, // @[:@46277.4]
  input         io_in_bits_0_wstrb_39, // @[:@46277.4]
  input         io_in_bits_0_wstrb_40, // @[:@46277.4]
  input         io_in_bits_0_wstrb_41, // @[:@46277.4]
  input         io_in_bits_0_wstrb_42, // @[:@46277.4]
  input         io_in_bits_0_wstrb_43, // @[:@46277.4]
  input         io_in_bits_0_wstrb_44, // @[:@46277.4]
  input         io_in_bits_0_wstrb_45, // @[:@46277.4]
  input         io_in_bits_0_wstrb_46, // @[:@46277.4]
  input         io_in_bits_0_wstrb_47, // @[:@46277.4]
  input         io_in_bits_0_wstrb_48, // @[:@46277.4]
  input         io_in_bits_0_wstrb_49, // @[:@46277.4]
  input         io_in_bits_0_wstrb_50, // @[:@46277.4]
  input         io_in_bits_0_wstrb_51, // @[:@46277.4]
  input         io_in_bits_0_wstrb_52, // @[:@46277.4]
  input         io_in_bits_0_wstrb_53, // @[:@46277.4]
  input         io_in_bits_0_wstrb_54, // @[:@46277.4]
  input         io_in_bits_0_wstrb_55, // @[:@46277.4]
  input         io_in_bits_0_wstrb_56, // @[:@46277.4]
  input         io_in_bits_0_wstrb_57, // @[:@46277.4]
  input         io_in_bits_0_wstrb_58, // @[:@46277.4]
  input         io_in_bits_0_wstrb_59, // @[:@46277.4]
  input         io_in_bits_0_wstrb_60, // @[:@46277.4]
  input         io_in_bits_0_wstrb_61, // @[:@46277.4]
  input         io_in_bits_0_wstrb_62, // @[:@46277.4]
  input         io_in_bits_0_wstrb_63, // @[:@46277.4]
  input         io_out_ready, // @[:@46277.4]
  output        io_out_valid, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_0, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_1, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_2, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_3, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_4, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_5, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_6, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_7, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_8, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_9, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_10, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_11, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_12, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_13, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_14, // @[:@46277.4]
  output [31:0] io_out_bits_wdata_15, // @[:@46277.4]
  output        io_out_bits_wstrb_0, // @[:@46277.4]
  output        io_out_bits_wstrb_1, // @[:@46277.4]
  output        io_out_bits_wstrb_2, // @[:@46277.4]
  output        io_out_bits_wstrb_3, // @[:@46277.4]
  output        io_out_bits_wstrb_4, // @[:@46277.4]
  output        io_out_bits_wstrb_5, // @[:@46277.4]
  output        io_out_bits_wstrb_6, // @[:@46277.4]
  output        io_out_bits_wstrb_7, // @[:@46277.4]
  output        io_out_bits_wstrb_8, // @[:@46277.4]
  output        io_out_bits_wstrb_9, // @[:@46277.4]
  output        io_out_bits_wstrb_10, // @[:@46277.4]
  output        io_out_bits_wstrb_11, // @[:@46277.4]
  output        io_out_bits_wstrb_12, // @[:@46277.4]
  output        io_out_bits_wstrb_13, // @[:@46277.4]
  output        io_out_bits_wstrb_14, // @[:@46277.4]
  output        io_out_bits_wstrb_15, // @[:@46277.4]
  output        io_out_bits_wstrb_16, // @[:@46277.4]
  output        io_out_bits_wstrb_17, // @[:@46277.4]
  output        io_out_bits_wstrb_18, // @[:@46277.4]
  output        io_out_bits_wstrb_19, // @[:@46277.4]
  output        io_out_bits_wstrb_20, // @[:@46277.4]
  output        io_out_bits_wstrb_21, // @[:@46277.4]
  output        io_out_bits_wstrb_22, // @[:@46277.4]
  output        io_out_bits_wstrb_23, // @[:@46277.4]
  output        io_out_bits_wstrb_24, // @[:@46277.4]
  output        io_out_bits_wstrb_25, // @[:@46277.4]
  output        io_out_bits_wstrb_26, // @[:@46277.4]
  output        io_out_bits_wstrb_27, // @[:@46277.4]
  output        io_out_bits_wstrb_28, // @[:@46277.4]
  output        io_out_bits_wstrb_29, // @[:@46277.4]
  output        io_out_bits_wstrb_30, // @[:@46277.4]
  output        io_out_bits_wstrb_31, // @[:@46277.4]
  output        io_out_bits_wstrb_32, // @[:@46277.4]
  output        io_out_bits_wstrb_33, // @[:@46277.4]
  output        io_out_bits_wstrb_34, // @[:@46277.4]
  output        io_out_bits_wstrb_35, // @[:@46277.4]
  output        io_out_bits_wstrb_36, // @[:@46277.4]
  output        io_out_bits_wstrb_37, // @[:@46277.4]
  output        io_out_bits_wstrb_38, // @[:@46277.4]
  output        io_out_bits_wstrb_39, // @[:@46277.4]
  output        io_out_bits_wstrb_40, // @[:@46277.4]
  output        io_out_bits_wstrb_41, // @[:@46277.4]
  output        io_out_bits_wstrb_42, // @[:@46277.4]
  output        io_out_bits_wstrb_43, // @[:@46277.4]
  output        io_out_bits_wstrb_44, // @[:@46277.4]
  output        io_out_bits_wstrb_45, // @[:@46277.4]
  output        io_out_bits_wstrb_46, // @[:@46277.4]
  output        io_out_bits_wstrb_47, // @[:@46277.4]
  output        io_out_bits_wstrb_48, // @[:@46277.4]
  output        io_out_bits_wstrb_49, // @[:@46277.4]
  output        io_out_bits_wstrb_50, // @[:@46277.4]
  output        io_out_bits_wstrb_51, // @[:@46277.4]
  output        io_out_bits_wstrb_52, // @[:@46277.4]
  output        io_out_bits_wstrb_53, // @[:@46277.4]
  output        io_out_bits_wstrb_54, // @[:@46277.4]
  output        io_out_bits_wstrb_55, // @[:@46277.4]
  output        io_out_bits_wstrb_56, // @[:@46277.4]
  output        io_out_bits_wstrb_57, // @[:@46277.4]
  output        io_out_bits_wstrb_58, // @[:@46277.4]
  output        io_out_bits_wstrb_59, // @[:@46277.4]
  output        io_out_bits_wstrb_60, // @[:@46277.4]
  output        io_out_bits_wstrb_61, // @[:@46277.4]
  output        io_out_bits_wstrb_62, // @[:@46277.4]
  output        io_out_bits_wstrb_63 // @[:@46277.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@46279.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@46279.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@46364.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@46363.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@46430.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@46431.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@46432.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@46433.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@46434.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@46435.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@46436.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@46437.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@46438.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@46439.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@46440.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@46441.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@46442.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@46443.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@46444.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@46445.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@46366.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@46367.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@46368.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@46369.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@46370.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@46371.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@46372.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@46373.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@46374.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@46375.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@46376.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@46377.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@46378.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@46379.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@46380.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@46381.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@46382.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@46383.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@46384.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@46385.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@46386.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@46387.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@46388.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@46389.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@46390.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@46391.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@46392.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@46393.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@46394.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@46395.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@46396.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@46397.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@46398.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@46399.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@46400.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@46401.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@46402.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@46403.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@46404.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@46405.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@46406.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@46407.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@46408.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@46409.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@46410.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@46411.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@46412.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@46413.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@46414.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@46415.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@46416.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@46417.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@46418.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@46419.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@46420.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@46421.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@46422.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@46423.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@46424.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@46425.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@46426.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@46427.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@46428.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@46429.4]
endmodule
module ElementCounter( // @[:@46447.2]
  input         clock, // @[:@46448.4]
  input         reset, // @[:@46449.4]
  input         io_reset, // @[:@46450.4]
  input         io_enable, // @[:@46450.4]
  output [31:0] io_out // @[:@46450.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@46452.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@46453.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@46454.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@46459.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@46455.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@46453.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@46454.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@46459.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@46455.4]
  assign io_out = count; // @[Counter.scala 47:10:@46462.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@46464.2]
  input         clock, // @[:@46465.4]
  input         reset, // @[:@46466.4]
  output        io_app_0_cmd_ready, // @[:@46467.4]
  input         io_app_0_cmd_valid, // @[:@46467.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@46467.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@46467.4]
  input         io_app_0_cmd_bits_isWr, // @[:@46467.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@46467.4]
  output        io_app_0_wdata_ready, // @[:@46467.4]
  input         io_app_0_wdata_valid, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@46467.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@46467.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@46467.4]
  input         io_app_0_rresp_ready, // @[:@46467.4]
  input         io_app_0_wresp_ready, // @[:@46467.4]
  output        io_app_0_wresp_valid, // @[:@46467.4]
  input         io_dram_cmd_ready, // @[:@46467.4]
  output        io_dram_cmd_valid, // @[:@46467.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@46467.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@46467.4]
  output        io_dram_cmd_bits_isWr, // @[:@46467.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@46467.4]
  input         io_dram_wdata_ready, // @[:@46467.4]
  output        io_dram_wdata_valid, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@46467.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@46467.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@46467.4]
  output        io_dram_rresp_ready, // @[:@46467.4]
  output        io_dram_wresp_ready, // @[:@46467.4]
  input         io_dram_wresp_valid, // @[:@46467.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@46467.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@46696.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@46696.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@46696.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@46696.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@46696.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@46703.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@46703.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@46703.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@46703.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@46703.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@46713.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@46713.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@46713.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@46713.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@46713.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@46713.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@46713.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@46713.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@46713.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@46713.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@46713.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@46713.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@46736.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@46736.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@46739.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@46739.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@46739.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@46739.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@46739.4]
  wire  _T_346; // @[package.scala 96:25:@46708.4 package.scala 96:25:@46709.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@46710.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@46712.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@46728.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@46730.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@46733.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@46742.4]
  wire [31:0] _T_365; // @[:@46746.4 :@46747.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@46748.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@46754.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@46757.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@46758.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@46945.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@46952.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@46957.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@46961.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@46962.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@46986.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@46696.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@46703.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@46713.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@46736.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@46739.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@46708.4 package.scala 96:25:@46709.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@46710.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@46712.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@46728.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@46730.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@46733.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@46742.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@46746.4 :@46747.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@46748.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@46754.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@46757.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@46758.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@46945.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@46952.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@46957.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@46961.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@46962.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@46986.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@46959.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@46965.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@46988.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@46848.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@46847.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@46846.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@46844.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@46843.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@46931.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@46915.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@46916.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@46917.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@46918.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@46919.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@46920.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@46921.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@46922.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@46923.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@46924.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@46925.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@46926.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@46927.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@46928.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@46929.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@46930.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@46851.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@46852.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@46853.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@46854.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@46855.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@46856.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@46857.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@46858.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@46859.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@46860.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@46861.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@46862.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@46863.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@46864.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@46865.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@46866.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@46867.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@46868.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@46869.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@46870.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@46871.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@46872.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@46873.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@46874.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@46875.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@46876.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@46877.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@46878.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@46879.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@46880.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@46881.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@46882.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@46883.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@46884.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@46885.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@46886.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@46887.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@46888.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@46889.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@46890.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@46891.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@46892.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@46893.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@46894.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@46895.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@46896.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@46897.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@46898.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@46899.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@46900.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@46901.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@46902.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@46903.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@46904.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@46905.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@46906.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@46907.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@46908.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@46909.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@46910.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@46911.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@46912.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@46913.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@46914.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@46992.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@46995.4]
  assign RetimeWrapper_clock = clock; // @[:@46697.4]
  assign RetimeWrapper_reset = reset; // @[:@46698.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@46700.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@46699.4]
  assign RetimeWrapper_1_clock = clock; // @[:@46704.4]
  assign RetimeWrapper_1_reset = reset; // @[:@46705.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@46707.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@46706.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@46716.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@46722.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@46721.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@46719.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@46718.4 FringeBundles.scala 115:32:@46735.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@46849.4 StreamArbiter.scala 57:23:@46955.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@46760.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@46827.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@46828.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@46829.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@46830.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@46831.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@46832.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@46833.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@46834.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@46835.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@46836.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@46837.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@46838.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@46839.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@46840.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@46841.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@46842.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@46763.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@46764.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@46765.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@46766.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@46767.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@46768.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@46769.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@46770.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@46771.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@46772.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@46773.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@46774.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@46775.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@46776.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@46777.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@46778.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@46779.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@46780.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@46781.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@46782.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@46783.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@46784.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@46785.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@46786.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@46787.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@46788.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@46789.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@46790.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@46791.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@46792.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@46793.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@46794.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@46795.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@46796.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@46797.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@46798.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@46799.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@46800.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@46801.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@46802.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@46803.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@46804.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@46805.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@46806.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@46807.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@46808.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@46809.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@46810.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@46811.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@46812.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@46813.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@46814.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@46815.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@46816.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@46817.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@46818.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@46819.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@46820.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@46821.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@46822.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@46823.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@46824.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@46825.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@46826.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@46932.4 StreamArbiter.scala 58:25:@46956.4]
  assign elementCtr_clock = clock; // @[:@46740.4]
  assign elementCtr_reset = reset; // @[:@46741.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@46744.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@46743.4]
endmodule
module Counter_72( // @[:@46997.2]
  input         clock, // @[:@46998.4]
  input         reset, // @[:@46999.4]
  input         io_reset, // @[:@47000.4]
  input         io_enable, // @[:@47000.4]
  input  [31:0] io_stride, // @[:@47000.4]
  output [31:0] io_out, // @[:@47000.4]
  output [31:0] io_next // @[:@47000.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@47002.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@47003.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@47004.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@47009.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@47005.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@47003.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@47004.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@47009.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@47005.4]
  assign io_out = count; // @[Counter.scala 25:10:@47012.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@47013.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@47015.2]
  input         clock, // @[:@47016.4]
  input         reset, // @[:@47017.4]
  output        io_in_cmd_ready, // @[:@47018.4]
  input         io_in_cmd_valid, // @[:@47018.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@47018.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@47018.4]
  input         io_in_cmd_bits_isWr, // @[:@47018.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@47018.4]
  output        io_in_wdata_ready, // @[:@47018.4]
  input         io_in_wdata_valid, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@47018.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@47018.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@47018.4]
  input         io_in_rresp_ready, // @[:@47018.4]
  input         io_in_wresp_ready, // @[:@47018.4]
  output        io_in_wresp_valid, // @[:@47018.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@47018.4]
  input         io_out_cmd_ready, // @[:@47018.4]
  output        io_out_cmd_valid, // @[:@47018.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@47018.4]
  output [31:0] io_out_cmd_bits_size, // @[:@47018.4]
  output        io_out_cmd_bits_isWr, // @[:@47018.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@47018.4]
  input         io_out_wdata_ready, // @[:@47018.4]
  output        io_out_wdata_valid, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@47018.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@47018.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@47018.4]
  output        io_out_rresp_ready, // @[:@47018.4]
  output        io_out_wresp_ready, // @[:@47018.4]
  input         io_out_wresp_valid, // @[:@47018.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@47018.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@47132.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@47132.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@47132.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@47132.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@47132.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@47132.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@47132.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@47135.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@47136.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@47137.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@47138.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@47141.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@47141.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@47142.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@47142.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@47143.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@47146.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@47153.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@47157.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@47160.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@47163.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@47174.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@47132.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@47135.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@47136.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@47137.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@47138.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@47141.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@47141.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@47142.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@47142.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@47143.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@47146.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@47153.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@47157.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@47160.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@47163.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@47174.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@47131.4 AXIProtocol.scala 38:19:@47165.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@47124.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@47021.4 AXIProtocol.scala 46:21:@47179.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@47020.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@47130.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@47129.4 AXIProtocol.scala 29:24:@47148.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@47128.4 AXIProtocol.scala 25:24:@47140.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@47126.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@47125.4 FringeBundles.scala 115:32:@47162.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@47123.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@47107.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@47108.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@47109.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@47110.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@47111.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@47112.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@47113.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@47114.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@47115.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@47116.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@47117.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@47118.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@47119.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@47120.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@47121.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@47122.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@47043.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@47044.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@47045.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@47046.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@47047.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@47048.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@47049.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@47050.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@47051.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@47052.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@47053.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@47054.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@47055.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@47056.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@47057.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@47058.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@47059.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@47060.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@47061.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@47062.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@47063.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@47064.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@47065.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@47066.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@47067.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@47068.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@47069.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@47070.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@47071.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@47072.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@47073.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@47074.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@47075.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@47076.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@47077.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@47078.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@47079.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@47080.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@47081.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@47082.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@47083.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@47084.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@47085.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@47086.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@47087.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@47088.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@47089.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@47090.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@47091.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@47092.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@47093.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@47094.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@47095.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@47096.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@47097.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@47098.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@47099.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@47100.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@47101.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@47102.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@47103.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@47104.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@47105.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@47106.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@47041.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@47022.4 AXIProtocol.scala 47:22:@47181.4]
  assign cmdSizeCounter_clock = clock; // @[:@47133.4]
  assign cmdSizeCounter_reset = reset; // @[:@47134.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@47166.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@47167.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@47168.4]
endmodule
module AXICmdIssue( // @[:@47201.2]
  input         clock, // @[:@47202.4]
  input         reset, // @[:@47203.4]
  output        io_in_cmd_ready, // @[:@47204.4]
  input         io_in_cmd_valid, // @[:@47204.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@47204.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@47204.4]
  input         io_in_cmd_bits_isWr, // @[:@47204.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@47204.4]
  output        io_in_wdata_ready, // @[:@47204.4]
  input         io_in_wdata_valid, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@47204.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@47204.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@47204.4]
  input         io_in_rresp_ready, // @[:@47204.4]
  input         io_in_wresp_ready, // @[:@47204.4]
  output        io_in_wresp_valid, // @[:@47204.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@47204.4]
  input         io_out_cmd_ready, // @[:@47204.4]
  output        io_out_cmd_valid, // @[:@47204.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@47204.4]
  output [31:0] io_out_cmd_bits_size, // @[:@47204.4]
  output        io_out_cmd_bits_isWr, // @[:@47204.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@47204.4]
  input         io_out_wdata_ready, // @[:@47204.4]
  output        io_out_wdata_valid, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@47204.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@47204.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@47204.4]
  output        io_out_wdata_bits_wlast, // @[:@47204.4]
  output        io_out_rresp_ready, // @[:@47204.4]
  output        io_out_wresp_ready, // @[:@47204.4]
  input         io_out_wresp_valid, // @[:@47204.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@47204.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@47318.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@47318.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@47318.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@47318.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@47318.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@47318.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@47318.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@47321.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@47322.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@47323.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@47324.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@47325.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@47331.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@47332.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@47327.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@47341.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@47342.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@47318.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@47322.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@47323.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@47324.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@47325.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@47331.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@47332.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@47327.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@47341.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@47342.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@47317.4 AXIProtocol.scala 81:19:@47339.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@47310.4 AXIProtocol.scala 82:21:@47340.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@47207.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@47206.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@47316.4 AXIProtocol.scala 84:20:@47344.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@47315.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@47314.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@47312.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@47311.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@47309.4 AXIProtocol.scala 86:22:@47346.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@47293.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@47294.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@47295.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@47296.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@47297.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@47298.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@47299.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@47300.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@47301.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@47302.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@47303.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@47304.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@47305.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@47306.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@47307.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@47308.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@47229.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@47230.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@47231.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@47232.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@47233.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@47234.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@47235.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@47236.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@47237.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@47238.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@47239.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@47240.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@47241.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@47242.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@47243.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@47244.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@47245.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@47246.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@47247.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@47248.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@47249.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@47250.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@47251.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@47252.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@47253.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@47254.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@47255.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@47256.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@47257.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@47258.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@47259.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@47260.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@47261.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@47262.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@47263.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@47264.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@47265.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@47266.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@47267.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@47268.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@47269.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@47270.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@47271.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@47272.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@47273.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@47274.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@47275.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@47276.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@47277.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@47278.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@47279.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@47280.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@47281.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@47282.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@47283.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@47284.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@47285.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@47286.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@47287.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@47288.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@47289.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@47290.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@47291.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@47292.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@47228.4 AXIProtocol.scala 87:27:@47347.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@47227.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@47208.4]
  assign wdataCounter_clock = clock; // @[:@47319.4]
  assign wdataCounter_reset = reset; // @[:@47320.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@47335.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@47336.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@47337.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@47349.2]
  input         clock, // @[:@47350.4]
  input         reset, // @[:@47351.4]
  input         io_enable, // @[:@47352.4]
  output        io_app_stores_0_cmd_ready, // @[:@47352.4]
  input         io_app_stores_0_cmd_valid, // @[:@47352.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@47352.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@47352.4]
  output        io_app_stores_0_data_ready, // @[:@47352.4]
  input         io_app_stores_0_data_valid, // @[:@47352.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@47352.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@47352.4]
  input         io_app_stores_0_wresp_ready, // @[:@47352.4]
  output        io_app_stores_0_wresp_valid, // @[:@47352.4]
  output        io_app_stores_0_wresp_bits, // @[:@47352.4]
  input         io_dram_cmd_ready, // @[:@47352.4]
  output        io_dram_cmd_valid, // @[:@47352.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@47352.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@47352.4]
  output        io_dram_cmd_bits_isWr, // @[:@47352.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@47352.4]
  input         io_dram_wdata_ready, // @[:@47352.4]
  output        io_dram_wdata_valid, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@47352.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@47352.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@47352.4]
  output        io_dram_wdata_bits_wlast, // @[:@47352.4]
  output        io_dram_rresp_ready, // @[:@47352.4]
  output        io_dram_wresp_ready, // @[:@47352.4]
  input         io_dram_wresp_valid, // @[:@47352.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@47352.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@48238.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@48252.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@48480.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@48595.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@48595.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@48238.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@48252.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@48480.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@48595.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@48251.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@48247.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@48242.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@48241.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@48820.4 DRAMArbiter.scala 100:23:@48823.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@48819.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@48818.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@48816.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@48815.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@48813.4 DRAMArbiter.scala 101:25:@48825.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@48797.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@48798.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@48799.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@48800.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@48801.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@48802.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@48803.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@48804.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@48805.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@48806.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@48807.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@48808.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@48809.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@48810.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@48811.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@48812.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@48733.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@48734.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@48735.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@48736.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@48737.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@48738.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@48739.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@48740.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@48741.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@48742.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@48743.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@48744.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@48745.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@48746.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@48747.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@48748.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@48749.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@48750.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@48751.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@48752.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@48753.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@48754.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@48755.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@48756.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@48757.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@48758.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@48759.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@48760.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@48761.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@48762.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@48763.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@48764.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@48765.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@48766.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@48767.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@48768.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@48769.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@48770.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@48771.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@48772.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@48773.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@48774.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@48775.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@48776.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@48777.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@48778.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@48779.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@48780.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@48781.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@48782.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@48783.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@48784.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@48785.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@48786.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@48787.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@48788.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@48789.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@48790.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@48791.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@48792.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@48793.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@48794.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@48795.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@48796.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@48732.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@48731.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@48712.4]
  assign StreamControllerStore_clock = clock; // @[:@48239.4]
  assign StreamControllerStore_reset = reset; // @[:@48240.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@48367.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@48360.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@48257.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@48250.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@48249.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@48248.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@48246.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@48245.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@48244.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@48243.4]
  assign StreamArbiter_clock = clock; // @[:@48253.4]
  assign StreamArbiter_reset = reset; // @[:@48254.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@48478.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@48477.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@48476.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@48474.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@48473.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@48471.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@48455.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@48456.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@48457.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@48458.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@48459.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@48460.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@48461.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@48462.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@48463.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@48464.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@48465.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@48466.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@48467.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@48468.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@48469.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@48470.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@48391.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@48392.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@48393.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@48394.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@48395.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@48396.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@48397.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@48398.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@48399.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@48400.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@48401.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@48402.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@48403.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@48404.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@48405.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@48406.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@48407.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@48408.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@48409.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@48410.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@48411.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@48412.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@48413.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@48414.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@48415.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@48416.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@48417.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@48418.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@48419.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@48420.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@48421.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@48422.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@48423.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@48424.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@48425.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@48426.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@48427.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@48428.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@48429.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@48430.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@48431.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@48432.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@48433.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@48434.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@48435.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@48436.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@48437.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@48438.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@48439.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@48440.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@48441.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@48442.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@48443.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@48444.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@48445.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@48446.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@48447.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@48448.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@48449.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@48450.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@48451.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@48452.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@48453.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@48454.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@48389.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@48370.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@48594.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@48587.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@48484.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@48483.4]
  assign AXICmdSplit_clock = clock; // @[:@48481.4]
  assign AXICmdSplit_reset = reset; // @[:@48482.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@48593.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@48592.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@48591.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@48589.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@48588.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@48586.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@48570.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@48571.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@48572.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@48573.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@48574.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@48575.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@48576.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@48577.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@48578.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@48579.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@48580.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@48581.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@48582.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@48583.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@48584.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@48585.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@48506.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@48507.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@48508.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@48509.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@48510.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@48511.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@48512.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@48513.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@48514.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@48515.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@48516.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@48517.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@48518.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@48519.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@48520.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@48521.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@48522.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@48523.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@48524.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@48525.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@48526.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@48527.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@48528.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@48529.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@48530.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@48531.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@48532.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@48533.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@48534.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@48535.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@48536.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@48537.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@48538.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@48539.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@48540.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@48541.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@48542.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@48543.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@48544.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@48545.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@48546.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@48547.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@48548.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@48549.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@48550.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@48551.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@48552.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@48553.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@48554.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@48555.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@48556.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@48557.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@48558.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@48559.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@48560.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@48561.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@48562.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@48563.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@48564.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@48565.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@48566.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@48567.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@48568.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@48569.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@48504.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@48485.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@48709.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@48702.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@48599.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@48598.4]
  assign AXICmdIssue_clock = clock; // @[:@48596.4]
  assign AXICmdIssue_reset = reset; // @[:@48597.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@48708.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@48707.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@48706.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@48704.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@48703.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@48701.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@48685.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@48686.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@48687.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@48688.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@48689.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@48690.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@48691.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@48692.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@48693.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@48694.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@48695.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@48696.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@48697.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@48698.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@48699.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@48700.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@48621.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@48622.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@48623.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@48624.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@48625.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@48626.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@48627.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@48628.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@48629.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@48630.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@48631.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@48632.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@48633.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@48634.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@48635.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@48636.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@48637.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@48638.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@48639.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@48640.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@48641.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@48642.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@48643.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@48644.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@48645.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@48646.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@48647.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@48648.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@48649.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@48650.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@48651.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@48652.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@48653.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@48654.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@48655.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@48656.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@48657.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@48658.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@48659.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@48660.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@48661.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@48662.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@48663.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@48664.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@48665.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@48666.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@48667.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@48668.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@48669.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@48670.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@48671.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@48672.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@48673.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@48674.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@48675.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@48676.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@48677.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@48678.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@48679.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@48680.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@48681.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@48682.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@48683.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@48684.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@48619.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@48600.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@48821.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@48814.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@48711.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@48710.4]
endmodule
module DRAMArbiter_1( // @[:@63050.2]
  input         clock, // @[:@63051.4]
  input         reset, // @[:@63052.4]
  input         io_enable, // @[:@63053.4]
  input         io_dram_cmd_ready, // @[:@63053.4]
  output        io_dram_cmd_valid, // @[:@63053.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@63053.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@63053.4]
  output        io_dram_cmd_bits_isWr, // @[:@63053.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@63053.4]
  input         io_dram_wdata_ready, // @[:@63053.4]
  output        io_dram_wdata_valid, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@63053.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@63053.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@63053.4]
  output        io_dram_wdata_bits_wlast, // @[:@63053.4]
  output        io_dram_rresp_ready, // @[:@63053.4]
  output        io_dram_wresp_ready, // @[:@63053.4]
  input         io_dram_wresp_valid, // @[:@63053.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@63053.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@63939.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@63953.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@64181.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@64296.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@64296.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@63939.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@63953.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@64181.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@64296.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@64521.4 DRAMArbiter.scala 100:23:@64524.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@64520.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@64519.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@64517.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@64516.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@64514.4 DRAMArbiter.scala 101:25:@64526.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@64498.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@64499.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@64500.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@64501.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@64502.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@64503.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@64504.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@64505.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@64506.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@64507.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@64508.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@64509.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@64510.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@64511.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@64512.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@64513.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@64434.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@64435.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@64436.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@64437.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@64438.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@64439.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@64440.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@64441.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@64442.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@64443.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@64444.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@64445.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@64446.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@64447.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@64448.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@64449.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@64450.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@64451.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@64452.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@64453.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@64454.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@64455.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@64456.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@64457.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@64458.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@64459.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@64460.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@64461.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@64462.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@64463.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@64464.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@64465.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@64466.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@64467.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@64468.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@64469.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@64470.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@64471.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@64472.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@64473.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@64474.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@64475.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@64476.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@64477.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@64478.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@64479.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@64480.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@64481.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@64482.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@64483.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@64484.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@64485.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@64486.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@64487.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@64488.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@64489.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@64490.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@64491.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@64492.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@64493.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@64494.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@64495.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@64496.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@64497.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@64433.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@64432.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@64413.4]
  assign StreamControllerStore_clock = clock; // @[:@63940.4]
  assign StreamControllerStore_reset = reset; // @[:@63941.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@64068.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@64061.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@63958.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@63951.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@63950.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@63949.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@63947.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@63946.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@63945.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@63944.4]
  assign StreamArbiter_clock = clock; // @[:@63954.4]
  assign StreamArbiter_reset = reset; // @[:@63955.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@64179.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@64178.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@64177.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@64175.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@64174.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@64172.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@64156.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@64157.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@64158.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@64159.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@64160.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@64161.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@64162.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@64163.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@64164.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@64165.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@64166.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@64167.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@64168.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@64169.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@64170.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@64171.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@64092.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@64093.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@64094.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@64095.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@64096.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@64097.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@64098.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@64099.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@64100.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@64101.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@64102.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@64103.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@64104.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@64105.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@64106.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@64107.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@64108.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@64109.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@64110.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@64111.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@64112.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@64113.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@64114.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@64115.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@64116.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@64117.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@64118.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@64119.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@64120.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@64121.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@64122.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@64123.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@64124.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@64125.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@64126.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@64127.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@64128.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@64129.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@64130.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@64131.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@64132.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@64133.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@64134.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@64135.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@64136.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@64137.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@64138.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@64139.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@64140.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@64141.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@64142.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@64143.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@64144.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@64145.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@64146.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@64147.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@64148.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@64149.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@64150.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@64151.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@64152.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@64153.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@64154.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@64155.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@64090.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@64071.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@64295.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@64288.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@64185.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@64184.4]
  assign AXICmdSplit_clock = clock; // @[:@64182.4]
  assign AXICmdSplit_reset = reset; // @[:@64183.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@64294.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@64293.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@64292.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@64290.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@64289.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@64287.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@64271.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@64272.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@64273.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@64274.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@64275.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@64276.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@64277.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@64278.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@64279.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@64280.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@64281.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@64282.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@64283.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@64284.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@64285.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@64286.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@64207.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@64208.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@64209.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@64210.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@64211.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@64212.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@64213.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@64214.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@64215.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@64216.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@64217.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@64218.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@64219.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@64220.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@64221.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@64222.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@64223.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@64224.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@64225.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@64226.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@64227.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@64228.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@64229.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@64230.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@64231.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@64232.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@64233.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@64234.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@64235.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@64236.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@64237.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@64238.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@64239.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@64240.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@64241.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@64242.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@64243.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@64244.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@64245.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@64246.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@64247.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@64248.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@64249.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@64250.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@64251.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@64252.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@64253.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@64254.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@64255.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@64256.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@64257.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@64258.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@64259.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@64260.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@64261.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@64262.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@64263.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@64264.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@64265.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@64266.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@64267.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@64268.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@64269.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@64270.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@64205.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@64186.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@64410.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@64403.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@64300.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@64299.4]
  assign AXICmdIssue_clock = clock; // @[:@64297.4]
  assign AXICmdIssue_reset = reset; // @[:@64298.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@64409.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@64408.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@64407.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@64405.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@64404.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@64402.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@64386.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@64387.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@64388.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@64389.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@64390.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@64391.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@64392.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@64393.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@64394.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@64395.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@64396.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@64397.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@64398.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@64399.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@64400.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@64401.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@64322.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@64323.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@64324.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@64325.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@64326.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@64327.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@64328.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@64329.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@64330.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@64331.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@64332.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@64333.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@64334.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@64335.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@64336.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@64337.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@64338.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@64339.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@64340.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@64341.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@64342.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@64343.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@64344.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@64345.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@64346.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@64347.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@64348.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@64349.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@64350.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@64351.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@64352.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@64353.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@64354.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@64355.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@64356.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@64357.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@64358.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@64359.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@64360.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@64361.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@64362.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@64363.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@64364.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@64365.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@64366.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@64367.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@64368.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@64369.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@64370.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@64371.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@64372.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@64373.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@64374.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@64375.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@64376.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@64377.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@64378.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@64379.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@64380.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@64381.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@64382.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@64383.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@64384.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@64385.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@64320.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@64301.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@64522.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@64515.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@64412.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@64411.4]
endmodule
module DRAMHeap( // @[:@95158.2]
  input         io_accel_0_req_valid, // @[:@95161.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@95161.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@95161.4]
  output        io_accel_0_resp_valid, // @[:@95161.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@95161.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@95161.4]
  output        io_host_0_req_valid, // @[:@95161.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@95161.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@95161.4]
  input         io_host_0_resp_valid, // @[:@95161.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@95161.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@95161.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@95168.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@95170.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@95169.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@95165.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@95164.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@95163.4]
endmodule
module FringeFF( // @[:@95204.2]
  input         clock, // @[:@95205.4]
  input         reset, // @[:@95206.4]
  input  [63:0] io_in, // @[:@95207.4]
  input         io_reset, // @[:@95207.4]
  output [63:0] io_out, // @[:@95207.4]
  input         io_enable // @[:@95207.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@95210.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@95210.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@95210.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@95210.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@95210.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@95215.4 package.scala 96:25:@95216.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@95221.6]
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@95210.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@95215.4 package.scala 96:25:@95216.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@95221.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@95227.4]
  assign RetimeWrapper_clock = clock; // @[:@95211.4]
  assign RetimeWrapper_reset = reset; // @[:@95212.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@95214.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@95213.4]
endmodule
module MuxN( // @[:@123843.2]
  input  [63:0] io_ins_0, // @[:@123846.4]
  input  [63:0] io_ins_1, // @[:@123846.4]
  input  [63:0] io_ins_2, // @[:@123846.4]
  input  [63:0] io_ins_3, // @[:@123846.4]
  input  [63:0] io_ins_4, // @[:@123846.4]
  input  [63:0] io_ins_5, // @[:@123846.4]
  input  [63:0] io_ins_6, // @[:@123846.4]
  input  [63:0] io_ins_7, // @[:@123846.4]
  input  [63:0] io_ins_8, // @[:@123846.4]
  input  [63:0] io_ins_9, // @[:@123846.4]
  input  [63:0] io_ins_10, // @[:@123846.4]
  input  [63:0] io_ins_11, // @[:@123846.4]
  input  [63:0] io_ins_12, // @[:@123846.4]
  input  [63:0] io_ins_13, // @[:@123846.4]
  input  [63:0] io_ins_14, // @[:@123846.4]
  input  [63:0] io_ins_15, // @[:@123846.4]
  input  [63:0] io_ins_16, // @[:@123846.4]
  input  [63:0] io_ins_17, // @[:@123846.4]
  input  [63:0] io_ins_18, // @[:@123846.4]
  input  [63:0] io_ins_19, // @[:@123846.4]
  input  [63:0] io_ins_20, // @[:@123846.4]
  input  [63:0] io_ins_21, // @[:@123846.4]
  input  [63:0] io_ins_22, // @[:@123846.4]
  input  [63:0] io_ins_23, // @[:@123846.4]
  input  [63:0] io_ins_24, // @[:@123846.4]
  input  [63:0] io_ins_25, // @[:@123846.4]
  input  [63:0] io_ins_26, // @[:@123846.4]
  input  [63:0] io_ins_27, // @[:@123846.4]
  input  [63:0] io_ins_28, // @[:@123846.4]
  input  [63:0] io_ins_29, // @[:@123846.4]
  input  [63:0] io_ins_30, // @[:@123846.4]
  input  [63:0] io_ins_31, // @[:@123846.4]
  input  [63:0] io_ins_32, // @[:@123846.4]
  input  [63:0] io_ins_33, // @[:@123846.4]
  input  [63:0] io_ins_34, // @[:@123846.4]
  input  [63:0] io_ins_35, // @[:@123846.4]
  input  [63:0] io_ins_36, // @[:@123846.4]
  input  [63:0] io_ins_37, // @[:@123846.4]
  input  [63:0] io_ins_38, // @[:@123846.4]
  input  [63:0] io_ins_39, // @[:@123846.4]
  input  [63:0] io_ins_40, // @[:@123846.4]
  input  [63:0] io_ins_41, // @[:@123846.4]
  input  [63:0] io_ins_42, // @[:@123846.4]
  input  [63:0] io_ins_43, // @[:@123846.4]
  input  [63:0] io_ins_44, // @[:@123846.4]
  input  [63:0] io_ins_45, // @[:@123846.4]
  input  [63:0] io_ins_46, // @[:@123846.4]
  input  [63:0] io_ins_47, // @[:@123846.4]
  input  [63:0] io_ins_48, // @[:@123846.4]
  input  [63:0] io_ins_49, // @[:@123846.4]
  input  [63:0] io_ins_50, // @[:@123846.4]
  input  [63:0] io_ins_51, // @[:@123846.4]
  input  [63:0] io_ins_52, // @[:@123846.4]
  input  [63:0] io_ins_53, // @[:@123846.4]
  input  [63:0] io_ins_54, // @[:@123846.4]
  input  [63:0] io_ins_55, // @[:@123846.4]
  input  [63:0] io_ins_56, // @[:@123846.4]
  input  [63:0] io_ins_57, // @[:@123846.4]
  input  [63:0] io_ins_58, // @[:@123846.4]
  input  [63:0] io_ins_59, // @[:@123846.4]
  input  [63:0] io_ins_60, // @[:@123846.4]
  input  [63:0] io_ins_61, // @[:@123846.4]
  input  [63:0] io_ins_62, // @[:@123846.4]
  input  [63:0] io_ins_63, // @[:@123846.4]
  input  [63:0] io_ins_64, // @[:@123846.4]
  input  [63:0] io_ins_65, // @[:@123846.4]
  input  [63:0] io_ins_66, // @[:@123846.4]
  input  [63:0] io_ins_67, // @[:@123846.4]
  input  [63:0] io_ins_68, // @[:@123846.4]
  input  [63:0] io_ins_69, // @[:@123846.4]
  input  [63:0] io_ins_70, // @[:@123846.4]
  input  [63:0] io_ins_71, // @[:@123846.4]
  input  [63:0] io_ins_72, // @[:@123846.4]
  input  [63:0] io_ins_73, // @[:@123846.4]
  input  [63:0] io_ins_74, // @[:@123846.4]
  input  [63:0] io_ins_75, // @[:@123846.4]
  input  [63:0] io_ins_76, // @[:@123846.4]
  input  [63:0] io_ins_77, // @[:@123846.4]
  input  [63:0] io_ins_78, // @[:@123846.4]
  input  [63:0] io_ins_79, // @[:@123846.4]
  input  [63:0] io_ins_80, // @[:@123846.4]
  input  [63:0] io_ins_81, // @[:@123846.4]
  input  [63:0] io_ins_82, // @[:@123846.4]
  input  [63:0] io_ins_83, // @[:@123846.4]
  input  [63:0] io_ins_84, // @[:@123846.4]
  input  [63:0] io_ins_85, // @[:@123846.4]
  input  [63:0] io_ins_86, // @[:@123846.4]
  input  [63:0] io_ins_87, // @[:@123846.4]
  input  [63:0] io_ins_88, // @[:@123846.4]
  input  [63:0] io_ins_89, // @[:@123846.4]
  input  [63:0] io_ins_90, // @[:@123846.4]
  input  [63:0] io_ins_91, // @[:@123846.4]
  input  [63:0] io_ins_92, // @[:@123846.4]
  input  [63:0] io_ins_93, // @[:@123846.4]
  input  [63:0] io_ins_94, // @[:@123846.4]
  input  [63:0] io_ins_95, // @[:@123846.4]
  input  [63:0] io_ins_96, // @[:@123846.4]
  input  [63:0] io_ins_97, // @[:@123846.4]
  input  [63:0] io_ins_98, // @[:@123846.4]
  input  [63:0] io_ins_99, // @[:@123846.4]
  input  [63:0] io_ins_100, // @[:@123846.4]
  input  [63:0] io_ins_101, // @[:@123846.4]
  input  [63:0] io_ins_102, // @[:@123846.4]
  input  [63:0] io_ins_103, // @[:@123846.4]
  input  [63:0] io_ins_104, // @[:@123846.4]
  input  [63:0] io_ins_105, // @[:@123846.4]
  input  [63:0] io_ins_106, // @[:@123846.4]
  input  [63:0] io_ins_107, // @[:@123846.4]
  input  [63:0] io_ins_108, // @[:@123846.4]
  input  [63:0] io_ins_109, // @[:@123846.4]
  input  [63:0] io_ins_110, // @[:@123846.4]
  input  [63:0] io_ins_111, // @[:@123846.4]
  input  [63:0] io_ins_112, // @[:@123846.4]
  input  [63:0] io_ins_113, // @[:@123846.4]
  input  [63:0] io_ins_114, // @[:@123846.4]
  input  [63:0] io_ins_115, // @[:@123846.4]
  input  [63:0] io_ins_116, // @[:@123846.4]
  input  [63:0] io_ins_117, // @[:@123846.4]
  input  [63:0] io_ins_118, // @[:@123846.4]
  input  [63:0] io_ins_119, // @[:@123846.4]
  input  [63:0] io_ins_120, // @[:@123846.4]
  input  [63:0] io_ins_121, // @[:@123846.4]
  input  [63:0] io_ins_122, // @[:@123846.4]
  input  [63:0] io_ins_123, // @[:@123846.4]
  input  [63:0] io_ins_124, // @[:@123846.4]
  input  [63:0] io_ins_125, // @[:@123846.4]
  input  [63:0] io_ins_126, // @[:@123846.4]
  input  [63:0] io_ins_127, // @[:@123846.4]
  input  [63:0] io_ins_128, // @[:@123846.4]
  input  [63:0] io_ins_129, // @[:@123846.4]
  input  [63:0] io_ins_130, // @[:@123846.4]
  input  [63:0] io_ins_131, // @[:@123846.4]
  input  [63:0] io_ins_132, // @[:@123846.4]
  input  [63:0] io_ins_133, // @[:@123846.4]
  input  [63:0] io_ins_134, // @[:@123846.4]
  input  [63:0] io_ins_135, // @[:@123846.4]
  input  [63:0] io_ins_136, // @[:@123846.4]
  input  [63:0] io_ins_137, // @[:@123846.4]
  input  [63:0] io_ins_138, // @[:@123846.4]
  input  [63:0] io_ins_139, // @[:@123846.4]
  input  [63:0] io_ins_140, // @[:@123846.4]
  input  [63:0] io_ins_141, // @[:@123846.4]
  input  [63:0] io_ins_142, // @[:@123846.4]
  input  [63:0] io_ins_143, // @[:@123846.4]
  input  [63:0] io_ins_144, // @[:@123846.4]
  input  [63:0] io_ins_145, // @[:@123846.4]
  input  [63:0] io_ins_146, // @[:@123846.4]
  input  [63:0] io_ins_147, // @[:@123846.4]
  input  [63:0] io_ins_148, // @[:@123846.4]
  input  [63:0] io_ins_149, // @[:@123846.4]
  input  [63:0] io_ins_150, // @[:@123846.4]
  input  [63:0] io_ins_151, // @[:@123846.4]
  input  [63:0] io_ins_152, // @[:@123846.4]
  input  [63:0] io_ins_153, // @[:@123846.4]
  input  [63:0] io_ins_154, // @[:@123846.4]
  input  [63:0] io_ins_155, // @[:@123846.4]
  input  [63:0] io_ins_156, // @[:@123846.4]
  input  [63:0] io_ins_157, // @[:@123846.4]
  input  [63:0] io_ins_158, // @[:@123846.4]
  input  [63:0] io_ins_159, // @[:@123846.4]
  input  [63:0] io_ins_160, // @[:@123846.4]
  input  [63:0] io_ins_161, // @[:@123846.4]
  input  [63:0] io_ins_162, // @[:@123846.4]
  input  [63:0] io_ins_163, // @[:@123846.4]
  input  [63:0] io_ins_164, // @[:@123846.4]
  input  [63:0] io_ins_165, // @[:@123846.4]
  input  [63:0] io_ins_166, // @[:@123846.4]
  input  [63:0] io_ins_167, // @[:@123846.4]
  input  [63:0] io_ins_168, // @[:@123846.4]
  input  [63:0] io_ins_169, // @[:@123846.4]
  input  [63:0] io_ins_170, // @[:@123846.4]
  input  [63:0] io_ins_171, // @[:@123846.4]
  input  [63:0] io_ins_172, // @[:@123846.4]
  input  [63:0] io_ins_173, // @[:@123846.4]
  input  [63:0] io_ins_174, // @[:@123846.4]
  input  [63:0] io_ins_175, // @[:@123846.4]
  input  [63:0] io_ins_176, // @[:@123846.4]
  input  [63:0] io_ins_177, // @[:@123846.4]
  input  [63:0] io_ins_178, // @[:@123846.4]
  input  [63:0] io_ins_179, // @[:@123846.4]
  input  [63:0] io_ins_180, // @[:@123846.4]
  input  [63:0] io_ins_181, // @[:@123846.4]
  input  [63:0] io_ins_182, // @[:@123846.4]
  input  [63:0] io_ins_183, // @[:@123846.4]
  input  [63:0] io_ins_184, // @[:@123846.4]
  input  [63:0] io_ins_185, // @[:@123846.4]
  input  [63:0] io_ins_186, // @[:@123846.4]
  input  [63:0] io_ins_187, // @[:@123846.4]
  input  [63:0] io_ins_188, // @[:@123846.4]
  input  [63:0] io_ins_189, // @[:@123846.4]
  input  [63:0] io_ins_190, // @[:@123846.4]
  input  [63:0] io_ins_191, // @[:@123846.4]
  input  [63:0] io_ins_192, // @[:@123846.4]
  input  [63:0] io_ins_193, // @[:@123846.4]
  input  [63:0] io_ins_194, // @[:@123846.4]
  input  [63:0] io_ins_195, // @[:@123846.4]
  input  [63:0] io_ins_196, // @[:@123846.4]
  input  [63:0] io_ins_197, // @[:@123846.4]
  input  [63:0] io_ins_198, // @[:@123846.4]
  input  [63:0] io_ins_199, // @[:@123846.4]
  input  [63:0] io_ins_200, // @[:@123846.4]
  input  [63:0] io_ins_201, // @[:@123846.4]
  input  [63:0] io_ins_202, // @[:@123846.4]
  input  [63:0] io_ins_203, // @[:@123846.4]
  input  [63:0] io_ins_204, // @[:@123846.4]
  input  [63:0] io_ins_205, // @[:@123846.4]
  input  [63:0] io_ins_206, // @[:@123846.4]
  input  [63:0] io_ins_207, // @[:@123846.4]
  input  [63:0] io_ins_208, // @[:@123846.4]
  input  [63:0] io_ins_209, // @[:@123846.4]
  input  [63:0] io_ins_210, // @[:@123846.4]
  input  [63:0] io_ins_211, // @[:@123846.4]
  input  [63:0] io_ins_212, // @[:@123846.4]
  input  [63:0] io_ins_213, // @[:@123846.4]
  input  [63:0] io_ins_214, // @[:@123846.4]
  input  [63:0] io_ins_215, // @[:@123846.4]
  input  [63:0] io_ins_216, // @[:@123846.4]
  input  [63:0] io_ins_217, // @[:@123846.4]
  input  [63:0] io_ins_218, // @[:@123846.4]
  input  [63:0] io_ins_219, // @[:@123846.4]
  input  [63:0] io_ins_220, // @[:@123846.4]
  input  [63:0] io_ins_221, // @[:@123846.4]
  input  [63:0] io_ins_222, // @[:@123846.4]
  input  [63:0] io_ins_223, // @[:@123846.4]
  input  [63:0] io_ins_224, // @[:@123846.4]
  input  [63:0] io_ins_225, // @[:@123846.4]
  input  [63:0] io_ins_226, // @[:@123846.4]
  input  [63:0] io_ins_227, // @[:@123846.4]
  input  [63:0] io_ins_228, // @[:@123846.4]
  input  [63:0] io_ins_229, // @[:@123846.4]
  input  [63:0] io_ins_230, // @[:@123846.4]
  input  [63:0] io_ins_231, // @[:@123846.4]
  input  [63:0] io_ins_232, // @[:@123846.4]
  input  [63:0] io_ins_233, // @[:@123846.4]
  input  [63:0] io_ins_234, // @[:@123846.4]
  input  [63:0] io_ins_235, // @[:@123846.4]
  input  [63:0] io_ins_236, // @[:@123846.4]
  input  [63:0] io_ins_237, // @[:@123846.4]
  input  [63:0] io_ins_238, // @[:@123846.4]
  input  [63:0] io_ins_239, // @[:@123846.4]
  input  [63:0] io_ins_240, // @[:@123846.4]
  input  [63:0] io_ins_241, // @[:@123846.4]
  input  [63:0] io_ins_242, // @[:@123846.4]
  input  [63:0] io_ins_243, // @[:@123846.4]
  input  [63:0] io_ins_244, // @[:@123846.4]
  input  [63:0] io_ins_245, // @[:@123846.4]
  input  [63:0] io_ins_246, // @[:@123846.4]
  input  [63:0] io_ins_247, // @[:@123846.4]
  input  [63:0] io_ins_248, // @[:@123846.4]
  input  [63:0] io_ins_249, // @[:@123846.4]
  input  [63:0] io_ins_250, // @[:@123846.4]
  input  [63:0] io_ins_251, // @[:@123846.4]
  input  [63:0] io_ins_252, // @[:@123846.4]
  input  [63:0] io_ins_253, // @[:@123846.4]
  input  [63:0] io_ins_254, // @[:@123846.4]
  input  [63:0] io_ins_255, // @[:@123846.4]
  input  [63:0] io_ins_256, // @[:@123846.4]
  input  [63:0] io_ins_257, // @[:@123846.4]
  input  [63:0] io_ins_258, // @[:@123846.4]
  input  [63:0] io_ins_259, // @[:@123846.4]
  input  [63:0] io_ins_260, // @[:@123846.4]
  input  [63:0] io_ins_261, // @[:@123846.4]
  input  [63:0] io_ins_262, // @[:@123846.4]
  input  [63:0] io_ins_263, // @[:@123846.4]
  input  [63:0] io_ins_264, // @[:@123846.4]
  input  [63:0] io_ins_265, // @[:@123846.4]
  input  [63:0] io_ins_266, // @[:@123846.4]
  input  [63:0] io_ins_267, // @[:@123846.4]
  input  [63:0] io_ins_268, // @[:@123846.4]
  input  [63:0] io_ins_269, // @[:@123846.4]
  input  [63:0] io_ins_270, // @[:@123846.4]
  input  [63:0] io_ins_271, // @[:@123846.4]
  input  [63:0] io_ins_272, // @[:@123846.4]
  input  [63:0] io_ins_273, // @[:@123846.4]
  input  [63:0] io_ins_274, // @[:@123846.4]
  input  [63:0] io_ins_275, // @[:@123846.4]
  input  [63:0] io_ins_276, // @[:@123846.4]
  input  [63:0] io_ins_277, // @[:@123846.4]
  input  [63:0] io_ins_278, // @[:@123846.4]
  input  [63:0] io_ins_279, // @[:@123846.4]
  input  [63:0] io_ins_280, // @[:@123846.4]
  input  [63:0] io_ins_281, // @[:@123846.4]
  input  [63:0] io_ins_282, // @[:@123846.4]
  input  [63:0] io_ins_283, // @[:@123846.4]
  input  [63:0] io_ins_284, // @[:@123846.4]
  input  [63:0] io_ins_285, // @[:@123846.4]
  input  [63:0] io_ins_286, // @[:@123846.4]
  input  [63:0] io_ins_287, // @[:@123846.4]
  input  [63:0] io_ins_288, // @[:@123846.4]
  input  [63:0] io_ins_289, // @[:@123846.4]
  input  [63:0] io_ins_290, // @[:@123846.4]
  input  [63:0] io_ins_291, // @[:@123846.4]
  input  [63:0] io_ins_292, // @[:@123846.4]
  input  [63:0] io_ins_293, // @[:@123846.4]
  input  [63:0] io_ins_294, // @[:@123846.4]
  input  [63:0] io_ins_295, // @[:@123846.4]
  input  [63:0] io_ins_296, // @[:@123846.4]
  input  [63:0] io_ins_297, // @[:@123846.4]
  input  [63:0] io_ins_298, // @[:@123846.4]
  input  [63:0] io_ins_299, // @[:@123846.4]
  input  [63:0] io_ins_300, // @[:@123846.4]
  input  [63:0] io_ins_301, // @[:@123846.4]
  input  [63:0] io_ins_302, // @[:@123846.4]
  input  [63:0] io_ins_303, // @[:@123846.4]
  input  [63:0] io_ins_304, // @[:@123846.4]
  input  [63:0] io_ins_305, // @[:@123846.4]
  input  [63:0] io_ins_306, // @[:@123846.4]
  input  [63:0] io_ins_307, // @[:@123846.4]
  input  [63:0] io_ins_308, // @[:@123846.4]
  input  [63:0] io_ins_309, // @[:@123846.4]
  input  [63:0] io_ins_310, // @[:@123846.4]
  input  [63:0] io_ins_311, // @[:@123846.4]
  input  [63:0] io_ins_312, // @[:@123846.4]
  input  [63:0] io_ins_313, // @[:@123846.4]
  input  [63:0] io_ins_314, // @[:@123846.4]
  input  [63:0] io_ins_315, // @[:@123846.4]
  input  [63:0] io_ins_316, // @[:@123846.4]
  input  [63:0] io_ins_317, // @[:@123846.4]
  input  [63:0] io_ins_318, // @[:@123846.4]
  input  [63:0] io_ins_319, // @[:@123846.4]
  input  [63:0] io_ins_320, // @[:@123846.4]
  input  [63:0] io_ins_321, // @[:@123846.4]
  input  [63:0] io_ins_322, // @[:@123846.4]
  input  [63:0] io_ins_323, // @[:@123846.4]
  input  [63:0] io_ins_324, // @[:@123846.4]
  input  [63:0] io_ins_325, // @[:@123846.4]
  input  [63:0] io_ins_326, // @[:@123846.4]
  input  [63:0] io_ins_327, // @[:@123846.4]
  input  [63:0] io_ins_328, // @[:@123846.4]
  input  [63:0] io_ins_329, // @[:@123846.4]
  input  [63:0] io_ins_330, // @[:@123846.4]
  input  [63:0] io_ins_331, // @[:@123846.4]
  input  [63:0] io_ins_332, // @[:@123846.4]
  input  [63:0] io_ins_333, // @[:@123846.4]
  input  [63:0] io_ins_334, // @[:@123846.4]
  input  [63:0] io_ins_335, // @[:@123846.4]
  input  [63:0] io_ins_336, // @[:@123846.4]
  input  [63:0] io_ins_337, // @[:@123846.4]
  input  [63:0] io_ins_338, // @[:@123846.4]
  input  [63:0] io_ins_339, // @[:@123846.4]
  input  [63:0] io_ins_340, // @[:@123846.4]
  input  [63:0] io_ins_341, // @[:@123846.4]
  input  [63:0] io_ins_342, // @[:@123846.4]
  input  [63:0] io_ins_343, // @[:@123846.4]
  input  [63:0] io_ins_344, // @[:@123846.4]
  input  [63:0] io_ins_345, // @[:@123846.4]
  input  [63:0] io_ins_346, // @[:@123846.4]
  input  [63:0] io_ins_347, // @[:@123846.4]
  input  [63:0] io_ins_348, // @[:@123846.4]
  input  [63:0] io_ins_349, // @[:@123846.4]
  input  [63:0] io_ins_350, // @[:@123846.4]
  input  [63:0] io_ins_351, // @[:@123846.4]
  input  [63:0] io_ins_352, // @[:@123846.4]
  input  [63:0] io_ins_353, // @[:@123846.4]
  input  [63:0] io_ins_354, // @[:@123846.4]
  input  [63:0] io_ins_355, // @[:@123846.4]
  input  [63:0] io_ins_356, // @[:@123846.4]
  input  [63:0] io_ins_357, // @[:@123846.4]
  input  [63:0] io_ins_358, // @[:@123846.4]
  input  [63:0] io_ins_359, // @[:@123846.4]
  input  [63:0] io_ins_360, // @[:@123846.4]
  input  [63:0] io_ins_361, // @[:@123846.4]
  input  [63:0] io_ins_362, // @[:@123846.4]
  input  [63:0] io_ins_363, // @[:@123846.4]
  input  [63:0] io_ins_364, // @[:@123846.4]
  input  [63:0] io_ins_365, // @[:@123846.4]
  input  [63:0] io_ins_366, // @[:@123846.4]
  input  [63:0] io_ins_367, // @[:@123846.4]
  input  [63:0] io_ins_368, // @[:@123846.4]
  input  [63:0] io_ins_369, // @[:@123846.4]
  input  [63:0] io_ins_370, // @[:@123846.4]
  input  [63:0] io_ins_371, // @[:@123846.4]
  input  [63:0] io_ins_372, // @[:@123846.4]
  input  [63:0] io_ins_373, // @[:@123846.4]
  input  [63:0] io_ins_374, // @[:@123846.4]
  input  [63:0] io_ins_375, // @[:@123846.4]
  input  [63:0] io_ins_376, // @[:@123846.4]
  input  [63:0] io_ins_377, // @[:@123846.4]
  input  [63:0] io_ins_378, // @[:@123846.4]
  input  [63:0] io_ins_379, // @[:@123846.4]
  input  [63:0] io_ins_380, // @[:@123846.4]
  input  [63:0] io_ins_381, // @[:@123846.4]
  input  [63:0] io_ins_382, // @[:@123846.4]
  input  [63:0] io_ins_383, // @[:@123846.4]
  input  [63:0] io_ins_384, // @[:@123846.4]
  input  [63:0] io_ins_385, // @[:@123846.4]
  input  [63:0] io_ins_386, // @[:@123846.4]
  input  [63:0] io_ins_387, // @[:@123846.4]
  input  [63:0] io_ins_388, // @[:@123846.4]
  input  [63:0] io_ins_389, // @[:@123846.4]
  input  [63:0] io_ins_390, // @[:@123846.4]
  input  [63:0] io_ins_391, // @[:@123846.4]
  input  [63:0] io_ins_392, // @[:@123846.4]
  input  [63:0] io_ins_393, // @[:@123846.4]
  input  [63:0] io_ins_394, // @[:@123846.4]
  input  [63:0] io_ins_395, // @[:@123846.4]
  input  [63:0] io_ins_396, // @[:@123846.4]
  input  [63:0] io_ins_397, // @[:@123846.4]
  input  [63:0] io_ins_398, // @[:@123846.4]
  input  [63:0] io_ins_399, // @[:@123846.4]
  input  [63:0] io_ins_400, // @[:@123846.4]
  input  [63:0] io_ins_401, // @[:@123846.4]
  input  [63:0] io_ins_402, // @[:@123846.4]
  input  [63:0] io_ins_403, // @[:@123846.4]
  input  [63:0] io_ins_404, // @[:@123846.4]
  input  [63:0] io_ins_405, // @[:@123846.4]
  input  [63:0] io_ins_406, // @[:@123846.4]
  input  [63:0] io_ins_407, // @[:@123846.4]
  input  [63:0] io_ins_408, // @[:@123846.4]
  input  [63:0] io_ins_409, // @[:@123846.4]
  input  [63:0] io_ins_410, // @[:@123846.4]
  input  [63:0] io_ins_411, // @[:@123846.4]
  input  [63:0] io_ins_412, // @[:@123846.4]
  input  [63:0] io_ins_413, // @[:@123846.4]
  input  [63:0] io_ins_414, // @[:@123846.4]
  input  [63:0] io_ins_415, // @[:@123846.4]
  input  [63:0] io_ins_416, // @[:@123846.4]
  input  [63:0] io_ins_417, // @[:@123846.4]
  input  [63:0] io_ins_418, // @[:@123846.4]
  input  [63:0] io_ins_419, // @[:@123846.4]
  input  [63:0] io_ins_420, // @[:@123846.4]
  input  [63:0] io_ins_421, // @[:@123846.4]
  input  [63:0] io_ins_422, // @[:@123846.4]
  input  [63:0] io_ins_423, // @[:@123846.4]
  input  [63:0] io_ins_424, // @[:@123846.4]
  input  [63:0] io_ins_425, // @[:@123846.4]
  input  [63:0] io_ins_426, // @[:@123846.4]
  input  [63:0] io_ins_427, // @[:@123846.4]
  input  [63:0] io_ins_428, // @[:@123846.4]
  input  [63:0] io_ins_429, // @[:@123846.4]
  input  [63:0] io_ins_430, // @[:@123846.4]
  input  [63:0] io_ins_431, // @[:@123846.4]
  input  [63:0] io_ins_432, // @[:@123846.4]
  input  [63:0] io_ins_433, // @[:@123846.4]
  input  [63:0] io_ins_434, // @[:@123846.4]
  input  [63:0] io_ins_435, // @[:@123846.4]
  input  [63:0] io_ins_436, // @[:@123846.4]
  input  [63:0] io_ins_437, // @[:@123846.4]
  input  [63:0] io_ins_438, // @[:@123846.4]
  input  [63:0] io_ins_439, // @[:@123846.4]
  input  [63:0] io_ins_440, // @[:@123846.4]
  input  [63:0] io_ins_441, // @[:@123846.4]
  input  [63:0] io_ins_442, // @[:@123846.4]
  input  [63:0] io_ins_443, // @[:@123846.4]
  input  [63:0] io_ins_444, // @[:@123846.4]
  input  [63:0] io_ins_445, // @[:@123846.4]
  input  [63:0] io_ins_446, // @[:@123846.4]
  input  [63:0] io_ins_447, // @[:@123846.4]
  input  [63:0] io_ins_448, // @[:@123846.4]
  input  [63:0] io_ins_449, // @[:@123846.4]
  input  [63:0] io_ins_450, // @[:@123846.4]
  input  [63:0] io_ins_451, // @[:@123846.4]
  input  [63:0] io_ins_452, // @[:@123846.4]
  input  [63:0] io_ins_453, // @[:@123846.4]
  input  [63:0] io_ins_454, // @[:@123846.4]
  input  [63:0] io_ins_455, // @[:@123846.4]
  input  [63:0] io_ins_456, // @[:@123846.4]
  input  [63:0] io_ins_457, // @[:@123846.4]
  input  [63:0] io_ins_458, // @[:@123846.4]
  input  [63:0] io_ins_459, // @[:@123846.4]
  input  [63:0] io_ins_460, // @[:@123846.4]
  input  [63:0] io_ins_461, // @[:@123846.4]
  input  [63:0] io_ins_462, // @[:@123846.4]
  input  [63:0] io_ins_463, // @[:@123846.4]
  input  [63:0] io_ins_464, // @[:@123846.4]
  input  [63:0] io_ins_465, // @[:@123846.4]
  input  [63:0] io_ins_466, // @[:@123846.4]
  input  [63:0] io_ins_467, // @[:@123846.4]
  input  [63:0] io_ins_468, // @[:@123846.4]
  input  [63:0] io_ins_469, // @[:@123846.4]
  input  [63:0] io_ins_470, // @[:@123846.4]
  input  [63:0] io_ins_471, // @[:@123846.4]
  input  [63:0] io_ins_472, // @[:@123846.4]
  input  [63:0] io_ins_473, // @[:@123846.4]
  input  [63:0] io_ins_474, // @[:@123846.4]
  input  [63:0] io_ins_475, // @[:@123846.4]
  input  [63:0] io_ins_476, // @[:@123846.4]
  input  [63:0] io_ins_477, // @[:@123846.4]
  input  [63:0] io_ins_478, // @[:@123846.4]
  input  [63:0] io_ins_479, // @[:@123846.4]
  input  [63:0] io_ins_480, // @[:@123846.4]
  input  [63:0] io_ins_481, // @[:@123846.4]
  input  [63:0] io_ins_482, // @[:@123846.4]
  input  [63:0] io_ins_483, // @[:@123846.4]
  input  [63:0] io_ins_484, // @[:@123846.4]
  input  [63:0] io_ins_485, // @[:@123846.4]
  input  [63:0] io_ins_486, // @[:@123846.4]
  input  [63:0] io_ins_487, // @[:@123846.4]
  input  [63:0] io_ins_488, // @[:@123846.4]
  input  [63:0] io_ins_489, // @[:@123846.4]
  input  [63:0] io_ins_490, // @[:@123846.4]
  input  [63:0] io_ins_491, // @[:@123846.4]
  input  [63:0] io_ins_492, // @[:@123846.4]
  input  [63:0] io_ins_493, // @[:@123846.4]
  input  [63:0] io_ins_494, // @[:@123846.4]
  input  [63:0] io_ins_495, // @[:@123846.4]
  input  [63:0] io_ins_496, // @[:@123846.4]
  input  [63:0] io_ins_497, // @[:@123846.4]
  input  [63:0] io_ins_498, // @[:@123846.4]
  input  [63:0] io_ins_499, // @[:@123846.4]
  input  [63:0] io_ins_500, // @[:@123846.4]
  input  [63:0] io_ins_501, // @[:@123846.4]
  input  [63:0] io_ins_502, // @[:@123846.4]
  input  [8:0]  io_sel, // @[:@123846.4]
  output [63:0] io_out // @[:@123846.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@123848.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@123848.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@123848.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@123848.4]
endmodule
module RegFile( // @[:@123850.2]
  input         clock, // @[:@123851.4]
  input         reset, // @[:@123852.4]
  input  [31:0] io_raddr, // @[:@123853.4]
  input         io_wen, // @[:@123853.4]
  input  [31:0] io_waddr, // @[:@123853.4]
  input  [63:0] io_wdata, // @[:@123853.4]
  output [63:0] io_rdata, // @[:@123853.4]
  input         io_reset, // @[:@123853.4]
  output [63:0] io_argIns_0, // @[:@123853.4]
  output [63:0] io_argIns_1, // @[:@123853.4]
  output [63:0] io_argIns_2, // @[:@123853.4]
  output [63:0] io_argIns_3, // @[:@123853.4]
  input         io_argOuts_0_valid, // @[:@123853.4]
  input  [63:0] io_argOuts_0_bits, // @[:@123853.4]
  input         io_argOuts_1_valid, // @[:@123853.4]
  input  [63:0] io_argOuts_1_bits // @[:@123853.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@125863.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@125863.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@125863.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@125863.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@125863.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@125863.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@125875.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@125875.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@125875.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@125875.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@125875.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@125875.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@125894.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@125894.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@125894.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@125894.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@125894.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@125894.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@125906.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@125906.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@125906.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@125906.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@125906.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@125906.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@125918.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@125918.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@125918.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@125918.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@125918.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@125918.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@125932.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@125932.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@125932.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@125932.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@125932.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@125932.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@125946.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@125946.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@125946.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@125946.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@125946.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@125946.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@125960.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@125960.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@125960.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@125960.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@125960.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@125960.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@125974.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@125974.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@125974.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@125974.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@125974.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@125974.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@125988.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@125988.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@125988.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@125988.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@125988.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@125988.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@126002.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@126002.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@126002.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@126002.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@126002.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@126002.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@126016.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@126016.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@126016.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@126016.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@126016.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@126016.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@126030.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@126030.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@126030.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@126030.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@126030.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@126030.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@126044.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@126044.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@126044.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@126044.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@126044.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@126044.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@126058.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@126058.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@126058.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@126058.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@126058.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@126058.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@126072.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@126072.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@126072.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@126072.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@126072.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@126072.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@126086.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@126086.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@126086.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@126086.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@126086.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@126086.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@126100.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@126100.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@126100.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@126100.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@126100.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@126100.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@126114.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@126114.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@126114.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@126114.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@126114.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@126114.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@126128.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@126128.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@126128.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@126128.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@126128.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@126128.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@126142.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@126142.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@126142.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@126142.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@126142.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@126142.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@126156.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@126156.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@126156.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@126156.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@126156.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@126156.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@126170.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@126170.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@126170.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@126170.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@126170.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@126170.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@126184.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@126184.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@126184.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@126184.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@126184.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@126184.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@126198.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@126198.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@126198.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@126198.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@126198.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@126198.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@126212.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@126212.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@126212.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@126212.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@126212.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@126212.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@126226.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@126226.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@126226.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@126226.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@126226.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@126226.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@126240.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@126240.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@126240.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@126240.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@126240.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@126240.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@126254.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@126254.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@126254.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@126254.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@126254.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@126254.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@126268.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@126268.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@126268.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@126268.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@126268.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@126268.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@126282.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@126282.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@126282.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@126282.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@126282.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@126282.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@126296.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@126296.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@126296.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@126296.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@126296.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@126296.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@126310.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@126310.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@126310.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@126310.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@126310.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@126310.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@126324.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@126324.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@126324.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@126324.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@126324.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@126324.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@126338.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@126338.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@126338.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@126338.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@126338.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@126338.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@126352.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@126352.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@126352.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@126352.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@126352.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@126352.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@126366.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@126366.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@126366.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@126366.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@126366.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@126366.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@126380.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@126380.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@126380.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@126380.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@126380.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@126380.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@126394.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@126394.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@126394.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@126394.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@126394.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@126394.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@126408.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@126408.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@126408.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@126408.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@126408.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@126408.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@126422.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@126422.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@126422.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@126422.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@126422.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@126422.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@126436.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@126436.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@126436.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@126436.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@126436.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@126436.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@126450.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@126450.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@126450.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@126450.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@126450.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@126450.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@126464.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@126464.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@126464.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@126464.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@126464.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@126464.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@126478.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@126478.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@126478.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@126478.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@126478.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@126478.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@126492.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@126492.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@126492.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@126492.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@126492.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@126492.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@126506.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@126506.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@126506.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@126506.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@126506.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@126506.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@126520.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@126520.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@126520.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@126520.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@126520.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@126520.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@126534.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@126534.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@126534.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@126534.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@126534.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@126534.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@126548.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@126548.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@126548.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@126548.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@126548.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@126548.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@126562.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@126562.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@126562.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@126562.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@126562.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@126562.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@126576.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@126576.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@126576.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@126576.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@126576.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@126576.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@126590.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@126590.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@126590.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@126590.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@126590.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@126590.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@126604.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@126604.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@126604.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@126604.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@126604.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@126604.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@126618.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@126618.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@126618.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@126618.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@126618.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@126618.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@126632.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@126632.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@126632.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@126632.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@126632.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@126632.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@126646.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@126646.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@126646.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@126646.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@126646.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@126646.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@126660.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@126660.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@126660.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@126660.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@126660.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@126660.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@126674.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@126674.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@126674.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@126674.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@126674.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@126674.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@126688.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@126688.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@126688.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@126688.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@126688.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@126688.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@126702.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@126702.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@126702.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@126702.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@126702.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@126702.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@126716.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@126716.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@126716.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@126716.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@126716.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@126716.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@126730.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@126730.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@126730.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@126730.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@126730.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@126730.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@126744.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@126744.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@126744.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@126744.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@126744.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@126744.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@126758.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@126758.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@126758.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@126758.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@126758.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@126758.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@126772.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@126772.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@126772.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@126772.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@126772.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@126772.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@126786.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@126786.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@126786.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@126786.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@126786.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@126786.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@126800.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@126800.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@126800.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@126800.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@126800.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@126800.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@126814.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@126814.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@126814.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@126814.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@126814.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@126814.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@126828.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@126828.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@126828.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@126828.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@126828.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@126828.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@126842.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@126842.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@126842.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@126842.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@126842.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@126842.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@126856.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@126856.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@126856.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@126856.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@126856.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@126856.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@126870.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@126870.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@126870.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@126870.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@126870.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@126870.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@126884.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@126884.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@126884.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@126884.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@126884.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@126884.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@126898.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@126898.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@126898.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@126898.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@126898.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@126898.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@126912.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@126912.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@126912.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@126926.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@126926.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@126926.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@126926.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@126926.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@126926.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@126940.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@126940.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@126954.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@126954.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@126954.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@126954.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@126954.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@126954.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@126968.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@126968.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@126968.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@126968.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@126968.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@126968.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@126982.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@126982.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@126982.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@126982.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@126982.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@126982.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@126996.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@126996.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@126996.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@126996.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@126996.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@126996.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@127010.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@127010.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@127010.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@127010.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@127010.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@127010.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@127024.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@127024.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@127024.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@127024.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@127024.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@127024.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@127038.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@127038.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@127038.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@127038.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@127038.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@127038.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@127052.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@127052.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@127052.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@127052.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@127052.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@127052.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@127066.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@127066.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@127066.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@127066.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@127066.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@127066.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@127080.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@127080.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@127080.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@127080.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@127080.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@127080.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@127094.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@127094.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@127094.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@127094.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@127094.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@127094.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@127108.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@127108.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@127108.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@127108.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@127108.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@127108.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@127122.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@127122.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@127122.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@127122.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@127122.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@127122.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@127136.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@127136.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@127136.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@127136.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@127136.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@127136.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@127150.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@127150.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@127150.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@127150.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@127150.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@127150.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@127164.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@127164.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@127164.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@127164.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@127164.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@127164.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@127178.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@127178.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@127178.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@127178.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@127178.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@127178.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@127192.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@127192.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@127192.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@127192.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@127192.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@127192.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@127206.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@127206.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@127206.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@127206.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@127206.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@127206.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@127220.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@127220.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@127220.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@127220.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@127220.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@127220.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@127234.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@127234.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@127234.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@127234.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@127234.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@127234.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@127248.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@127248.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@127248.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@127248.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@127248.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@127248.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@127262.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@127262.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@127262.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@127262.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@127262.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@127262.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@127276.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@127276.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@127276.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@127276.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@127276.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@127276.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@127290.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@127290.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@127290.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@127290.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@127290.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@127290.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@127304.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@127304.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@127304.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@127304.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@127304.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@127304.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@127318.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@127318.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@127318.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@127318.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@127318.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@127318.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@127332.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@127332.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@127332.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@127332.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@127332.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@127332.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@127346.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@127346.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@127346.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@127346.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@127346.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@127346.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@127360.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@127360.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@127360.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@127360.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@127360.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@127360.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@127374.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@127374.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@127374.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@127374.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@127374.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@127374.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@127388.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@127388.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@127388.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@127388.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@127388.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@127388.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@127402.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@127402.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@127402.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@127402.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@127402.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@127402.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@127416.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@127416.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@127416.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@127416.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@127416.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@127416.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@127430.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@127430.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@127430.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@127430.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@127430.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@127430.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@127444.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@127444.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@127444.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@127444.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@127444.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@127444.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@127458.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@127458.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@127458.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@127458.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@127458.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@127458.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@127472.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@127472.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@127472.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@127472.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@127472.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@127472.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@127486.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@127486.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@127486.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@127486.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@127486.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@127486.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@127500.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@127500.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@127500.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@127500.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@127500.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@127500.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@127514.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@127514.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@127514.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@127514.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@127514.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@127514.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@127528.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@127528.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@127528.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@127528.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@127528.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@127528.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@127542.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@127542.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@127542.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@127542.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@127542.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@127542.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@127556.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@127556.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@127556.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@127556.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@127556.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@127556.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@127570.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@127570.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@127570.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@127570.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@127570.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@127570.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@127584.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@127584.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@127584.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@127584.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@127584.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@127584.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@127598.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@127598.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@127598.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@127598.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@127598.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@127598.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@127612.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@127612.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@127612.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@127612.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@127612.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@127612.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@127626.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@127626.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@127626.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@127626.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@127626.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@127626.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@127640.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@127640.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@127640.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@127640.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@127640.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@127640.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@127654.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@127654.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@127654.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@127654.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@127654.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@127654.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@127668.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@127668.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@127668.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@127668.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@127668.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@127668.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@127682.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@127682.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@127682.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@127682.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@127682.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@127682.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@127696.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@127696.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@127696.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@127696.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@127696.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@127696.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@127710.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@127710.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@127710.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@127710.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@127710.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@127710.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@127724.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@127724.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@127724.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@127724.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@127724.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@127724.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@127738.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@127738.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@127738.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@127738.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@127738.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@127738.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@127752.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@127752.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@127752.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@127752.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@127752.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@127752.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@127766.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@127766.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@127766.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@127766.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@127766.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@127766.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@127780.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@127780.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@127780.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@127780.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@127780.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@127780.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@127794.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@127794.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@127794.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@127794.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@127794.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@127794.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@127808.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@127808.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@127808.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@127808.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@127808.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@127808.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@127822.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@127822.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@127822.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@127822.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@127822.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@127822.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@127836.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@127836.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@127836.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@127836.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@127836.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@127836.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@127850.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@127850.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@127850.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@127850.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@127850.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@127850.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@127864.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@127864.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@127864.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@127864.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@127864.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@127864.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@127878.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@127878.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@127878.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@127878.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@127878.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@127878.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@127892.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@127892.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@127892.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@127892.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@127892.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@127892.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@127906.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@127906.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@127906.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@127906.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@127906.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@127906.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@127920.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@127920.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@127920.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@127920.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@127920.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@127920.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@127934.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@127934.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@127934.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@127934.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@127934.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@127934.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@127948.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@127948.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@127948.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@127948.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@127948.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@127948.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@127962.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@127962.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@127962.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@127962.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@127962.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@127962.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@127976.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@127976.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@127976.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@127976.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@127976.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@127976.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@127990.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@127990.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@127990.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@127990.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@127990.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@127990.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@128004.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@128004.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@128004.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@128004.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@128004.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@128004.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@128018.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@128018.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@128018.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@128018.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@128018.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@128018.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@128032.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@128032.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@128032.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@128032.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@128032.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@128032.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@128046.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@128046.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@128046.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@128046.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@128046.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@128046.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@128060.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@128060.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@128060.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@128060.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@128060.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@128060.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@128074.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@128074.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@128074.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@128074.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@128074.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@128074.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@128088.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@128088.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@128088.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@128088.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@128088.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@128088.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@128102.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@128102.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@128102.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@128102.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@128102.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@128102.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@128116.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@128116.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@128116.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@128116.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@128116.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@128116.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@128130.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@128130.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@128130.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@128130.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@128130.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@128130.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@128144.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@128144.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@128144.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@128144.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@128144.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@128144.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@128158.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@128158.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@128158.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@128158.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@128158.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@128158.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@128172.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@128172.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@128172.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@128172.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@128172.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@128172.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@128186.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@128186.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@128186.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@128186.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@128186.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@128186.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@128200.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@128200.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@128200.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@128200.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@128200.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@128200.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@128214.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@128214.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@128214.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@128214.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@128214.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@128214.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@128228.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@128228.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@128228.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@128228.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@128228.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@128228.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@128242.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@128242.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@128242.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@128242.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@128242.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@128242.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@128256.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@128256.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@128256.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@128256.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@128256.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@128256.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@128270.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@128270.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@128270.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@128270.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@128270.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@128270.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@128284.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@128284.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@128284.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@128284.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@128284.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@128284.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@128298.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@128298.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@128298.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@128298.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@128298.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@128298.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@128312.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@128312.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@128312.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@128312.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@128312.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@128312.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@128326.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@128326.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@128326.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@128326.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@128326.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@128326.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@128340.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@128340.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@128340.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@128340.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@128340.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@128340.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@128354.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@128354.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@128354.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@128354.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@128354.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@128354.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@128368.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@128368.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@128368.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@128368.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@128368.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@128368.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@128382.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@128382.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@128382.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@128382.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@128382.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@128382.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@128396.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@128396.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@128396.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@128396.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@128396.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@128396.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@128410.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@128410.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@128410.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@128410.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@128410.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@128410.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@128424.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@128424.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@128424.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@128424.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@128424.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@128424.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@128438.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@128438.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@128438.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@128438.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@128438.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@128438.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@128452.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@128452.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@128452.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@128452.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@128452.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@128452.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@128466.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@128466.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@128466.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@128466.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@128466.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@128466.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@128480.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@128480.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@128480.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@128480.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@128480.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@128480.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@128494.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@128494.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@128494.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@128494.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@128494.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@128494.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@128508.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@128508.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@128508.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@128508.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@128508.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@128508.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@128522.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@128522.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@128522.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@128522.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@128522.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@128522.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@128536.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@128536.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@128536.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@128536.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@128536.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@128536.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@128550.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@128550.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@128550.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@128550.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@128550.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@128550.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@128564.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@128564.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@128564.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@128564.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@128564.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@128564.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@128578.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@128578.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@128578.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@128578.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@128578.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@128578.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@128592.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@128592.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@128592.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@128592.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@128592.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@128592.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@128606.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@128606.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@128606.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@128606.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@128606.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@128606.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@128620.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@128620.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@128620.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@128620.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@128620.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@128620.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@128634.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@128634.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@128634.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@128634.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@128634.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@128634.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@128648.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@128648.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@128648.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@128648.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@128648.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@128648.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@128662.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@128662.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@128662.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@128662.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@128662.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@128662.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@128676.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@128676.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@128676.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@128676.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@128676.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@128676.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@128690.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@128690.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@128690.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@128690.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@128690.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@128690.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@128704.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@128704.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@128704.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@128704.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@128704.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@128704.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@128718.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@128718.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@128718.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@128718.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@128718.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@128718.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@128732.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@128732.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@128732.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@128732.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@128732.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@128732.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@128746.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@128746.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@128746.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@128746.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@128746.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@128746.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@128760.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@128760.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@128760.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@128760.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@128760.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@128760.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@128774.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@128774.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@128774.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@128774.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@128774.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@128774.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@128788.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@128788.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@128788.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@128788.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@128788.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@128788.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@128802.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@128802.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@128802.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@128802.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@128802.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@128802.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@128816.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@128816.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@128816.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@128816.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@128816.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@128816.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@128830.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@128830.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@128830.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@128830.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@128830.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@128830.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@128844.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@128844.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@128844.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@128844.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@128844.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@128844.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@128858.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@128858.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@128858.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@128858.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@128858.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@128858.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@128872.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@128872.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@128872.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@128872.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@128872.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@128872.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@128886.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@128886.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@128886.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@128886.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@128886.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@128886.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@128900.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@128900.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@128900.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@128900.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@128900.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@128900.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@128914.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@128914.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@128914.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@128914.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@128914.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@128914.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@128928.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@128928.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@128928.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@128928.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@128928.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@128928.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@128942.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@128942.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@128942.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@128942.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@128942.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@128942.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@128956.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@128956.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@128956.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@128956.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@128956.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@128956.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@128970.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@128970.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@128970.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@128970.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@128970.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@128970.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@128984.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@128984.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@128984.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@128984.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@128984.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@128984.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@128998.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@128998.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@128998.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@128998.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@128998.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@128998.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@129012.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@129012.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@129012.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@129012.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@129012.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@129012.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@129026.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@129026.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@129026.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@129026.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@129026.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@129026.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@129040.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@129040.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@129040.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@129040.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@129040.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@129040.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@129054.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@129054.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@129054.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@129054.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@129054.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@129054.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@129068.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@129068.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@129068.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@129068.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@129068.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@129068.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@129082.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@129082.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@129082.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@129082.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@129082.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@129082.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@129096.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@129096.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@129096.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@129096.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@129096.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@129096.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@129110.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@129110.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@129110.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@129110.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@129110.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@129110.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@129124.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@129124.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@129124.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@129124.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@129124.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@129124.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@129138.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@129138.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@129138.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@129138.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@129138.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@129138.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@129152.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@129152.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@129152.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@129152.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@129152.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@129152.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@129166.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@129166.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@129166.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@129166.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@129166.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@129166.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@129180.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@129180.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@129180.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@129180.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@129180.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@129180.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@129194.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@129194.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@129194.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@129194.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@129194.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@129194.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@129208.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@129208.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@129208.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@129208.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@129208.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@129208.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@129222.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@129222.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@129222.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@129222.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@129222.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@129222.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@129236.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@129236.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@129236.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@129236.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@129236.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@129236.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@129250.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@129250.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@129250.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@129250.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@129250.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@129250.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@129264.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@129264.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@129264.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@129264.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@129264.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@129264.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@129278.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@129278.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@129278.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@129278.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@129278.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@129278.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@129292.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@129292.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@129292.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@129292.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@129292.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@129292.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@129306.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@129306.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@129306.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@129306.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@129306.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@129306.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@129320.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@129320.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@129320.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@129320.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@129320.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@129320.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@129334.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@129334.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@129334.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@129334.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@129334.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@129334.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@129348.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@129348.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@129348.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@129348.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@129348.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@129348.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@129362.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@129362.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@129362.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@129362.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@129362.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@129362.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@129376.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@129376.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@129376.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@129376.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@129376.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@129376.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@129390.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@129390.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@129390.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@129390.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@129390.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@129390.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@129404.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@129404.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@129404.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@129404.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@129404.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@129404.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@129418.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@129418.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@129418.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@129418.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@129418.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@129418.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@129432.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@129432.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@129432.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@129432.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@129432.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@129432.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@129446.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@129446.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@129446.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@129446.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@129446.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@129446.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@129460.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@129460.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@129460.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@129460.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@129460.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@129460.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@129474.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@129474.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@129474.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@129474.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@129474.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@129474.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@129488.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@129488.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@129488.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@129488.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@129488.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@129488.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@129502.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@129502.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@129502.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@129502.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@129502.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@129502.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@129516.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@129516.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@129516.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@129516.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@129516.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@129516.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@129530.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@129530.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@129530.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@129530.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@129530.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@129530.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@129544.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@129544.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@129544.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@129544.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@129544.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@129544.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@129558.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@129558.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@129558.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@129558.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@129558.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@129558.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@129572.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@129572.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@129572.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@129572.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@129572.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@129572.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@129586.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@129586.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@129586.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@129586.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@129586.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@129586.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@129600.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@129600.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@129600.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@129600.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@129600.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@129600.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@129614.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@129614.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@129614.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@129614.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@129614.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@129614.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@129628.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@129628.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@129628.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@129628.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@129628.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@129628.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@129642.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@129642.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@129642.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@129642.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@129642.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@129642.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@129656.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@129656.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@129656.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@129656.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@129656.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@129656.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@129670.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@129670.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@129670.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@129670.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@129670.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@129670.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@129684.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@129684.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@129684.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@129684.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@129684.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@129684.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@129698.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@129698.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@129698.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@129698.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@129698.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@129698.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@129712.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@129712.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@129712.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@129712.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@129712.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@129712.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@129726.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@129726.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@129726.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@129726.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@129726.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@129726.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@129740.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@129740.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@129740.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@129740.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@129740.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@129740.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@129754.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@129754.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@129754.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@129754.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@129754.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@129754.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@129768.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@129768.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@129768.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@129768.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@129768.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@129768.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@129782.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@129782.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@129782.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@129782.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@129782.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@129782.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@129796.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@129796.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@129796.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@129796.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@129796.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@129796.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@129810.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@129810.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@129810.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@129810.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@129810.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@129810.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@129824.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@129824.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@129824.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@129824.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@129824.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@129824.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@129838.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@129838.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@129838.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@129838.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@129838.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@129838.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@129852.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@129852.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@129852.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@129852.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@129852.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@129852.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@129866.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@129866.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@129866.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@129866.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@129866.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@129866.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@129880.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@129880.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@129880.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@129880.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@129880.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@129880.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@129894.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@129894.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@129894.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@129894.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@129894.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@129894.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@129908.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@129908.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@129908.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@129908.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@129908.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@129908.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@129922.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@129922.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@129922.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@129922.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@129922.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@129922.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@129936.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@129936.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@129936.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@129936.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@129936.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@129936.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@129950.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@129950.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@129950.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@129950.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@129950.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@129950.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@129964.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@129964.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@129964.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@129964.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@129964.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@129964.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@129978.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@129978.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@129978.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@129978.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@129978.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@129978.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@129992.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@129992.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@129992.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@129992.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@129992.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@129992.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@130006.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@130006.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@130006.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@130006.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@130006.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@130006.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@130020.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@130020.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@130020.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@130020.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@130020.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@130020.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@130034.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@130034.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@130034.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@130034.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@130034.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@130034.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@130048.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@130048.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@130048.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@130048.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@130048.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@130048.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@130062.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@130062.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@130062.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@130062.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@130062.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@130062.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@130076.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@130076.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@130076.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@130076.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@130076.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@130076.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@130090.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@130090.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@130090.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@130090.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@130090.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@130090.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@130104.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@130104.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@130104.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@130104.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@130104.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@130104.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@130118.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@130118.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@130118.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@130118.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@130118.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@130118.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@130132.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@130132.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@130132.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@130132.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@130132.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@130132.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@130146.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@130146.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@130146.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@130146.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@130146.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@130146.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@130160.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@130160.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@130160.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@130160.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@130160.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@130160.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@130174.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@130174.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@130174.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@130174.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@130174.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@130174.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@130188.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@130188.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@130188.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@130188.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@130188.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@130188.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@130202.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@130202.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@130202.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@130202.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@130202.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@130202.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@130216.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@130216.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@130216.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@130216.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@130216.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@130216.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@130230.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@130230.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@130230.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@130230.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@130230.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@130230.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@130244.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@130244.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@130244.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@130244.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@130244.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@130244.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@130258.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@130258.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@130258.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@130258.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@130258.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@130258.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@130272.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@130272.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@130272.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@130272.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@130272.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@130272.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@130286.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@130286.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@130286.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@130286.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@130286.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@130286.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@130300.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@130300.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@130300.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@130300.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@130300.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@130300.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@130314.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@130314.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@130314.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@130314.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@130314.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@130314.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@130328.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@130328.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@130328.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@130328.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@130328.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@130328.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@130342.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@130342.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@130342.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@130342.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@130342.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@130342.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@130356.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@130356.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@130356.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@130356.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@130356.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@130356.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@130370.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@130370.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@130370.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@130370.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@130370.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@130370.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@130384.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@130384.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@130384.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@130384.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@130384.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@130384.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@130398.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@130398.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@130398.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@130398.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@130398.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@130398.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@130412.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@130412.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@130412.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@130412.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@130412.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@130412.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@130426.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@130426.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@130426.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@130426.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@130426.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@130426.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@130440.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@130440.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@130440.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@130440.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@130440.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@130440.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@130454.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@130454.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@130454.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@130454.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@130454.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@130454.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@130468.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@130468.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@130468.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@130468.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@130468.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@130468.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@130482.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@130482.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@130482.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@130482.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@130482.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@130482.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@130496.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@130496.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@130496.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@130496.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@130496.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@130496.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@130510.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@130510.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@130510.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@130510.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@130510.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@130510.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@130524.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@130524.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@130524.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@130524.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@130524.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@130524.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@130538.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@130538.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@130538.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@130538.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@130538.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@130538.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@130552.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@130552.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@130552.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@130552.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@130552.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@130552.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@130566.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@130566.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@130566.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@130566.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@130566.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@130566.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@130580.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@130580.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@130580.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@130580.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@130580.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@130580.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@130594.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@130594.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@130594.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@130594.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@130594.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@130594.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@130608.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@130608.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@130608.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@130608.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@130608.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@130608.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@130622.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@130622.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@130622.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@130622.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@130622.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@130622.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@130636.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@130636.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@130636.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@130636.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@130636.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@130636.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@130650.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@130650.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@130650.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@130650.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@130650.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@130650.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@130664.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@130664.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@130664.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@130664.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@130664.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@130664.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@130678.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@130678.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@130678.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@130678.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@130678.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@130678.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@130692.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@130692.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@130692.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@130692.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@130692.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@130692.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@130706.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@130706.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@130706.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@130706.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@130706.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@130706.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@130720.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@130720.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@130720.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@130720.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@130720.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@130720.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@130734.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@130734.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@130734.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@130734.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@130734.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@130734.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@130748.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@130748.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@130748.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@130748.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@130748.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@130748.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@130762.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@130762.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@130762.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@130762.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@130762.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@130762.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@130776.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@130776.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@130776.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@130776.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@130776.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@130776.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@130790.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@130790.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@130790.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@130790.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@130790.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@130790.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@130804.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@130804.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@130804.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@130804.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@130804.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@130804.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@130818.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@130818.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@130818.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@130818.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@130818.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@130818.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@130832.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@130832.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@130832.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@130832.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@130832.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@130832.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@130846.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@130846.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@130846.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@130846.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@130846.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@130846.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@130860.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@130860.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@130860.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@130860.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@130860.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@130860.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@130874.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@130874.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@130874.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@130874.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@130874.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@130874.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@130888.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@130888.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@130888.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@130888.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@130888.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@130888.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@130902.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@130902.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@130902.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@130902.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@130902.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@130902.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@130916.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@130916.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@130916.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@130916.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@130916.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@130916.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@130930.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@130930.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@130930.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@130930.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@130930.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@130930.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@130944.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@130944.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@130944.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@130944.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@130944.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@130944.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@130958.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@130958.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@130958.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@130958.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@130958.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@130958.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@130972.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@130972.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@130972.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@130972.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@130972.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@130972.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@130986.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@130986.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@130986.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@130986.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@130986.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@130986.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@131000.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@131000.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@131000.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@131000.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@131000.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@131000.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@131014.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@131014.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@131014.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@131014.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@131014.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@131014.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@131028.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@131028.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@131028.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@131028.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@131028.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@131028.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@131042.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@131042.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@131042.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@131042.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@131042.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@131042.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@131056.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@131056.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@131056.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@131056.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@131056.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@131056.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@131070.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@131070.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@131070.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@131070.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@131070.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@131070.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@131084.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@131084.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@131084.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@131084.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@131084.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@131084.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@131098.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@131098.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@131098.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@131098.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@131098.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@131098.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@131112.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@131112.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@131112.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@131112.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@131112.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@131112.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@131126.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@131126.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@131126.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@131126.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@131126.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@131126.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@131140.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@131140.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@131140.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@131140.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@131140.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@131140.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@131154.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@131154.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@131154.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@131154.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@131154.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@131154.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@131168.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@131168.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@131168.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@131168.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@131168.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@131168.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@131182.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@131182.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@131182.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@131182.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@131182.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@131182.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@131196.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@131196.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@131196.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@131196.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@131196.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@131196.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@131210.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@131210.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@131210.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@131210.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@131210.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@131210.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@131224.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@131224.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@131224.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@131224.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@131224.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@131224.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@131238.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@131238.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@131238.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@131238.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@131238.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@131238.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@131252.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@131252.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@131252.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@131252.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@131252.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@131252.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@131266.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@131266.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@131266.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@131266.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@131266.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@131266.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@131280.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@131280.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@131280.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@131280.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@131280.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@131280.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@131294.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@131294.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@131294.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@131294.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@131294.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@131294.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@131308.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@131308.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@131308.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@131308.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@131308.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@131308.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@131322.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@131322.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@131322.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@131322.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@131322.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@131322.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@131336.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@131336.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@131336.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@131336.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@131336.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@131336.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@131350.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@131350.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@131350.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@131350.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@131350.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@131350.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@131364.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@131364.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@131364.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@131364.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@131364.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@131364.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@131378.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@131378.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@131378.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@131378.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@131378.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@131378.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@131392.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@131392.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@131392.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@131392.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@131392.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@131392.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@131406.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@131406.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@131406.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@131406.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@131406.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@131406.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@131420.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@131420.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@131420.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@131420.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@131420.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@131420.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@131434.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@131434.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@131434.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@131434.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@131434.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@131434.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@131448.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@131448.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@131448.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@131448.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@131448.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@131448.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@131462.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@131462.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@131462.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@131462.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@131462.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@131462.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@131476.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@131476.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@131476.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@131476.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@131476.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@131476.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@131490.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@131490.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@131490.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@131490.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@131490.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@131490.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@131504.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@131504.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@131504.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@131504.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@131504.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@131504.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@131518.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@131518.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@131518.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@131518.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@131518.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@131518.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@131532.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@131532.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@131532.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@131532.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@131532.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@131532.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@131546.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@131546.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@131546.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@131546.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@131546.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@131546.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@131560.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@131560.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@131560.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@131560.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@131560.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@131560.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@131574.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@131574.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@131574.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@131574.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@131574.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@131574.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@131588.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@131588.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@131588.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@131588.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@131588.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@131588.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@131602.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@131602.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@131602.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@131602.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@131602.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@131602.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@131616.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@131616.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@131616.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@131616.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@131616.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@131616.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@131630.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@131630.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@131630.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@131630.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@131630.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@131630.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@131644.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@131644.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@131644.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@131644.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@131644.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@131644.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@131658.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@131658.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@131658.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@131658.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@131658.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@131658.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@131672.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@131672.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@131672.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@131672.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@131672.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@131672.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@131686.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@131686.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@131686.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@131686.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@131686.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@131686.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@131700.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@131700.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@131700.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@131700.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@131700.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@131700.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@131714.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@131714.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@131714.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@131714.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@131714.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@131714.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@131728.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@131728.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@131728.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@131728.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@131728.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@131728.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@131742.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@131742.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@131742.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@131742.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@131742.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@131742.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@131756.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@131756.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@131756.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@131756.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@131756.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@131756.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@131770.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@131770.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@131770.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@131770.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@131770.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@131770.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@131784.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@131784.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@131784.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@131784.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@131784.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@131784.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@131798.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@131798.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@131798.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@131798.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@131798.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@131798.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@131812.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@131812.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@131812.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@131812.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@131812.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@131812.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@131826.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@131826.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@131826.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@131826.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@131826.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@131826.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@131840.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@131840.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@131840.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@131840.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@131840.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@131840.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@131854.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@131854.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@131854.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@131854.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@131854.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@131854.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@131868.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@131868.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@131868.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@131868.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@131868.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@131868.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@131882.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@131882.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@131882.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@131882.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@131882.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@131882.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@131896.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@131896.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@131896.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@131896.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@131896.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@131896.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@131910.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@131910.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@131910.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@131910.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@131910.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@131910.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@131924.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@131924.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@131924.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@131924.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@131924.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@131924.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@131938.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@131938.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@131938.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@131938.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@131938.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@131938.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@131952.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@131952.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@131952.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@131952.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@131952.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@131952.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@131966.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@131966.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@131966.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@131966.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@131966.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@131966.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@131980.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@131980.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@131980.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@131980.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@131980.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@131980.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@131994.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@131994.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@131994.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@131994.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@131994.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@131994.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@132008.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@132008.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@132008.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@132008.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@132008.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@132008.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@132022.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@132022.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@132022.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@132022.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@132022.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@132022.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@132036.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@132036.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@132036.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@132036.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@132036.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@132036.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@132050.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@132050.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@132050.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@132050.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@132050.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@132050.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@132064.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@132064.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@132064.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@132064.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@132064.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@132064.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@132078.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@132078.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@132078.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@132078.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@132078.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@132078.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@132092.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@132092.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@132092.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@132092.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@132092.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@132092.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@132106.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@132106.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@132106.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@132106.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@132106.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@132106.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@132120.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@132120.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@132120.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@132120.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@132120.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@132120.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@132134.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@132134.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@132134.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@132134.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@132134.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@132134.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@132148.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@132148.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@132148.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@132148.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@132148.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@132148.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@132162.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@132162.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@132162.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@132162.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@132162.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@132162.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@132176.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@132176.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@132176.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@132176.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@132176.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@132176.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@132190.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@132190.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@132190.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@132190.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@132190.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@132190.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@132204.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@132204.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@132204.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@132204.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@132204.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@132204.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@132218.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@132218.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@132218.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@132218.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@132218.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@132218.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@132232.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@132232.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@132232.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@132232.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@132232.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@132232.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@132246.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@132246.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@132246.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@132246.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@132246.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@132246.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@132260.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@132260.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@132260.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@132260.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@132260.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@132260.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@132274.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@132274.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@132274.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@132274.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@132274.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@132274.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@132288.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@132288.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@132288.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@132288.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@132288.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@132288.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@132302.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@132302.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@132302.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@132302.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@132302.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@132302.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@132316.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@132316.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@132316.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@132316.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@132316.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@132316.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@132330.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@132330.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@132330.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@132330.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@132330.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@132330.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@132344.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@132344.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@132344.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@132344.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@132344.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@132344.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@132358.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@132358.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@132358.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@132358.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@132358.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@132358.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@132372.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@132372.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@132372.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@132372.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@132372.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@132372.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@132386.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@132386.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@132386.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@132386.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@132386.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@132386.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@132400.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@132400.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@132400.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@132400.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@132400.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@132400.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@132414.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@132414.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@132414.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@132414.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@132414.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@132414.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@132428.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@132428.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@132428.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@132428.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@132428.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@132428.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@132442.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@132442.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@132442.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@132442.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@132442.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@132442.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@132456.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@132456.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@132456.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@132456.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@132456.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@132456.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@132470.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@132470.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@132470.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@132470.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@132470.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@132470.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@132484.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@132484.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@132484.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@132484.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@132484.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@132484.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@132498.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@132498.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@132498.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@132498.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@132498.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@132498.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@132512.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@132512.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@132512.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@132512.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@132512.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@132512.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@132526.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@132526.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@132526.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@132526.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@132526.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@132526.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@132540.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@132540.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@132540.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@132540.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@132540.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@132540.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@132554.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@132554.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@132554.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@132554.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@132554.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@132554.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@132568.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@132568.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@132568.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@132568.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@132568.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@132568.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@132582.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@132582.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@132582.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@132582.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@132582.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@132582.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@132596.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@132596.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@132596.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@132596.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@132596.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@132596.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@132610.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@132610.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@132610.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@132610.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@132610.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@132610.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@132624.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@132624.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@132624.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@132624.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@132624.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@132624.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@132638.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@132638.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@132638.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@132638.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@132638.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@132638.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@132652.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@132652.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@132652.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@132652.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@132652.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@132652.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@132666.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@132666.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@132666.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@132666.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@132666.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@132666.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@132680.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@132680.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@132680.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@132680.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@132680.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@132680.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@132694.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@132694.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@132694.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@132694.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@132694.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@132694.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@132708.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@132708.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@132708.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@132708.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@132708.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@132708.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@132722.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@132722.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@132722.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@132722.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@132722.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@132722.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@132736.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@132736.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@132736.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@132736.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@132736.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@132736.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@132750.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@132750.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@132750.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@132750.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@132750.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@132750.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@132764.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@132764.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@132764.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@132764.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@132764.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@132764.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@132778.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@132778.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@132778.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@132792.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@132792.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@132792.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@132806.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@132806.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@132806.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@132820.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@132820.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@132820.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@132834.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@132834.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@132834.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@132848.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@132848.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@132848.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@132862.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@132862.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@132862.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@132876.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@132876.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@132876.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@132890.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@132890.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@132890.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@132890.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@132904.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@132904.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@132904.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@125866.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@125878.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@125879.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@125897.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@125909.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@125921.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@125922.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@125863.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@125875.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@125894.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@125906.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@125918.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@125932.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@125946.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@125960.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@125974.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@125988.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@126002.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@126016.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@126030.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@126044.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@126058.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@126072.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@126086.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@126100.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@126114.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@126128.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@126142.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@126156.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@126170.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@126184.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@126198.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@126212.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@126226.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@126240.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@126254.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@126268.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@126282.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@126296.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@126310.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@126324.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@126338.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@126352.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@126366.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@126380.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@126394.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@126408.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@126422.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@126436.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@126450.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@126464.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@126478.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@126492.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@126506.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@126520.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@126534.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@126548.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@126562.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@126576.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@126590.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@126604.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@126618.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@126632.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@126646.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@126660.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@126674.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@126688.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@126702.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@126716.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@126730.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@126744.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@126758.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@126772.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@126786.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@126800.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@126814.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@126828.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@126842.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@126856.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@126870.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@126884.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@126898.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@126912.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@126926.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@126940.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@126954.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@126968.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@126982.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@126996.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@127010.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@127024.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@127038.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@127052.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@127066.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@127080.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@127094.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@127108.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@127122.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@127136.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@127150.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@127164.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@127178.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@127192.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@127206.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@127220.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@127234.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@127248.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@127262.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@127276.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@127290.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@127304.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@127318.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@127332.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@127346.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@127360.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@127374.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@127388.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@127402.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@127416.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@127430.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@127444.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@127458.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@127472.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@127486.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@127500.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@127514.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@127528.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@127542.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@127556.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@127570.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@127584.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@127598.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@127612.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@127626.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@127640.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@127654.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@127668.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@127682.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@127696.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@127710.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@127724.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@127738.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@127752.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@127766.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@127780.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@127794.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@127808.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@127822.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@127836.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@127850.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@127864.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@127878.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@127892.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@127906.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@127920.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@127934.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@127948.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@127962.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@127976.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@127990.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@128004.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@128018.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@128032.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@128046.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@128060.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@128074.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@128088.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@128102.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@128116.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@128130.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@128144.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@128158.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@128172.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@128186.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@128200.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@128214.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@128228.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@128242.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@128256.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@128270.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@128284.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@128298.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@128312.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@128326.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@128340.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@128354.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@128368.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@128382.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@128396.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@128410.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@128424.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@128438.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@128452.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@128466.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@128480.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@128494.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@128508.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@128522.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@128536.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@128550.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@128564.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@128578.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@128592.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@128606.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@128620.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@128634.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@128648.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@128662.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@128676.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@128690.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@128704.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@128718.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@128732.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@128746.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@128760.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@128774.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@128788.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@128802.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@128816.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@128830.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@128844.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@128858.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@128872.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@128886.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@128900.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@128914.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@128928.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@128942.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@128956.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@128970.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@128984.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@128998.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@129012.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@129026.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@129040.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@129054.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@129068.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@129082.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@129096.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@129110.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@129124.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@129138.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@129152.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@129166.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@129180.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@129194.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@129208.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@129222.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@129236.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@129250.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@129264.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@129278.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@129292.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@129306.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@129320.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@129334.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@129348.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@129362.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@129376.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@129390.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@129404.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@129418.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@129432.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@129446.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@129460.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@129474.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@129488.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@129502.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@129516.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@129530.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@129544.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@129558.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@129572.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@129586.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@129600.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@129614.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@129628.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@129642.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@129656.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@129670.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@129684.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@129698.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@129712.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@129726.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@129740.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@129754.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@129768.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@129782.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@129796.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@129810.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@129824.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@129838.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@129852.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@129866.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@129880.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@129894.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@129908.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@129922.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@129936.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@129950.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@129964.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@129978.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@129992.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@130006.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@130020.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@130034.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@130048.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@130062.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@130076.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@130090.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@130104.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@130118.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@130132.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@130146.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@130160.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@130174.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@130188.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@130202.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@130216.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@130230.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@130244.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@130258.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@130272.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@130286.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@130300.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@130314.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@130328.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@130342.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@130356.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@130370.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@130384.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@130398.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@130412.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@130426.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@130440.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@130454.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@130468.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@130482.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@130496.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@130510.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@130524.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@130538.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@130552.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@130566.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@130580.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@130594.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@130608.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@130622.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@130636.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@130650.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@130664.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@130678.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@130692.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@130706.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@130720.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@130734.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@130748.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@130762.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@130776.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@130790.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@130804.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@130818.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@130832.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@130846.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@130860.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@130874.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@130888.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@130902.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@130916.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@130930.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@130944.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@130958.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@130972.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@130986.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@131000.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@131014.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@131028.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@131042.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@131056.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@131070.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@131084.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@131098.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@131112.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@131126.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@131140.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@131154.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@131168.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@131182.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@131196.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@131210.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@131224.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@131238.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@131252.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@131266.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@131280.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@131294.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@131308.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@131322.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@131336.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@131350.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@131364.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@131378.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@131392.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@131406.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@131420.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@131434.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@131448.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@131462.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@131476.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@131490.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@131504.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@131518.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@131532.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@131546.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@131560.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@131574.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@131588.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@131602.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@131616.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@131630.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@131644.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@131658.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@131672.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@131686.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@131700.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@131714.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@131728.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@131742.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@131756.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@131770.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@131784.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@131798.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@131812.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@131826.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@131840.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@131854.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@131868.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@131882.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@131896.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@131910.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@131924.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@131938.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@131952.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@131966.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@131980.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@131994.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@132008.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@132022.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@132036.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@132050.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@132064.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@132078.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@132092.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@132106.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@132120.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@132134.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@132148.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@132162.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@132176.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@132190.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@132204.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@132218.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@132232.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@132246.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@132260.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@132274.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@132288.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@132302.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@132316.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@132330.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@132344.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@132358.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@132372.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@132386.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@132400.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@132414.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@132428.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@132442.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@132456.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@132470.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@132484.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@132498.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@132512.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@132526.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@132540.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@132554.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@132568.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@132582.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@132596.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@132610.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@132624.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@132638.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@132652.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@132666.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@132680.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@132694.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@132708.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@132722.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@132736.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@132750.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@132764.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@132778.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@132792.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@132806.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@132820.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@132834.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@132848.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@132862.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@132876.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@132890.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@132904.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@125866.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@125878.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@125879.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@125897.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@125909.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@125921.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@125922.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@133915.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@133921.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@133922.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@133923.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@133924.4]
  assign regs_0_clock = clock; // @[:@125864.4]
  assign regs_0_reset = reset; // @[:@125865.4 RegFile.scala 82:16:@125871.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@125869.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@125873.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@125868.4]
  assign regs_1_clock = clock; // @[:@125876.4]
  assign regs_1_reset = reset; // @[:@125877.4 RegFile.scala 70:16:@125889.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@125887.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@125892.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@125883.4]
  assign regs_2_clock = clock; // @[:@125895.4]
  assign regs_2_reset = reset; // @[:@125896.4 RegFile.scala 82:16:@125902.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@125900.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@125904.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@125899.4]
  assign regs_3_clock = clock; // @[:@125907.4]
  assign regs_3_reset = reset; // @[:@125908.4 RegFile.scala 82:16:@125914.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@125912.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@125916.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@125911.4]
  assign regs_4_clock = clock; // @[:@125919.4]
  assign regs_4_reset = io_reset; // @[:@125920.4 RegFile.scala 76:16:@125927.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@125926.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@125930.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@125924.4]
  assign regs_5_clock = clock; // @[:@125933.4]
  assign regs_5_reset = io_reset; // @[:@125934.4 RegFile.scala 76:16:@125941.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@125940.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@125944.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@125938.4]
  assign regs_6_clock = clock; // @[:@125947.4]
  assign regs_6_reset = io_reset; // @[:@125948.4 RegFile.scala 76:16:@125955.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@125954.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@125958.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@125952.4]
  assign regs_7_clock = clock; // @[:@125961.4]
  assign regs_7_reset = io_reset; // @[:@125962.4 RegFile.scala 76:16:@125969.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@125968.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@125972.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@125966.4]
  assign regs_8_clock = clock; // @[:@125975.4]
  assign regs_8_reset = io_reset; // @[:@125976.4 RegFile.scala 76:16:@125983.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@125982.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@125986.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@125980.4]
  assign regs_9_clock = clock; // @[:@125989.4]
  assign regs_9_reset = io_reset; // @[:@125990.4 RegFile.scala 76:16:@125997.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@125996.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@126000.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@125994.4]
  assign regs_10_clock = clock; // @[:@126003.4]
  assign regs_10_reset = io_reset; // @[:@126004.4 RegFile.scala 76:16:@126011.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@126010.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@126014.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@126008.4]
  assign regs_11_clock = clock; // @[:@126017.4]
  assign regs_11_reset = io_reset; // @[:@126018.4 RegFile.scala 76:16:@126025.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@126024.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@126028.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@126022.4]
  assign regs_12_clock = clock; // @[:@126031.4]
  assign regs_12_reset = io_reset; // @[:@126032.4 RegFile.scala 76:16:@126039.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@126038.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@126042.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@126036.4]
  assign regs_13_clock = clock; // @[:@126045.4]
  assign regs_13_reset = io_reset; // @[:@126046.4 RegFile.scala 76:16:@126053.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@126052.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@126056.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@126050.4]
  assign regs_14_clock = clock; // @[:@126059.4]
  assign regs_14_reset = io_reset; // @[:@126060.4 RegFile.scala 76:16:@126067.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@126066.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@126070.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@126064.4]
  assign regs_15_clock = clock; // @[:@126073.4]
  assign regs_15_reset = io_reset; // @[:@126074.4 RegFile.scala 76:16:@126081.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@126080.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@126084.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@126078.4]
  assign regs_16_clock = clock; // @[:@126087.4]
  assign regs_16_reset = io_reset; // @[:@126088.4 RegFile.scala 76:16:@126095.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@126094.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@126098.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@126092.4]
  assign regs_17_clock = clock; // @[:@126101.4]
  assign regs_17_reset = io_reset; // @[:@126102.4 RegFile.scala 76:16:@126109.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@126108.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@126112.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@126106.4]
  assign regs_18_clock = clock; // @[:@126115.4]
  assign regs_18_reset = io_reset; // @[:@126116.4 RegFile.scala 76:16:@126123.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@126122.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@126126.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@126120.4]
  assign regs_19_clock = clock; // @[:@126129.4]
  assign regs_19_reset = io_reset; // @[:@126130.4 RegFile.scala 76:16:@126137.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@126136.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@126140.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@126134.4]
  assign regs_20_clock = clock; // @[:@126143.4]
  assign regs_20_reset = io_reset; // @[:@126144.4 RegFile.scala 76:16:@126151.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@126150.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@126154.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@126148.4]
  assign regs_21_clock = clock; // @[:@126157.4]
  assign regs_21_reset = io_reset; // @[:@126158.4 RegFile.scala 76:16:@126165.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@126164.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@126168.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@126162.4]
  assign regs_22_clock = clock; // @[:@126171.4]
  assign regs_22_reset = io_reset; // @[:@126172.4 RegFile.scala 76:16:@126179.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@126178.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@126182.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@126176.4]
  assign regs_23_clock = clock; // @[:@126185.4]
  assign regs_23_reset = io_reset; // @[:@126186.4 RegFile.scala 76:16:@126193.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@126192.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@126196.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@126190.4]
  assign regs_24_clock = clock; // @[:@126199.4]
  assign regs_24_reset = io_reset; // @[:@126200.4 RegFile.scala 76:16:@126207.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@126206.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@126210.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@126204.4]
  assign regs_25_clock = clock; // @[:@126213.4]
  assign regs_25_reset = io_reset; // @[:@126214.4 RegFile.scala 76:16:@126221.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@126220.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@126224.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@126218.4]
  assign regs_26_clock = clock; // @[:@126227.4]
  assign regs_26_reset = io_reset; // @[:@126228.4 RegFile.scala 76:16:@126235.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@126234.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@126238.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@126232.4]
  assign regs_27_clock = clock; // @[:@126241.4]
  assign regs_27_reset = io_reset; // @[:@126242.4 RegFile.scala 76:16:@126249.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@126248.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@126252.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@126246.4]
  assign regs_28_clock = clock; // @[:@126255.4]
  assign regs_28_reset = io_reset; // @[:@126256.4 RegFile.scala 76:16:@126263.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@126262.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@126266.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@126260.4]
  assign regs_29_clock = clock; // @[:@126269.4]
  assign regs_29_reset = io_reset; // @[:@126270.4 RegFile.scala 76:16:@126277.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@126276.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@126280.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@126274.4]
  assign regs_30_clock = clock; // @[:@126283.4]
  assign regs_30_reset = io_reset; // @[:@126284.4 RegFile.scala 76:16:@126291.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@126290.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@126294.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@126288.4]
  assign regs_31_clock = clock; // @[:@126297.4]
  assign regs_31_reset = io_reset; // @[:@126298.4 RegFile.scala 76:16:@126305.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@126304.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@126308.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@126302.4]
  assign regs_32_clock = clock; // @[:@126311.4]
  assign regs_32_reset = io_reset; // @[:@126312.4 RegFile.scala 76:16:@126319.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@126318.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@126322.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@126316.4]
  assign regs_33_clock = clock; // @[:@126325.4]
  assign regs_33_reset = io_reset; // @[:@126326.4 RegFile.scala 76:16:@126333.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@126332.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@126336.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@126330.4]
  assign regs_34_clock = clock; // @[:@126339.4]
  assign regs_34_reset = io_reset; // @[:@126340.4 RegFile.scala 76:16:@126347.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@126346.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@126350.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@126344.4]
  assign regs_35_clock = clock; // @[:@126353.4]
  assign regs_35_reset = io_reset; // @[:@126354.4 RegFile.scala 76:16:@126361.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@126360.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@126364.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@126358.4]
  assign regs_36_clock = clock; // @[:@126367.4]
  assign regs_36_reset = io_reset; // @[:@126368.4 RegFile.scala 76:16:@126375.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@126374.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@126378.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@126372.4]
  assign regs_37_clock = clock; // @[:@126381.4]
  assign regs_37_reset = io_reset; // @[:@126382.4 RegFile.scala 76:16:@126389.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@126388.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@126392.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@126386.4]
  assign regs_38_clock = clock; // @[:@126395.4]
  assign regs_38_reset = io_reset; // @[:@126396.4 RegFile.scala 76:16:@126403.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@126402.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@126406.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@126400.4]
  assign regs_39_clock = clock; // @[:@126409.4]
  assign regs_39_reset = io_reset; // @[:@126410.4 RegFile.scala 76:16:@126417.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@126416.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@126420.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@126414.4]
  assign regs_40_clock = clock; // @[:@126423.4]
  assign regs_40_reset = io_reset; // @[:@126424.4 RegFile.scala 76:16:@126431.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@126430.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@126434.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@126428.4]
  assign regs_41_clock = clock; // @[:@126437.4]
  assign regs_41_reset = io_reset; // @[:@126438.4 RegFile.scala 76:16:@126445.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@126444.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@126448.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@126442.4]
  assign regs_42_clock = clock; // @[:@126451.4]
  assign regs_42_reset = io_reset; // @[:@126452.4 RegFile.scala 76:16:@126459.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@126458.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@126462.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@126456.4]
  assign regs_43_clock = clock; // @[:@126465.4]
  assign regs_43_reset = io_reset; // @[:@126466.4 RegFile.scala 76:16:@126473.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@126472.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@126476.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@126470.4]
  assign regs_44_clock = clock; // @[:@126479.4]
  assign regs_44_reset = io_reset; // @[:@126480.4 RegFile.scala 76:16:@126487.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@126486.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@126490.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@126484.4]
  assign regs_45_clock = clock; // @[:@126493.4]
  assign regs_45_reset = io_reset; // @[:@126494.4 RegFile.scala 76:16:@126501.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@126500.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@126504.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@126498.4]
  assign regs_46_clock = clock; // @[:@126507.4]
  assign regs_46_reset = io_reset; // @[:@126508.4 RegFile.scala 76:16:@126515.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@126514.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@126518.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@126512.4]
  assign regs_47_clock = clock; // @[:@126521.4]
  assign regs_47_reset = io_reset; // @[:@126522.4 RegFile.scala 76:16:@126529.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@126528.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@126532.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@126526.4]
  assign regs_48_clock = clock; // @[:@126535.4]
  assign regs_48_reset = io_reset; // @[:@126536.4 RegFile.scala 76:16:@126543.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@126542.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@126546.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@126540.4]
  assign regs_49_clock = clock; // @[:@126549.4]
  assign regs_49_reset = io_reset; // @[:@126550.4 RegFile.scala 76:16:@126557.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@126556.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@126560.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@126554.4]
  assign regs_50_clock = clock; // @[:@126563.4]
  assign regs_50_reset = io_reset; // @[:@126564.4 RegFile.scala 76:16:@126571.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@126570.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@126574.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@126568.4]
  assign regs_51_clock = clock; // @[:@126577.4]
  assign regs_51_reset = io_reset; // @[:@126578.4 RegFile.scala 76:16:@126585.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@126584.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@126588.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@126582.4]
  assign regs_52_clock = clock; // @[:@126591.4]
  assign regs_52_reset = io_reset; // @[:@126592.4 RegFile.scala 76:16:@126599.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@126598.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@126602.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@126596.4]
  assign regs_53_clock = clock; // @[:@126605.4]
  assign regs_53_reset = io_reset; // @[:@126606.4 RegFile.scala 76:16:@126613.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@126612.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@126616.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@126610.4]
  assign regs_54_clock = clock; // @[:@126619.4]
  assign regs_54_reset = io_reset; // @[:@126620.4 RegFile.scala 76:16:@126627.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@126626.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@126630.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@126624.4]
  assign regs_55_clock = clock; // @[:@126633.4]
  assign regs_55_reset = io_reset; // @[:@126634.4 RegFile.scala 76:16:@126641.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@126640.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@126644.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@126638.4]
  assign regs_56_clock = clock; // @[:@126647.4]
  assign regs_56_reset = io_reset; // @[:@126648.4 RegFile.scala 76:16:@126655.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@126654.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@126658.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@126652.4]
  assign regs_57_clock = clock; // @[:@126661.4]
  assign regs_57_reset = io_reset; // @[:@126662.4 RegFile.scala 76:16:@126669.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@126668.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@126672.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@126666.4]
  assign regs_58_clock = clock; // @[:@126675.4]
  assign regs_58_reset = io_reset; // @[:@126676.4 RegFile.scala 76:16:@126683.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@126682.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@126686.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@126680.4]
  assign regs_59_clock = clock; // @[:@126689.4]
  assign regs_59_reset = io_reset; // @[:@126690.4 RegFile.scala 76:16:@126697.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@126696.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@126700.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@126694.4]
  assign regs_60_clock = clock; // @[:@126703.4]
  assign regs_60_reset = io_reset; // @[:@126704.4 RegFile.scala 76:16:@126711.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@126710.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@126714.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@126708.4]
  assign regs_61_clock = clock; // @[:@126717.4]
  assign regs_61_reset = io_reset; // @[:@126718.4 RegFile.scala 76:16:@126725.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@126724.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@126728.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@126722.4]
  assign regs_62_clock = clock; // @[:@126731.4]
  assign regs_62_reset = io_reset; // @[:@126732.4 RegFile.scala 76:16:@126739.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@126738.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@126742.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@126736.4]
  assign regs_63_clock = clock; // @[:@126745.4]
  assign regs_63_reset = io_reset; // @[:@126746.4 RegFile.scala 76:16:@126753.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@126752.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@126756.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@126750.4]
  assign regs_64_clock = clock; // @[:@126759.4]
  assign regs_64_reset = io_reset; // @[:@126760.4 RegFile.scala 76:16:@126767.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@126766.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@126770.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@126764.4]
  assign regs_65_clock = clock; // @[:@126773.4]
  assign regs_65_reset = io_reset; // @[:@126774.4 RegFile.scala 76:16:@126781.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@126780.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@126784.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@126778.4]
  assign regs_66_clock = clock; // @[:@126787.4]
  assign regs_66_reset = io_reset; // @[:@126788.4 RegFile.scala 76:16:@126795.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@126794.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@126798.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@126792.4]
  assign regs_67_clock = clock; // @[:@126801.4]
  assign regs_67_reset = io_reset; // @[:@126802.4 RegFile.scala 76:16:@126809.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@126808.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@126812.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@126806.4]
  assign regs_68_clock = clock; // @[:@126815.4]
  assign regs_68_reset = io_reset; // @[:@126816.4 RegFile.scala 76:16:@126823.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@126822.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@126826.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@126820.4]
  assign regs_69_clock = clock; // @[:@126829.4]
  assign regs_69_reset = io_reset; // @[:@126830.4 RegFile.scala 76:16:@126837.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@126836.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@126840.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@126834.4]
  assign regs_70_clock = clock; // @[:@126843.4]
  assign regs_70_reset = io_reset; // @[:@126844.4 RegFile.scala 76:16:@126851.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@126850.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@126854.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@126848.4]
  assign regs_71_clock = clock; // @[:@126857.4]
  assign regs_71_reset = io_reset; // @[:@126858.4 RegFile.scala 76:16:@126865.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@126864.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@126868.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@126862.4]
  assign regs_72_clock = clock; // @[:@126871.4]
  assign regs_72_reset = io_reset; // @[:@126872.4 RegFile.scala 76:16:@126879.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@126878.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@126882.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@126876.4]
  assign regs_73_clock = clock; // @[:@126885.4]
  assign regs_73_reset = io_reset; // @[:@126886.4 RegFile.scala 76:16:@126893.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@126892.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@126896.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@126890.4]
  assign regs_74_clock = clock; // @[:@126899.4]
  assign regs_74_reset = io_reset; // @[:@126900.4 RegFile.scala 76:16:@126907.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@126906.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@126910.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@126904.4]
  assign regs_75_clock = clock; // @[:@126913.4]
  assign regs_75_reset = io_reset; // @[:@126914.4 RegFile.scala 76:16:@126921.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@126920.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@126924.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@126918.4]
  assign regs_76_clock = clock; // @[:@126927.4]
  assign regs_76_reset = io_reset; // @[:@126928.4 RegFile.scala 76:16:@126935.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@126934.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@126938.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@126932.4]
  assign regs_77_clock = clock; // @[:@126941.4]
  assign regs_77_reset = io_reset; // @[:@126942.4 RegFile.scala 76:16:@126949.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@126948.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@126952.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@126946.4]
  assign regs_78_clock = clock; // @[:@126955.4]
  assign regs_78_reset = io_reset; // @[:@126956.4 RegFile.scala 76:16:@126963.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@126962.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@126966.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@126960.4]
  assign regs_79_clock = clock; // @[:@126969.4]
  assign regs_79_reset = io_reset; // @[:@126970.4 RegFile.scala 76:16:@126977.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@126976.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@126980.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@126974.4]
  assign regs_80_clock = clock; // @[:@126983.4]
  assign regs_80_reset = io_reset; // @[:@126984.4 RegFile.scala 76:16:@126991.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@126990.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@126994.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@126988.4]
  assign regs_81_clock = clock; // @[:@126997.4]
  assign regs_81_reset = io_reset; // @[:@126998.4 RegFile.scala 76:16:@127005.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@127004.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@127008.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@127002.4]
  assign regs_82_clock = clock; // @[:@127011.4]
  assign regs_82_reset = io_reset; // @[:@127012.4 RegFile.scala 76:16:@127019.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@127018.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@127022.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@127016.4]
  assign regs_83_clock = clock; // @[:@127025.4]
  assign regs_83_reset = io_reset; // @[:@127026.4 RegFile.scala 76:16:@127033.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@127032.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@127036.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@127030.4]
  assign regs_84_clock = clock; // @[:@127039.4]
  assign regs_84_reset = io_reset; // @[:@127040.4 RegFile.scala 76:16:@127047.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@127046.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@127050.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@127044.4]
  assign regs_85_clock = clock; // @[:@127053.4]
  assign regs_85_reset = io_reset; // @[:@127054.4 RegFile.scala 76:16:@127061.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@127060.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@127064.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@127058.4]
  assign regs_86_clock = clock; // @[:@127067.4]
  assign regs_86_reset = io_reset; // @[:@127068.4 RegFile.scala 76:16:@127075.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@127074.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@127078.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@127072.4]
  assign regs_87_clock = clock; // @[:@127081.4]
  assign regs_87_reset = io_reset; // @[:@127082.4 RegFile.scala 76:16:@127089.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@127088.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@127092.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@127086.4]
  assign regs_88_clock = clock; // @[:@127095.4]
  assign regs_88_reset = io_reset; // @[:@127096.4 RegFile.scala 76:16:@127103.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@127102.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@127106.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@127100.4]
  assign regs_89_clock = clock; // @[:@127109.4]
  assign regs_89_reset = io_reset; // @[:@127110.4 RegFile.scala 76:16:@127117.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@127116.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@127120.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@127114.4]
  assign regs_90_clock = clock; // @[:@127123.4]
  assign regs_90_reset = io_reset; // @[:@127124.4 RegFile.scala 76:16:@127131.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@127130.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@127134.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@127128.4]
  assign regs_91_clock = clock; // @[:@127137.4]
  assign regs_91_reset = io_reset; // @[:@127138.4 RegFile.scala 76:16:@127145.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@127144.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@127148.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@127142.4]
  assign regs_92_clock = clock; // @[:@127151.4]
  assign regs_92_reset = io_reset; // @[:@127152.4 RegFile.scala 76:16:@127159.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@127158.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@127162.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@127156.4]
  assign regs_93_clock = clock; // @[:@127165.4]
  assign regs_93_reset = io_reset; // @[:@127166.4 RegFile.scala 76:16:@127173.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@127172.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@127176.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@127170.4]
  assign regs_94_clock = clock; // @[:@127179.4]
  assign regs_94_reset = io_reset; // @[:@127180.4 RegFile.scala 76:16:@127187.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@127186.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@127190.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@127184.4]
  assign regs_95_clock = clock; // @[:@127193.4]
  assign regs_95_reset = io_reset; // @[:@127194.4 RegFile.scala 76:16:@127201.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@127200.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@127204.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@127198.4]
  assign regs_96_clock = clock; // @[:@127207.4]
  assign regs_96_reset = io_reset; // @[:@127208.4 RegFile.scala 76:16:@127215.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@127214.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@127218.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@127212.4]
  assign regs_97_clock = clock; // @[:@127221.4]
  assign regs_97_reset = io_reset; // @[:@127222.4 RegFile.scala 76:16:@127229.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@127228.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@127232.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@127226.4]
  assign regs_98_clock = clock; // @[:@127235.4]
  assign regs_98_reset = io_reset; // @[:@127236.4 RegFile.scala 76:16:@127243.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@127242.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@127246.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@127240.4]
  assign regs_99_clock = clock; // @[:@127249.4]
  assign regs_99_reset = io_reset; // @[:@127250.4 RegFile.scala 76:16:@127257.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@127256.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@127260.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@127254.4]
  assign regs_100_clock = clock; // @[:@127263.4]
  assign regs_100_reset = io_reset; // @[:@127264.4 RegFile.scala 76:16:@127271.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@127270.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@127274.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@127268.4]
  assign regs_101_clock = clock; // @[:@127277.4]
  assign regs_101_reset = io_reset; // @[:@127278.4 RegFile.scala 76:16:@127285.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@127284.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@127288.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@127282.4]
  assign regs_102_clock = clock; // @[:@127291.4]
  assign regs_102_reset = io_reset; // @[:@127292.4 RegFile.scala 76:16:@127299.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@127298.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@127302.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@127296.4]
  assign regs_103_clock = clock; // @[:@127305.4]
  assign regs_103_reset = io_reset; // @[:@127306.4 RegFile.scala 76:16:@127313.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@127312.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@127316.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@127310.4]
  assign regs_104_clock = clock; // @[:@127319.4]
  assign regs_104_reset = io_reset; // @[:@127320.4 RegFile.scala 76:16:@127327.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@127326.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@127330.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@127324.4]
  assign regs_105_clock = clock; // @[:@127333.4]
  assign regs_105_reset = io_reset; // @[:@127334.4 RegFile.scala 76:16:@127341.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@127340.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@127344.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@127338.4]
  assign regs_106_clock = clock; // @[:@127347.4]
  assign regs_106_reset = io_reset; // @[:@127348.4 RegFile.scala 76:16:@127355.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@127354.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@127358.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@127352.4]
  assign regs_107_clock = clock; // @[:@127361.4]
  assign regs_107_reset = io_reset; // @[:@127362.4 RegFile.scala 76:16:@127369.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@127368.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@127372.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@127366.4]
  assign regs_108_clock = clock; // @[:@127375.4]
  assign regs_108_reset = io_reset; // @[:@127376.4 RegFile.scala 76:16:@127383.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@127382.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@127386.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@127380.4]
  assign regs_109_clock = clock; // @[:@127389.4]
  assign regs_109_reset = io_reset; // @[:@127390.4 RegFile.scala 76:16:@127397.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@127396.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@127400.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@127394.4]
  assign regs_110_clock = clock; // @[:@127403.4]
  assign regs_110_reset = io_reset; // @[:@127404.4 RegFile.scala 76:16:@127411.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@127410.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@127414.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@127408.4]
  assign regs_111_clock = clock; // @[:@127417.4]
  assign regs_111_reset = io_reset; // @[:@127418.4 RegFile.scala 76:16:@127425.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@127424.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@127428.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@127422.4]
  assign regs_112_clock = clock; // @[:@127431.4]
  assign regs_112_reset = io_reset; // @[:@127432.4 RegFile.scala 76:16:@127439.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@127438.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@127442.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@127436.4]
  assign regs_113_clock = clock; // @[:@127445.4]
  assign regs_113_reset = io_reset; // @[:@127446.4 RegFile.scala 76:16:@127453.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@127452.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@127456.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@127450.4]
  assign regs_114_clock = clock; // @[:@127459.4]
  assign regs_114_reset = io_reset; // @[:@127460.4 RegFile.scala 76:16:@127467.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@127466.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@127470.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@127464.4]
  assign regs_115_clock = clock; // @[:@127473.4]
  assign regs_115_reset = io_reset; // @[:@127474.4 RegFile.scala 76:16:@127481.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@127480.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@127484.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@127478.4]
  assign regs_116_clock = clock; // @[:@127487.4]
  assign regs_116_reset = io_reset; // @[:@127488.4 RegFile.scala 76:16:@127495.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@127494.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@127498.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@127492.4]
  assign regs_117_clock = clock; // @[:@127501.4]
  assign regs_117_reset = io_reset; // @[:@127502.4 RegFile.scala 76:16:@127509.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@127508.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@127512.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@127506.4]
  assign regs_118_clock = clock; // @[:@127515.4]
  assign regs_118_reset = io_reset; // @[:@127516.4 RegFile.scala 76:16:@127523.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@127522.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@127526.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@127520.4]
  assign regs_119_clock = clock; // @[:@127529.4]
  assign regs_119_reset = io_reset; // @[:@127530.4 RegFile.scala 76:16:@127537.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@127536.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@127540.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@127534.4]
  assign regs_120_clock = clock; // @[:@127543.4]
  assign regs_120_reset = io_reset; // @[:@127544.4 RegFile.scala 76:16:@127551.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@127550.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@127554.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@127548.4]
  assign regs_121_clock = clock; // @[:@127557.4]
  assign regs_121_reset = io_reset; // @[:@127558.4 RegFile.scala 76:16:@127565.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@127564.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@127568.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@127562.4]
  assign regs_122_clock = clock; // @[:@127571.4]
  assign regs_122_reset = io_reset; // @[:@127572.4 RegFile.scala 76:16:@127579.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@127578.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@127582.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@127576.4]
  assign regs_123_clock = clock; // @[:@127585.4]
  assign regs_123_reset = io_reset; // @[:@127586.4 RegFile.scala 76:16:@127593.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@127592.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@127596.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@127590.4]
  assign regs_124_clock = clock; // @[:@127599.4]
  assign regs_124_reset = io_reset; // @[:@127600.4 RegFile.scala 76:16:@127607.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@127606.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@127610.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@127604.4]
  assign regs_125_clock = clock; // @[:@127613.4]
  assign regs_125_reset = io_reset; // @[:@127614.4 RegFile.scala 76:16:@127621.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@127620.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@127624.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@127618.4]
  assign regs_126_clock = clock; // @[:@127627.4]
  assign regs_126_reset = io_reset; // @[:@127628.4 RegFile.scala 76:16:@127635.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@127634.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@127638.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@127632.4]
  assign regs_127_clock = clock; // @[:@127641.4]
  assign regs_127_reset = io_reset; // @[:@127642.4 RegFile.scala 76:16:@127649.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@127648.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@127652.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@127646.4]
  assign regs_128_clock = clock; // @[:@127655.4]
  assign regs_128_reset = io_reset; // @[:@127656.4 RegFile.scala 76:16:@127663.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@127662.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@127666.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@127660.4]
  assign regs_129_clock = clock; // @[:@127669.4]
  assign regs_129_reset = io_reset; // @[:@127670.4 RegFile.scala 76:16:@127677.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@127676.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@127680.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@127674.4]
  assign regs_130_clock = clock; // @[:@127683.4]
  assign regs_130_reset = io_reset; // @[:@127684.4 RegFile.scala 76:16:@127691.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@127690.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@127694.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@127688.4]
  assign regs_131_clock = clock; // @[:@127697.4]
  assign regs_131_reset = io_reset; // @[:@127698.4 RegFile.scala 76:16:@127705.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@127704.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@127708.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@127702.4]
  assign regs_132_clock = clock; // @[:@127711.4]
  assign regs_132_reset = io_reset; // @[:@127712.4 RegFile.scala 76:16:@127719.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@127718.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@127722.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@127716.4]
  assign regs_133_clock = clock; // @[:@127725.4]
  assign regs_133_reset = io_reset; // @[:@127726.4 RegFile.scala 76:16:@127733.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@127732.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@127736.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@127730.4]
  assign regs_134_clock = clock; // @[:@127739.4]
  assign regs_134_reset = io_reset; // @[:@127740.4 RegFile.scala 76:16:@127747.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@127746.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@127750.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@127744.4]
  assign regs_135_clock = clock; // @[:@127753.4]
  assign regs_135_reset = io_reset; // @[:@127754.4 RegFile.scala 76:16:@127761.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@127760.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@127764.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@127758.4]
  assign regs_136_clock = clock; // @[:@127767.4]
  assign regs_136_reset = io_reset; // @[:@127768.4 RegFile.scala 76:16:@127775.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@127774.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@127778.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@127772.4]
  assign regs_137_clock = clock; // @[:@127781.4]
  assign regs_137_reset = io_reset; // @[:@127782.4 RegFile.scala 76:16:@127789.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@127788.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@127792.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@127786.4]
  assign regs_138_clock = clock; // @[:@127795.4]
  assign regs_138_reset = io_reset; // @[:@127796.4 RegFile.scala 76:16:@127803.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@127802.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@127806.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@127800.4]
  assign regs_139_clock = clock; // @[:@127809.4]
  assign regs_139_reset = io_reset; // @[:@127810.4 RegFile.scala 76:16:@127817.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@127816.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@127820.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@127814.4]
  assign regs_140_clock = clock; // @[:@127823.4]
  assign regs_140_reset = io_reset; // @[:@127824.4 RegFile.scala 76:16:@127831.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@127830.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@127834.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@127828.4]
  assign regs_141_clock = clock; // @[:@127837.4]
  assign regs_141_reset = io_reset; // @[:@127838.4 RegFile.scala 76:16:@127845.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@127844.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@127848.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@127842.4]
  assign regs_142_clock = clock; // @[:@127851.4]
  assign regs_142_reset = io_reset; // @[:@127852.4 RegFile.scala 76:16:@127859.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@127858.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@127862.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@127856.4]
  assign regs_143_clock = clock; // @[:@127865.4]
  assign regs_143_reset = io_reset; // @[:@127866.4 RegFile.scala 76:16:@127873.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@127872.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@127876.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@127870.4]
  assign regs_144_clock = clock; // @[:@127879.4]
  assign regs_144_reset = io_reset; // @[:@127880.4 RegFile.scala 76:16:@127887.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@127886.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@127890.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@127884.4]
  assign regs_145_clock = clock; // @[:@127893.4]
  assign regs_145_reset = io_reset; // @[:@127894.4 RegFile.scala 76:16:@127901.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@127900.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@127904.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@127898.4]
  assign regs_146_clock = clock; // @[:@127907.4]
  assign regs_146_reset = io_reset; // @[:@127908.4 RegFile.scala 76:16:@127915.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@127914.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@127918.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@127912.4]
  assign regs_147_clock = clock; // @[:@127921.4]
  assign regs_147_reset = io_reset; // @[:@127922.4 RegFile.scala 76:16:@127929.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@127928.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@127932.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@127926.4]
  assign regs_148_clock = clock; // @[:@127935.4]
  assign regs_148_reset = io_reset; // @[:@127936.4 RegFile.scala 76:16:@127943.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@127942.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@127946.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@127940.4]
  assign regs_149_clock = clock; // @[:@127949.4]
  assign regs_149_reset = io_reset; // @[:@127950.4 RegFile.scala 76:16:@127957.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@127956.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@127960.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@127954.4]
  assign regs_150_clock = clock; // @[:@127963.4]
  assign regs_150_reset = io_reset; // @[:@127964.4 RegFile.scala 76:16:@127971.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@127970.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@127974.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@127968.4]
  assign regs_151_clock = clock; // @[:@127977.4]
  assign regs_151_reset = io_reset; // @[:@127978.4 RegFile.scala 76:16:@127985.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@127984.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@127988.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@127982.4]
  assign regs_152_clock = clock; // @[:@127991.4]
  assign regs_152_reset = io_reset; // @[:@127992.4 RegFile.scala 76:16:@127999.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@127998.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@128002.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@127996.4]
  assign regs_153_clock = clock; // @[:@128005.4]
  assign regs_153_reset = io_reset; // @[:@128006.4 RegFile.scala 76:16:@128013.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@128012.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@128016.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@128010.4]
  assign regs_154_clock = clock; // @[:@128019.4]
  assign regs_154_reset = io_reset; // @[:@128020.4 RegFile.scala 76:16:@128027.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@128026.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@128030.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@128024.4]
  assign regs_155_clock = clock; // @[:@128033.4]
  assign regs_155_reset = io_reset; // @[:@128034.4 RegFile.scala 76:16:@128041.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@128040.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@128044.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@128038.4]
  assign regs_156_clock = clock; // @[:@128047.4]
  assign regs_156_reset = io_reset; // @[:@128048.4 RegFile.scala 76:16:@128055.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@128054.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@128058.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@128052.4]
  assign regs_157_clock = clock; // @[:@128061.4]
  assign regs_157_reset = io_reset; // @[:@128062.4 RegFile.scala 76:16:@128069.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@128068.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@128072.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@128066.4]
  assign regs_158_clock = clock; // @[:@128075.4]
  assign regs_158_reset = io_reset; // @[:@128076.4 RegFile.scala 76:16:@128083.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@128082.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@128086.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@128080.4]
  assign regs_159_clock = clock; // @[:@128089.4]
  assign regs_159_reset = io_reset; // @[:@128090.4 RegFile.scala 76:16:@128097.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@128096.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@128100.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@128094.4]
  assign regs_160_clock = clock; // @[:@128103.4]
  assign regs_160_reset = io_reset; // @[:@128104.4 RegFile.scala 76:16:@128111.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@128110.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@128114.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@128108.4]
  assign regs_161_clock = clock; // @[:@128117.4]
  assign regs_161_reset = io_reset; // @[:@128118.4 RegFile.scala 76:16:@128125.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@128124.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@128128.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@128122.4]
  assign regs_162_clock = clock; // @[:@128131.4]
  assign regs_162_reset = io_reset; // @[:@128132.4 RegFile.scala 76:16:@128139.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@128138.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@128142.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@128136.4]
  assign regs_163_clock = clock; // @[:@128145.4]
  assign regs_163_reset = io_reset; // @[:@128146.4 RegFile.scala 76:16:@128153.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@128152.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@128156.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@128150.4]
  assign regs_164_clock = clock; // @[:@128159.4]
  assign regs_164_reset = io_reset; // @[:@128160.4 RegFile.scala 76:16:@128167.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@128166.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@128170.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@128164.4]
  assign regs_165_clock = clock; // @[:@128173.4]
  assign regs_165_reset = io_reset; // @[:@128174.4 RegFile.scala 76:16:@128181.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@128180.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@128184.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@128178.4]
  assign regs_166_clock = clock; // @[:@128187.4]
  assign regs_166_reset = io_reset; // @[:@128188.4 RegFile.scala 76:16:@128195.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@128194.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@128198.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@128192.4]
  assign regs_167_clock = clock; // @[:@128201.4]
  assign regs_167_reset = io_reset; // @[:@128202.4 RegFile.scala 76:16:@128209.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@128208.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@128212.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@128206.4]
  assign regs_168_clock = clock; // @[:@128215.4]
  assign regs_168_reset = io_reset; // @[:@128216.4 RegFile.scala 76:16:@128223.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@128222.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@128226.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@128220.4]
  assign regs_169_clock = clock; // @[:@128229.4]
  assign regs_169_reset = io_reset; // @[:@128230.4 RegFile.scala 76:16:@128237.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@128236.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@128240.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@128234.4]
  assign regs_170_clock = clock; // @[:@128243.4]
  assign regs_170_reset = io_reset; // @[:@128244.4 RegFile.scala 76:16:@128251.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@128250.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@128254.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@128248.4]
  assign regs_171_clock = clock; // @[:@128257.4]
  assign regs_171_reset = io_reset; // @[:@128258.4 RegFile.scala 76:16:@128265.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@128264.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@128268.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@128262.4]
  assign regs_172_clock = clock; // @[:@128271.4]
  assign regs_172_reset = io_reset; // @[:@128272.4 RegFile.scala 76:16:@128279.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@128278.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@128282.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@128276.4]
  assign regs_173_clock = clock; // @[:@128285.4]
  assign regs_173_reset = io_reset; // @[:@128286.4 RegFile.scala 76:16:@128293.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@128292.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@128296.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@128290.4]
  assign regs_174_clock = clock; // @[:@128299.4]
  assign regs_174_reset = io_reset; // @[:@128300.4 RegFile.scala 76:16:@128307.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@128306.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@128310.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@128304.4]
  assign regs_175_clock = clock; // @[:@128313.4]
  assign regs_175_reset = io_reset; // @[:@128314.4 RegFile.scala 76:16:@128321.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@128320.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@128324.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@128318.4]
  assign regs_176_clock = clock; // @[:@128327.4]
  assign regs_176_reset = io_reset; // @[:@128328.4 RegFile.scala 76:16:@128335.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@128334.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@128338.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@128332.4]
  assign regs_177_clock = clock; // @[:@128341.4]
  assign regs_177_reset = io_reset; // @[:@128342.4 RegFile.scala 76:16:@128349.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@128348.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@128352.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@128346.4]
  assign regs_178_clock = clock; // @[:@128355.4]
  assign regs_178_reset = io_reset; // @[:@128356.4 RegFile.scala 76:16:@128363.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@128362.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@128366.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@128360.4]
  assign regs_179_clock = clock; // @[:@128369.4]
  assign regs_179_reset = io_reset; // @[:@128370.4 RegFile.scala 76:16:@128377.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@128376.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@128380.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@128374.4]
  assign regs_180_clock = clock; // @[:@128383.4]
  assign regs_180_reset = io_reset; // @[:@128384.4 RegFile.scala 76:16:@128391.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@128390.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@128394.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@128388.4]
  assign regs_181_clock = clock; // @[:@128397.4]
  assign regs_181_reset = io_reset; // @[:@128398.4 RegFile.scala 76:16:@128405.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@128404.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@128408.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@128402.4]
  assign regs_182_clock = clock; // @[:@128411.4]
  assign regs_182_reset = io_reset; // @[:@128412.4 RegFile.scala 76:16:@128419.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@128418.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@128422.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@128416.4]
  assign regs_183_clock = clock; // @[:@128425.4]
  assign regs_183_reset = io_reset; // @[:@128426.4 RegFile.scala 76:16:@128433.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@128432.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@128436.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@128430.4]
  assign regs_184_clock = clock; // @[:@128439.4]
  assign regs_184_reset = io_reset; // @[:@128440.4 RegFile.scala 76:16:@128447.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@128446.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@128450.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@128444.4]
  assign regs_185_clock = clock; // @[:@128453.4]
  assign regs_185_reset = io_reset; // @[:@128454.4 RegFile.scala 76:16:@128461.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@128460.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@128464.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@128458.4]
  assign regs_186_clock = clock; // @[:@128467.4]
  assign regs_186_reset = io_reset; // @[:@128468.4 RegFile.scala 76:16:@128475.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@128474.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@128478.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@128472.4]
  assign regs_187_clock = clock; // @[:@128481.4]
  assign regs_187_reset = io_reset; // @[:@128482.4 RegFile.scala 76:16:@128489.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@128488.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@128492.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@128486.4]
  assign regs_188_clock = clock; // @[:@128495.4]
  assign regs_188_reset = io_reset; // @[:@128496.4 RegFile.scala 76:16:@128503.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@128502.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@128506.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@128500.4]
  assign regs_189_clock = clock; // @[:@128509.4]
  assign regs_189_reset = io_reset; // @[:@128510.4 RegFile.scala 76:16:@128517.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@128516.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@128520.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@128514.4]
  assign regs_190_clock = clock; // @[:@128523.4]
  assign regs_190_reset = io_reset; // @[:@128524.4 RegFile.scala 76:16:@128531.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@128530.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@128534.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@128528.4]
  assign regs_191_clock = clock; // @[:@128537.4]
  assign regs_191_reset = io_reset; // @[:@128538.4 RegFile.scala 76:16:@128545.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@128544.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@128548.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@128542.4]
  assign regs_192_clock = clock; // @[:@128551.4]
  assign regs_192_reset = io_reset; // @[:@128552.4 RegFile.scala 76:16:@128559.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@128558.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@128562.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@128556.4]
  assign regs_193_clock = clock; // @[:@128565.4]
  assign regs_193_reset = io_reset; // @[:@128566.4 RegFile.scala 76:16:@128573.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@128572.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@128576.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@128570.4]
  assign regs_194_clock = clock; // @[:@128579.4]
  assign regs_194_reset = io_reset; // @[:@128580.4 RegFile.scala 76:16:@128587.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@128586.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@128590.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@128584.4]
  assign regs_195_clock = clock; // @[:@128593.4]
  assign regs_195_reset = io_reset; // @[:@128594.4 RegFile.scala 76:16:@128601.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@128600.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@128604.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@128598.4]
  assign regs_196_clock = clock; // @[:@128607.4]
  assign regs_196_reset = io_reset; // @[:@128608.4 RegFile.scala 76:16:@128615.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@128614.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@128618.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@128612.4]
  assign regs_197_clock = clock; // @[:@128621.4]
  assign regs_197_reset = io_reset; // @[:@128622.4 RegFile.scala 76:16:@128629.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@128628.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@128632.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@128626.4]
  assign regs_198_clock = clock; // @[:@128635.4]
  assign regs_198_reset = io_reset; // @[:@128636.4 RegFile.scala 76:16:@128643.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@128642.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@128646.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@128640.4]
  assign regs_199_clock = clock; // @[:@128649.4]
  assign regs_199_reset = io_reset; // @[:@128650.4 RegFile.scala 76:16:@128657.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@128656.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@128660.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@128654.4]
  assign regs_200_clock = clock; // @[:@128663.4]
  assign regs_200_reset = io_reset; // @[:@128664.4 RegFile.scala 76:16:@128671.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@128670.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@128674.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@128668.4]
  assign regs_201_clock = clock; // @[:@128677.4]
  assign regs_201_reset = io_reset; // @[:@128678.4 RegFile.scala 76:16:@128685.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@128684.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@128688.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@128682.4]
  assign regs_202_clock = clock; // @[:@128691.4]
  assign regs_202_reset = io_reset; // @[:@128692.4 RegFile.scala 76:16:@128699.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@128698.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@128702.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@128696.4]
  assign regs_203_clock = clock; // @[:@128705.4]
  assign regs_203_reset = io_reset; // @[:@128706.4 RegFile.scala 76:16:@128713.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@128712.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@128716.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@128710.4]
  assign regs_204_clock = clock; // @[:@128719.4]
  assign regs_204_reset = io_reset; // @[:@128720.4 RegFile.scala 76:16:@128727.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@128726.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@128730.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@128724.4]
  assign regs_205_clock = clock; // @[:@128733.4]
  assign regs_205_reset = io_reset; // @[:@128734.4 RegFile.scala 76:16:@128741.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@128740.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@128744.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@128738.4]
  assign regs_206_clock = clock; // @[:@128747.4]
  assign regs_206_reset = io_reset; // @[:@128748.4 RegFile.scala 76:16:@128755.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@128754.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@128758.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@128752.4]
  assign regs_207_clock = clock; // @[:@128761.4]
  assign regs_207_reset = io_reset; // @[:@128762.4 RegFile.scala 76:16:@128769.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@128768.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@128772.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@128766.4]
  assign regs_208_clock = clock; // @[:@128775.4]
  assign regs_208_reset = io_reset; // @[:@128776.4 RegFile.scala 76:16:@128783.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@128782.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@128786.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@128780.4]
  assign regs_209_clock = clock; // @[:@128789.4]
  assign regs_209_reset = io_reset; // @[:@128790.4 RegFile.scala 76:16:@128797.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@128796.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@128800.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@128794.4]
  assign regs_210_clock = clock; // @[:@128803.4]
  assign regs_210_reset = io_reset; // @[:@128804.4 RegFile.scala 76:16:@128811.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@128810.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@128814.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@128808.4]
  assign regs_211_clock = clock; // @[:@128817.4]
  assign regs_211_reset = io_reset; // @[:@128818.4 RegFile.scala 76:16:@128825.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@128824.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@128828.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@128822.4]
  assign regs_212_clock = clock; // @[:@128831.4]
  assign regs_212_reset = io_reset; // @[:@128832.4 RegFile.scala 76:16:@128839.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@128838.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@128842.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@128836.4]
  assign regs_213_clock = clock; // @[:@128845.4]
  assign regs_213_reset = io_reset; // @[:@128846.4 RegFile.scala 76:16:@128853.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@128852.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@128856.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@128850.4]
  assign regs_214_clock = clock; // @[:@128859.4]
  assign regs_214_reset = io_reset; // @[:@128860.4 RegFile.scala 76:16:@128867.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@128866.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@128870.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@128864.4]
  assign regs_215_clock = clock; // @[:@128873.4]
  assign regs_215_reset = io_reset; // @[:@128874.4 RegFile.scala 76:16:@128881.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@128880.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@128884.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@128878.4]
  assign regs_216_clock = clock; // @[:@128887.4]
  assign regs_216_reset = io_reset; // @[:@128888.4 RegFile.scala 76:16:@128895.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@128894.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@128898.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@128892.4]
  assign regs_217_clock = clock; // @[:@128901.4]
  assign regs_217_reset = io_reset; // @[:@128902.4 RegFile.scala 76:16:@128909.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@128908.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@128912.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@128906.4]
  assign regs_218_clock = clock; // @[:@128915.4]
  assign regs_218_reset = io_reset; // @[:@128916.4 RegFile.scala 76:16:@128923.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@128922.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@128926.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@128920.4]
  assign regs_219_clock = clock; // @[:@128929.4]
  assign regs_219_reset = io_reset; // @[:@128930.4 RegFile.scala 76:16:@128937.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@128936.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@128940.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@128934.4]
  assign regs_220_clock = clock; // @[:@128943.4]
  assign regs_220_reset = io_reset; // @[:@128944.4 RegFile.scala 76:16:@128951.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@128950.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@128954.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@128948.4]
  assign regs_221_clock = clock; // @[:@128957.4]
  assign regs_221_reset = io_reset; // @[:@128958.4 RegFile.scala 76:16:@128965.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@128964.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@128968.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@128962.4]
  assign regs_222_clock = clock; // @[:@128971.4]
  assign regs_222_reset = io_reset; // @[:@128972.4 RegFile.scala 76:16:@128979.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@128978.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@128982.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@128976.4]
  assign regs_223_clock = clock; // @[:@128985.4]
  assign regs_223_reset = io_reset; // @[:@128986.4 RegFile.scala 76:16:@128993.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@128992.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@128996.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@128990.4]
  assign regs_224_clock = clock; // @[:@128999.4]
  assign regs_224_reset = io_reset; // @[:@129000.4 RegFile.scala 76:16:@129007.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@129006.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@129010.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@129004.4]
  assign regs_225_clock = clock; // @[:@129013.4]
  assign regs_225_reset = io_reset; // @[:@129014.4 RegFile.scala 76:16:@129021.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@129020.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@129024.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@129018.4]
  assign regs_226_clock = clock; // @[:@129027.4]
  assign regs_226_reset = io_reset; // @[:@129028.4 RegFile.scala 76:16:@129035.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@129034.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@129038.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@129032.4]
  assign regs_227_clock = clock; // @[:@129041.4]
  assign regs_227_reset = io_reset; // @[:@129042.4 RegFile.scala 76:16:@129049.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@129048.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@129052.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@129046.4]
  assign regs_228_clock = clock; // @[:@129055.4]
  assign regs_228_reset = io_reset; // @[:@129056.4 RegFile.scala 76:16:@129063.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@129062.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@129066.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@129060.4]
  assign regs_229_clock = clock; // @[:@129069.4]
  assign regs_229_reset = io_reset; // @[:@129070.4 RegFile.scala 76:16:@129077.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@129076.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@129080.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@129074.4]
  assign regs_230_clock = clock; // @[:@129083.4]
  assign regs_230_reset = io_reset; // @[:@129084.4 RegFile.scala 76:16:@129091.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@129090.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@129094.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@129088.4]
  assign regs_231_clock = clock; // @[:@129097.4]
  assign regs_231_reset = io_reset; // @[:@129098.4 RegFile.scala 76:16:@129105.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@129104.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@129108.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@129102.4]
  assign regs_232_clock = clock; // @[:@129111.4]
  assign regs_232_reset = io_reset; // @[:@129112.4 RegFile.scala 76:16:@129119.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@129118.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@129122.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@129116.4]
  assign regs_233_clock = clock; // @[:@129125.4]
  assign regs_233_reset = io_reset; // @[:@129126.4 RegFile.scala 76:16:@129133.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@129132.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@129136.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@129130.4]
  assign regs_234_clock = clock; // @[:@129139.4]
  assign regs_234_reset = io_reset; // @[:@129140.4 RegFile.scala 76:16:@129147.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@129146.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@129150.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@129144.4]
  assign regs_235_clock = clock; // @[:@129153.4]
  assign regs_235_reset = io_reset; // @[:@129154.4 RegFile.scala 76:16:@129161.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@129160.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@129164.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@129158.4]
  assign regs_236_clock = clock; // @[:@129167.4]
  assign regs_236_reset = io_reset; // @[:@129168.4 RegFile.scala 76:16:@129175.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@129174.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@129178.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@129172.4]
  assign regs_237_clock = clock; // @[:@129181.4]
  assign regs_237_reset = io_reset; // @[:@129182.4 RegFile.scala 76:16:@129189.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@129188.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@129192.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@129186.4]
  assign regs_238_clock = clock; // @[:@129195.4]
  assign regs_238_reset = io_reset; // @[:@129196.4 RegFile.scala 76:16:@129203.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@129202.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@129206.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@129200.4]
  assign regs_239_clock = clock; // @[:@129209.4]
  assign regs_239_reset = io_reset; // @[:@129210.4 RegFile.scala 76:16:@129217.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@129216.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@129220.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@129214.4]
  assign regs_240_clock = clock; // @[:@129223.4]
  assign regs_240_reset = io_reset; // @[:@129224.4 RegFile.scala 76:16:@129231.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@129230.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@129234.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@129228.4]
  assign regs_241_clock = clock; // @[:@129237.4]
  assign regs_241_reset = io_reset; // @[:@129238.4 RegFile.scala 76:16:@129245.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@129244.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@129248.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@129242.4]
  assign regs_242_clock = clock; // @[:@129251.4]
  assign regs_242_reset = io_reset; // @[:@129252.4 RegFile.scala 76:16:@129259.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@129258.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@129262.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@129256.4]
  assign regs_243_clock = clock; // @[:@129265.4]
  assign regs_243_reset = io_reset; // @[:@129266.4 RegFile.scala 76:16:@129273.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@129272.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@129276.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@129270.4]
  assign regs_244_clock = clock; // @[:@129279.4]
  assign regs_244_reset = io_reset; // @[:@129280.4 RegFile.scala 76:16:@129287.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@129286.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@129290.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@129284.4]
  assign regs_245_clock = clock; // @[:@129293.4]
  assign regs_245_reset = io_reset; // @[:@129294.4 RegFile.scala 76:16:@129301.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@129300.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@129304.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@129298.4]
  assign regs_246_clock = clock; // @[:@129307.4]
  assign regs_246_reset = io_reset; // @[:@129308.4 RegFile.scala 76:16:@129315.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@129314.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@129318.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@129312.4]
  assign regs_247_clock = clock; // @[:@129321.4]
  assign regs_247_reset = io_reset; // @[:@129322.4 RegFile.scala 76:16:@129329.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@129328.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@129332.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@129326.4]
  assign regs_248_clock = clock; // @[:@129335.4]
  assign regs_248_reset = io_reset; // @[:@129336.4 RegFile.scala 76:16:@129343.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@129342.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@129346.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@129340.4]
  assign regs_249_clock = clock; // @[:@129349.4]
  assign regs_249_reset = io_reset; // @[:@129350.4 RegFile.scala 76:16:@129357.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@129356.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@129360.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@129354.4]
  assign regs_250_clock = clock; // @[:@129363.4]
  assign regs_250_reset = io_reset; // @[:@129364.4 RegFile.scala 76:16:@129371.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@129370.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@129374.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@129368.4]
  assign regs_251_clock = clock; // @[:@129377.4]
  assign regs_251_reset = io_reset; // @[:@129378.4 RegFile.scala 76:16:@129385.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@129384.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@129388.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@129382.4]
  assign regs_252_clock = clock; // @[:@129391.4]
  assign regs_252_reset = io_reset; // @[:@129392.4 RegFile.scala 76:16:@129399.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@129398.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@129402.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@129396.4]
  assign regs_253_clock = clock; // @[:@129405.4]
  assign regs_253_reset = io_reset; // @[:@129406.4 RegFile.scala 76:16:@129413.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@129412.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@129416.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@129410.4]
  assign regs_254_clock = clock; // @[:@129419.4]
  assign regs_254_reset = io_reset; // @[:@129420.4 RegFile.scala 76:16:@129427.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@129426.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@129430.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@129424.4]
  assign regs_255_clock = clock; // @[:@129433.4]
  assign regs_255_reset = io_reset; // @[:@129434.4 RegFile.scala 76:16:@129441.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@129440.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@129444.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@129438.4]
  assign regs_256_clock = clock; // @[:@129447.4]
  assign regs_256_reset = io_reset; // @[:@129448.4 RegFile.scala 76:16:@129455.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@129454.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@129458.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@129452.4]
  assign regs_257_clock = clock; // @[:@129461.4]
  assign regs_257_reset = io_reset; // @[:@129462.4 RegFile.scala 76:16:@129469.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@129468.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@129472.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@129466.4]
  assign regs_258_clock = clock; // @[:@129475.4]
  assign regs_258_reset = io_reset; // @[:@129476.4 RegFile.scala 76:16:@129483.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@129482.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@129486.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@129480.4]
  assign regs_259_clock = clock; // @[:@129489.4]
  assign regs_259_reset = io_reset; // @[:@129490.4 RegFile.scala 76:16:@129497.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@129496.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@129500.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@129494.4]
  assign regs_260_clock = clock; // @[:@129503.4]
  assign regs_260_reset = io_reset; // @[:@129504.4 RegFile.scala 76:16:@129511.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@129510.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@129514.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@129508.4]
  assign regs_261_clock = clock; // @[:@129517.4]
  assign regs_261_reset = io_reset; // @[:@129518.4 RegFile.scala 76:16:@129525.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@129524.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@129528.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@129522.4]
  assign regs_262_clock = clock; // @[:@129531.4]
  assign regs_262_reset = io_reset; // @[:@129532.4 RegFile.scala 76:16:@129539.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@129538.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@129542.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@129536.4]
  assign regs_263_clock = clock; // @[:@129545.4]
  assign regs_263_reset = io_reset; // @[:@129546.4 RegFile.scala 76:16:@129553.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@129552.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@129556.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@129550.4]
  assign regs_264_clock = clock; // @[:@129559.4]
  assign regs_264_reset = io_reset; // @[:@129560.4 RegFile.scala 76:16:@129567.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@129566.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@129570.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@129564.4]
  assign regs_265_clock = clock; // @[:@129573.4]
  assign regs_265_reset = io_reset; // @[:@129574.4 RegFile.scala 76:16:@129581.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@129580.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@129584.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@129578.4]
  assign regs_266_clock = clock; // @[:@129587.4]
  assign regs_266_reset = io_reset; // @[:@129588.4 RegFile.scala 76:16:@129595.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@129594.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@129598.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@129592.4]
  assign regs_267_clock = clock; // @[:@129601.4]
  assign regs_267_reset = io_reset; // @[:@129602.4 RegFile.scala 76:16:@129609.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@129608.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@129612.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@129606.4]
  assign regs_268_clock = clock; // @[:@129615.4]
  assign regs_268_reset = io_reset; // @[:@129616.4 RegFile.scala 76:16:@129623.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@129622.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@129626.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@129620.4]
  assign regs_269_clock = clock; // @[:@129629.4]
  assign regs_269_reset = io_reset; // @[:@129630.4 RegFile.scala 76:16:@129637.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@129636.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@129640.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@129634.4]
  assign regs_270_clock = clock; // @[:@129643.4]
  assign regs_270_reset = io_reset; // @[:@129644.4 RegFile.scala 76:16:@129651.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@129650.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@129654.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@129648.4]
  assign regs_271_clock = clock; // @[:@129657.4]
  assign regs_271_reset = io_reset; // @[:@129658.4 RegFile.scala 76:16:@129665.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@129664.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@129668.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@129662.4]
  assign regs_272_clock = clock; // @[:@129671.4]
  assign regs_272_reset = io_reset; // @[:@129672.4 RegFile.scala 76:16:@129679.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@129678.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@129682.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@129676.4]
  assign regs_273_clock = clock; // @[:@129685.4]
  assign regs_273_reset = io_reset; // @[:@129686.4 RegFile.scala 76:16:@129693.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@129692.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@129696.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@129690.4]
  assign regs_274_clock = clock; // @[:@129699.4]
  assign regs_274_reset = io_reset; // @[:@129700.4 RegFile.scala 76:16:@129707.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@129706.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@129710.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@129704.4]
  assign regs_275_clock = clock; // @[:@129713.4]
  assign regs_275_reset = io_reset; // @[:@129714.4 RegFile.scala 76:16:@129721.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@129720.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@129724.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@129718.4]
  assign regs_276_clock = clock; // @[:@129727.4]
  assign regs_276_reset = io_reset; // @[:@129728.4 RegFile.scala 76:16:@129735.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@129734.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@129738.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@129732.4]
  assign regs_277_clock = clock; // @[:@129741.4]
  assign regs_277_reset = io_reset; // @[:@129742.4 RegFile.scala 76:16:@129749.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@129748.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@129752.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@129746.4]
  assign regs_278_clock = clock; // @[:@129755.4]
  assign regs_278_reset = io_reset; // @[:@129756.4 RegFile.scala 76:16:@129763.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@129762.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@129766.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@129760.4]
  assign regs_279_clock = clock; // @[:@129769.4]
  assign regs_279_reset = io_reset; // @[:@129770.4 RegFile.scala 76:16:@129777.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@129776.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@129780.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@129774.4]
  assign regs_280_clock = clock; // @[:@129783.4]
  assign regs_280_reset = io_reset; // @[:@129784.4 RegFile.scala 76:16:@129791.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@129790.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@129794.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@129788.4]
  assign regs_281_clock = clock; // @[:@129797.4]
  assign regs_281_reset = io_reset; // @[:@129798.4 RegFile.scala 76:16:@129805.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@129804.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@129808.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@129802.4]
  assign regs_282_clock = clock; // @[:@129811.4]
  assign regs_282_reset = io_reset; // @[:@129812.4 RegFile.scala 76:16:@129819.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@129818.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@129822.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@129816.4]
  assign regs_283_clock = clock; // @[:@129825.4]
  assign regs_283_reset = io_reset; // @[:@129826.4 RegFile.scala 76:16:@129833.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@129832.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@129836.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@129830.4]
  assign regs_284_clock = clock; // @[:@129839.4]
  assign regs_284_reset = io_reset; // @[:@129840.4 RegFile.scala 76:16:@129847.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@129846.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@129850.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@129844.4]
  assign regs_285_clock = clock; // @[:@129853.4]
  assign regs_285_reset = io_reset; // @[:@129854.4 RegFile.scala 76:16:@129861.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@129860.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@129864.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@129858.4]
  assign regs_286_clock = clock; // @[:@129867.4]
  assign regs_286_reset = io_reset; // @[:@129868.4 RegFile.scala 76:16:@129875.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@129874.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@129878.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@129872.4]
  assign regs_287_clock = clock; // @[:@129881.4]
  assign regs_287_reset = io_reset; // @[:@129882.4 RegFile.scala 76:16:@129889.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@129888.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@129892.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@129886.4]
  assign regs_288_clock = clock; // @[:@129895.4]
  assign regs_288_reset = io_reset; // @[:@129896.4 RegFile.scala 76:16:@129903.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@129902.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@129906.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@129900.4]
  assign regs_289_clock = clock; // @[:@129909.4]
  assign regs_289_reset = io_reset; // @[:@129910.4 RegFile.scala 76:16:@129917.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@129916.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@129920.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@129914.4]
  assign regs_290_clock = clock; // @[:@129923.4]
  assign regs_290_reset = io_reset; // @[:@129924.4 RegFile.scala 76:16:@129931.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@129930.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@129934.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@129928.4]
  assign regs_291_clock = clock; // @[:@129937.4]
  assign regs_291_reset = io_reset; // @[:@129938.4 RegFile.scala 76:16:@129945.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@129944.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@129948.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@129942.4]
  assign regs_292_clock = clock; // @[:@129951.4]
  assign regs_292_reset = io_reset; // @[:@129952.4 RegFile.scala 76:16:@129959.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@129958.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@129962.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@129956.4]
  assign regs_293_clock = clock; // @[:@129965.4]
  assign regs_293_reset = io_reset; // @[:@129966.4 RegFile.scala 76:16:@129973.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@129972.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@129976.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@129970.4]
  assign regs_294_clock = clock; // @[:@129979.4]
  assign regs_294_reset = io_reset; // @[:@129980.4 RegFile.scala 76:16:@129987.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@129986.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@129990.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@129984.4]
  assign regs_295_clock = clock; // @[:@129993.4]
  assign regs_295_reset = io_reset; // @[:@129994.4 RegFile.scala 76:16:@130001.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@130000.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@130004.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@129998.4]
  assign regs_296_clock = clock; // @[:@130007.4]
  assign regs_296_reset = io_reset; // @[:@130008.4 RegFile.scala 76:16:@130015.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@130014.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@130018.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@130012.4]
  assign regs_297_clock = clock; // @[:@130021.4]
  assign regs_297_reset = io_reset; // @[:@130022.4 RegFile.scala 76:16:@130029.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@130028.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@130032.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@130026.4]
  assign regs_298_clock = clock; // @[:@130035.4]
  assign regs_298_reset = io_reset; // @[:@130036.4 RegFile.scala 76:16:@130043.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@130042.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@130046.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@130040.4]
  assign regs_299_clock = clock; // @[:@130049.4]
  assign regs_299_reset = io_reset; // @[:@130050.4 RegFile.scala 76:16:@130057.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@130056.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@130060.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@130054.4]
  assign regs_300_clock = clock; // @[:@130063.4]
  assign regs_300_reset = io_reset; // @[:@130064.4 RegFile.scala 76:16:@130071.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@130070.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@130074.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@130068.4]
  assign regs_301_clock = clock; // @[:@130077.4]
  assign regs_301_reset = io_reset; // @[:@130078.4 RegFile.scala 76:16:@130085.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@130084.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@130088.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@130082.4]
  assign regs_302_clock = clock; // @[:@130091.4]
  assign regs_302_reset = io_reset; // @[:@130092.4 RegFile.scala 76:16:@130099.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@130098.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@130102.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@130096.4]
  assign regs_303_clock = clock; // @[:@130105.4]
  assign regs_303_reset = io_reset; // @[:@130106.4 RegFile.scala 76:16:@130113.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@130112.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@130116.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@130110.4]
  assign regs_304_clock = clock; // @[:@130119.4]
  assign regs_304_reset = io_reset; // @[:@130120.4 RegFile.scala 76:16:@130127.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@130126.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@130130.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@130124.4]
  assign regs_305_clock = clock; // @[:@130133.4]
  assign regs_305_reset = io_reset; // @[:@130134.4 RegFile.scala 76:16:@130141.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@130140.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@130144.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@130138.4]
  assign regs_306_clock = clock; // @[:@130147.4]
  assign regs_306_reset = io_reset; // @[:@130148.4 RegFile.scala 76:16:@130155.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@130154.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@130158.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@130152.4]
  assign regs_307_clock = clock; // @[:@130161.4]
  assign regs_307_reset = io_reset; // @[:@130162.4 RegFile.scala 76:16:@130169.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@130168.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@130172.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@130166.4]
  assign regs_308_clock = clock; // @[:@130175.4]
  assign regs_308_reset = io_reset; // @[:@130176.4 RegFile.scala 76:16:@130183.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@130182.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@130186.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@130180.4]
  assign regs_309_clock = clock; // @[:@130189.4]
  assign regs_309_reset = io_reset; // @[:@130190.4 RegFile.scala 76:16:@130197.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@130196.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@130200.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@130194.4]
  assign regs_310_clock = clock; // @[:@130203.4]
  assign regs_310_reset = io_reset; // @[:@130204.4 RegFile.scala 76:16:@130211.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@130210.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@130214.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@130208.4]
  assign regs_311_clock = clock; // @[:@130217.4]
  assign regs_311_reset = io_reset; // @[:@130218.4 RegFile.scala 76:16:@130225.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@130224.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@130228.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@130222.4]
  assign regs_312_clock = clock; // @[:@130231.4]
  assign regs_312_reset = io_reset; // @[:@130232.4 RegFile.scala 76:16:@130239.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@130238.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@130242.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@130236.4]
  assign regs_313_clock = clock; // @[:@130245.4]
  assign regs_313_reset = io_reset; // @[:@130246.4 RegFile.scala 76:16:@130253.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@130252.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@130256.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@130250.4]
  assign regs_314_clock = clock; // @[:@130259.4]
  assign regs_314_reset = io_reset; // @[:@130260.4 RegFile.scala 76:16:@130267.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@130266.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@130270.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@130264.4]
  assign regs_315_clock = clock; // @[:@130273.4]
  assign regs_315_reset = io_reset; // @[:@130274.4 RegFile.scala 76:16:@130281.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@130280.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@130284.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@130278.4]
  assign regs_316_clock = clock; // @[:@130287.4]
  assign regs_316_reset = io_reset; // @[:@130288.4 RegFile.scala 76:16:@130295.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@130294.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@130298.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@130292.4]
  assign regs_317_clock = clock; // @[:@130301.4]
  assign regs_317_reset = io_reset; // @[:@130302.4 RegFile.scala 76:16:@130309.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@130308.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@130312.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@130306.4]
  assign regs_318_clock = clock; // @[:@130315.4]
  assign regs_318_reset = io_reset; // @[:@130316.4 RegFile.scala 76:16:@130323.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@130322.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@130326.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@130320.4]
  assign regs_319_clock = clock; // @[:@130329.4]
  assign regs_319_reset = io_reset; // @[:@130330.4 RegFile.scala 76:16:@130337.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@130336.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@130340.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@130334.4]
  assign regs_320_clock = clock; // @[:@130343.4]
  assign regs_320_reset = io_reset; // @[:@130344.4 RegFile.scala 76:16:@130351.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@130350.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@130354.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@130348.4]
  assign regs_321_clock = clock; // @[:@130357.4]
  assign regs_321_reset = io_reset; // @[:@130358.4 RegFile.scala 76:16:@130365.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@130364.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@130368.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@130362.4]
  assign regs_322_clock = clock; // @[:@130371.4]
  assign regs_322_reset = io_reset; // @[:@130372.4 RegFile.scala 76:16:@130379.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@130378.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@130382.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@130376.4]
  assign regs_323_clock = clock; // @[:@130385.4]
  assign regs_323_reset = io_reset; // @[:@130386.4 RegFile.scala 76:16:@130393.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@130392.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@130396.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@130390.4]
  assign regs_324_clock = clock; // @[:@130399.4]
  assign regs_324_reset = io_reset; // @[:@130400.4 RegFile.scala 76:16:@130407.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@130406.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@130410.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@130404.4]
  assign regs_325_clock = clock; // @[:@130413.4]
  assign regs_325_reset = io_reset; // @[:@130414.4 RegFile.scala 76:16:@130421.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@130420.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@130424.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@130418.4]
  assign regs_326_clock = clock; // @[:@130427.4]
  assign regs_326_reset = io_reset; // @[:@130428.4 RegFile.scala 76:16:@130435.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@130434.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@130438.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@130432.4]
  assign regs_327_clock = clock; // @[:@130441.4]
  assign regs_327_reset = io_reset; // @[:@130442.4 RegFile.scala 76:16:@130449.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@130448.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@130452.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@130446.4]
  assign regs_328_clock = clock; // @[:@130455.4]
  assign regs_328_reset = io_reset; // @[:@130456.4 RegFile.scala 76:16:@130463.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@130462.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@130466.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@130460.4]
  assign regs_329_clock = clock; // @[:@130469.4]
  assign regs_329_reset = io_reset; // @[:@130470.4 RegFile.scala 76:16:@130477.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@130476.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@130480.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@130474.4]
  assign regs_330_clock = clock; // @[:@130483.4]
  assign regs_330_reset = io_reset; // @[:@130484.4 RegFile.scala 76:16:@130491.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@130490.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@130494.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@130488.4]
  assign regs_331_clock = clock; // @[:@130497.4]
  assign regs_331_reset = io_reset; // @[:@130498.4 RegFile.scala 76:16:@130505.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@130504.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@130508.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@130502.4]
  assign regs_332_clock = clock; // @[:@130511.4]
  assign regs_332_reset = io_reset; // @[:@130512.4 RegFile.scala 76:16:@130519.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@130518.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@130522.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@130516.4]
  assign regs_333_clock = clock; // @[:@130525.4]
  assign regs_333_reset = io_reset; // @[:@130526.4 RegFile.scala 76:16:@130533.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@130532.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@130536.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@130530.4]
  assign regs_334_clock = clock; // @[:@130539.4]
  assign regs_334_reset = io_reset; // @[:@130540.4 RegFile.scala 76:16:@130547.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@130546.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@130550.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@130544.4]
  assign regs_335_clock = clock; // @[:@130553.4]
  assign regs_335_reset = io_reset; // @[:@130554.4 RegFile.scala 76:16:@130561.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@130560.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@130564.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@130558.4]
  assign regs_336_clock = clock; // @[:@130567.4]
  assign regs_336_reset = io_reset; // @[:@130568.4 RegFile.scala 76:16:@130575.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@130574.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@130578.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@130572.4]
  assign regs_337_clock = clock; // @[:@130581.4]
  assign regs_337_reset = io_reset; // @[:@130582.4 RegFile.scala 76:16:@130589.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@130588.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@130592.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@130586.4]
  assign regs_338_clock = clock; // @[:@130595.4]
  assign regs_338_reset = io_reset; // @[:@130596.4 RegFile.scala 76:16:@130603.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@130602.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@130606.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@130600.4]
  assign regs_339_clock = clock; // @[:@130609.4]
  assign regs_339_reset = io_reset; // @[:@130610.4 RegFile.scala 76:16:@130617.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@130616.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@130620.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@130614.4]
  assign regs_340_clock = clock; // @[:@130623.4]
  assign regs_340_reset = io_reset; // @[:@130624.4 RegFile.scala 76:16:@130631.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@130630.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@130634.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@130628.4]
  assign regs_341_clock = clock; // @[:@130637.4]
  assign regs_341_reset = io_reset; // @[:@130638.4 RegFile.scala 76:16:@130645.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@130644.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@130648.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@130642.4]
  assign regs_342_clock = clock; // @[:@130651.4]
  assign regs_342_reset = io_reset; // @[:@130652.4 RegFile.scala 76:16:@130659.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@130658.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@130662.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@130656.4]
  assign regs_343_clock = clock; // @[:@130665.4]
  assign regs_343_reset = io_reset; // @[:@130666.4 RegFile.scala 76:16:@130673.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@130672.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@130676.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@130670.4]
  assign regs_344_clock = clock; // @[:@130679.4]
  assign regs_344_reset = io_reset; // @[:@130680.4 RegFile.scala 76:16:@130687.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@130686.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@130690.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@130684.4]
  assign regs_345_clock = clock; // @[:@130693.4]
  assign regs_345_reset = io_reset; // @[:@130694.4 RegFile.scala 76:16:@130701.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@130700.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@130704.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@130698.4]
  assign regs_346_clock = clock; // @[:@130707.4]
  assign regs_346_reset = io_reset; // @[:@130708.4 RegFile.scala 76:16:@130715.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@130714.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@130718.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@130712.4]
  assign regs_347_clock = clock; // @[:@130721.4]
  assign regs_347_reset = io_reset; // @[:@130722.4 RegFile.scala 76:16:@130729.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@130728.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@130732.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@130726.4]
  assign regs_348_clock = clock; // @[:@130735.4]
  assign regs_348_reset = io_reset; // @[:@130736.4 RegFile.scala 76:16:@130743.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@130742.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@130746.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@130740.4]
  assign regs_349_clock = clock; // @[:@130749.4]
  assign regs_349_reset = io_reset; // @[:@130750.4 RegFile.scala 76:16:@130757.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@130756.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@130760.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@130754.4]
  assign regs_350_clock = clock; // @[:@130763.4]
  assign regs_350_reset = io_reset; // @[:@130764.4 RegFile.scala 76:16:@130771.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@130770.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@130774.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@130768.4]
  assign regs_351_clock = clock; // @[:@130777.4]
  assign regs_351_reset = io_reset; // @[:@130778.4 RegFile.scala 76:16:@130785.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@130784.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@130788.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@130782.4]
  assign regs_352_clock = clock; // @[:@130791.4]
  assign regs_352_reset = io_reset; // @[:@130792.4 RegFile.scala 76:16:@130799.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@130798.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@130802.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@130796.4]
  assign regs_353_clock = clock; // @[:@130805.4]
  assign regs_353_reset = io_reset; // @[:@130806.4 RegFile.scala 76:16:@130813.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@130812.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@130816.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@130810.4]
  assign regs_354_clock = clock; // @[:@130819.4]
  assign regs_354_reset = io_reset; // @[:@130820.4 RegFile.scala 76:16:@130827.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@130826.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@130830.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@130824.4]
  assign regs_355_clock = clock; // @[:@130833.4]
  assign regs_355_reset = io_reset; // @[:@130834.4 RegFile.scala 76:16:@130841.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@130840.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@130844.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@130838.4]
  assign regs_356_clock = clock; // @[:@130847.4]
  assign regs_356_reset = io_reset; // @[:@130848.4 RegFile.scala 76:16:@130855.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@130854.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@130858.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@130852.4]
  assign regs_357_clock = clock; // @[:@130861.4]
  assign regs_357_reset = io_reset; // @[:@130862.4 RegFile.scala 76:16:@130869.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@130868.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@130872.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@130866.4]
  assign regs_358_clock = clock; // @[:@130875.4]
  assign regs_358_reset = io_reset; // @[:@130876.4 RegFile.scala 76:16:@130883.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@130882.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@130886.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@130880.4]
  assign regs_359_clock = clock; // @[:@130889.4]
  assign regs_359_reset = io_reset; // @[:@130890.4 RegFile.scala 76:16:@130897.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@130896.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@130900.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@130894.4]
  assign regs_360_clock = clock; // @[:@130903.4]
  assign regs_360_reset = io_reset; // @[:@130904.4 RegFile.scala 76:16:@130911.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@130910.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@130914.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@130908.4]
  assign regs_361_clock = clock; // @[:@130917.4]
  assign regs_361_reset = io_reset; // @[:@130918.4 RegFile.scala 76:16:@130925.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@130924.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@130928.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@130922.4]
  assign regs_362_clock = clock; // @[:@130931.4]
  assign regs_362_reset = io_reset; // @[:@130932.4 RegFile.scala 76:16:@130939.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@130938.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@130942.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@130936.4]
  assign regs_363_clock = clock; // @[:@130945.4]
  assign regs_363_reset = io_reset; // @[:@130946.4 RegFile.scala 76:16:@130953.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@130952.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@130956.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@130950.4]
  assign regs_364_clock = clock; // @[:@130959.4]
  assign regs_364_reset = io_reset; // @[:@130960.4 RegFile.scala 76:16:@130967.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@130966.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@130970.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@130964.4]
  assign regs_365_clock = clock; // @[:@130973.4]
  assign regs_365_reset = io_reset; // @[:@130974.4 RegFile.scala 76:16:@130981.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@130980.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@130984.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@130978.4]
  assign regs_366_clock = clock; // @[:@130987.4]
  assign regs_366_reset = io_reset; // @[:@130988.4 RegFile.scala 76:16:@130995.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@130994.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@130998.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@130992.4]
  assign regs_367_clock = clock; // @[:@131001.4]
  assign regs_367_reset = io_reset; // @[:@131002.4 RegFile.scala 76:16:@131009.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@131008.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@131012.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@131006.4]
  assign regs_368_clock = clock; // @[:@131015.4]
  assign regs_368_reset = io_reset; // @[:@131016.4 RegFile.scala 76:16:@131023.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@131022.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@131026.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@131020.4]
  assign regs_369_clock = clock; // @[:@131029.4]
  assign regs_369_reset = io_reset; // @[:@131030.4 RegFile.scala 76:16:@131037.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@131036.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@131040.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@131034.4]
  assign regs_370_clock = clock; // @[:@131043.4]
  assign regs_370_reset = io_reset; // @[:@131044.4 RegFile.scala 76:16:@131051.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@131050.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@131054.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@131048.4]
  assign regs_371_clock = clock; // @[:@131057.4]
  assign regs_371_reset = io_reset; // @[:@131058.4 RegFile.scala 76:16:@131065.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@131064.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@131068.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@131062.4]
  assign regs_372_clock = clock; // @[:@131071.4]
  assign regs_372_reset = io_reset; // @[:@131072.4 RegFile.scala 76:16:@131079.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@131078.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@131082.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@131076.4]
  assign regs_373_clock = clock; // @[:@131085.4]
  assign regs_373_reset = io_reset; // @[:@131086.4 RegFile.scala 76:16:@131093.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@131092.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@131096.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@131090.4]
  assign regs_374_clock = clock; // @[:@131099.4]
  assign regs_374_reset = io_reset; // @[:@131100.4 RegFile.scala 76:16:@131107.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@131106.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@131110.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@131104.4]
  assign regs_375_clock = clock; // @[:@131113.4]
  assign regs_375_reset = io_reset; // @[:@131114.4 RegFile.scala 76:16:@131121.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@131120.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@131124.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@131118.4]
  assign regs_376_clock = clock; // @[:@131127.4]
  assign regs_376_reset = io_reset; // @[:@131128.4 RegFile.scala 76:16:@131135.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@131134.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@131138.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@131132.4]
  assign regs_377_clock = clock; // @[:@131141.4]
  assign regs_377_reset = io_reset; // @[:@131142.4 RegFile.scala 76:16:@131149.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@131148.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@131152.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@131146.4]
  assign regs_378_clock = clock; // @[:@131155.4]
  assign regs_378_reset = io_reset; // @[:@131156.4 RegFile.scala 76:16:@131163.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@131162.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@131166.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@131160.4]
  assign regs_379_clock = clock; // @[:@131169.4]
  assign regs_379_reset = io_reset; // @[:@131170.4 RegFile.scala 76:16:@131177.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@131176.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@131180.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@131174.4]
  assign regs_380_clock = clock; // @[:@131183.4]
  assign regs_380_reset = io_reset; // @[:@131184.4 RegFile.scala 76:16:@131191.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@131190.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@131194.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@131188.4]
  assign regs_381_clock = clock; // @[:@131197.4]
  assign regs_381_reset = io_reset; // @[:@131198.4 RegFile.scala 76:16:@131205.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@131204.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@131208.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@131202.4]
  assign regs_382_clock = clock; // @[:@131211.4]
  assign regs_382_reset = io_reset; // @[:@131212.4 RegFile.scala 76:16:@131219.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@131218.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@131222.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@131216.4]
  assign regs_383_clock = clock; // @[:@131225.4]
  assign regs_383_reset = io_reset; // @[:@131226.4 RegFile.scala 76:16:@131233.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@131232.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@131236.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@131230.4]
  assign regs_384_clock = clock; // @[:@131239.4]
  assign regs_384_reset = io_reset; // @[:@131240.4 RegFile.scala 76:16:@131247.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@131246.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@131250.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@131244.4]
  assign regs_385_clock = clock; // @[:@131253.4]
  assign regs_385_reset = io_reset; // @[:@131254.4 RegFile.scala 76:16:@131261.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@131260.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@131264.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@131258.4]
  assign regs_386_clock = clock; // @[:@131267.4]
  assign regs_386_reset = io_reset; // @[:@131268.4 RegFile.scala 76:16:@131275.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@131274.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@131278.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@131272.4]
  assign regs_387_clock = clock; // @[:@131281.4]
  assign regs_387_reset = io_reset; // @[:@131282.4 RegFile.scala 76:16:@131289.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@131288.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@131292.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@131286.4]
  assign regs_388_clock = clock; // @[:@131295.4]
  assign regs_388_reset = io_reset; // @[:@131296.4 RegFile.scala 76:16:@131303.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@131302.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@131306.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@131300.4]
  assign regs_389_clock = clock; // @[:@131309.4]
  assign regs_389_reset = io_reset; // @[:@131310.4 RegFile.scala 76:16:@131317.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@131316.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@131320.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@131314.4]
  assign regs_390_clock = clock; // @[:@131323.4]
  assign regs_390_reset = io_reset; // @[:@131324.4 RegFile.scala 76:16:@131331.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@131330.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@131334.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@131328.4]
  assign regs_391_clock = clock; // @[:@131337.4]
  assign regs_391_reset = io_reset; // @[:@131338.4 RegFile.scala 76:16:@131345.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@131344.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@131348.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@131342.4]
  assign regs_392_clock = clock; // @[:@131351.4]
  assign regs_392_reset = io_reset; // @[:@131352.4 RegFile.scala 76:16:@131359.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@131358.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@131362.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@131356.4]
  assign regs_393_clock = clock; // @[:@131365.4]
  assign regs_393_reset = io_reset; // @[:@131366.4 RegFile.scala 76:16:@131373.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@131372.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@131376.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@131370.4]
  assign regs_394_clock = clock; // @[:@131379.4]
  assign regs_394_reset = io_reset; // @[:@131380.4 RegFile.scala 76:16:@131387.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@131386.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@131390.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@131384.4]
  assign regs_395_clock = clock; // @[:@131393.4]
  assign regs_395_reset = io_reset; // @[:@131394.4 RegFile.scala 76:16:@131401.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@131400.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@131404.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@131398.4]
  assign regs_396_clock = clock; // @[:@131407.4]
  assign regs_396_reset = io_reset; // @[:@131408.4 RegFile.scala 76:16:@131415.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@131414.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@131418.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@131412.4]
  assign regs_397_clock = clock; // @[:@131421.4]
  assign regs_397_reset = io_reset; // @[:@131422.4 RegFile.scala 76:16:@131429.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@131428.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@131432.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@131426.4]
  assign regs_398_clock = clock; // @[:@131435.4]
  assign regs_398_reset = io_reset; // @[:@131436.4 RegFile.scala 76:16:@131443.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@131442.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@131446.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@131440.4]
  assign regs_399_clock = clock; // @[:@131449.4]
  assign regs_399_reset = io_reset; // @[:@131450.4 RegFile.scala 76:16:@131457.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@131456.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@131460.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@131454.4]
  assign regs_400_clock = clock; // @[:@131463.4]
  assign regs_400_reset = io_reset; // @[:@131464.4 RegFile.scala 76:16:@131471.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@131470.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@131474.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@131468.4]
  assign regs_401_clock = clock; // @[:@131477.4]
  assign regs_401_reset = io_reset; // @[:@131478.4 RegFile.scala 76:16:@131485.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@131484.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@131488.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@131482.4]
  assign regs_402_clock = clock; // @[:@131491.4]
  assign regs_402_reset = io_reset; // @[:@131492.4 RegFile.scala 76:16:@131499.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@131498.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@131502.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@131496.4]
  assign regs_403_clock = clock; // @[:@131505.4]
  assign regs_403_reset = io_reset; // @[:@131506.4 RegFile.scala 76:16:@131513.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@131512.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@131516.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@131510.4]
  assign regs_404_clock = clock; // @[:@131519.4]
  assign regs_404_reset = io_reset; // @[:@131520.4 RegFile.scala 76:16:@131527.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@131526.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@131530.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@131524.4]
  assign regs_405_clock = clock; // @[:@131533.4]
  assign regs_405_reset = io_reset; // @[:@131534.4 RegFile.scala 76:16:@131541.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@131540.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@131544.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@131538.4]
  assign regs_406_clock = clock; // @[:@131547.4]
  assign regs_406_reset = io_reset; // @[:@131548.4 RegFile.scala 76:16:@131555.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@131554.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@131558.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@131552.4]
  assign regs_407_clock = clock; // @[:@131561.4]
  assign regs_407_reset = io_reset; // @[:@131562.4 RegFile.scala 76:16:@131569.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@131568.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@131572.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@131566.4]
  assign regs_408_clock = clock; // @[:@131575.4]
  assign regs_408_reset = io_reset; // @[:@131576.4 RegFile.scala 76:16:@131583.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@131582.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@131586.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@131580.4]
  assign regs_409_clock = clock; // @[:@131589.4]
  assign regs_409_reset = io_reset; // @[:@131590.4 RegFile.scala 76:16:@131597.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@131596.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@131600.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@131594.4]
  assign regs_410_clock = clock; // @[:@131603.4]
  assign regs_410_reset = io_reset; // @[:@131604.4 RegFile.scala 76:16:@131611.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@131610.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@131614.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@131608.4]
  assign regs_411_clock = clock; // @[:@131617.4]
  assign regs_411_reset = io_reset; // @[:@131618.4 RegFile.scala 76:16:@131625.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@131624.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@131628.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@131622.4]
  assign regs_412_clock = clock; // @[:@131631.4]
  assign regs_412_reset = io_reset; // @[:@131632.4 RegFile.scala 76:16:@131639.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@131638.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@131642.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@131636.4]
  assign regs_413_clock = clock; // @[:@131645.4]
  assign regs_413_reset = io_reset; // @[:@131646.4 RegFile.scala 76:16:@131653.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@131652.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@131656.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@131650.4]
  assign regs_414_clock = clock; // @[:@131659.4]
  assign regs_414_reset = io_reset; // @[:@131660.4 RegFile.scala 76:16:@131667.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@131666.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@131670.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@131664.4]
  assign regs_415_clock = clock; // @[:@131673.4]
  assign regs_415_reset = io_reset; // @[:@131674.4 RegFile.scala 76:16:@131681.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@131680.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@131684.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@131678.4]
  assign regs_416_clock = clock; // @[:@131687.4]
  assign regs_416_reset = io_reset; // @[:@131688.4 RegFile.scala 76:16:@131695.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@131694.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@131698.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@131692.4]
  assign regs_417_clock = clock; // @[:@131701.4]
  assign regs_417_reset = io_reset; // @[:@131702.4 RegFile.scala 76:16:@131709.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@131708.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@131712.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@131706.4]
  assign regs_418_clock = clock; // @[:@131715.4]
  assign regs_418_reset = io_reset; // @[:@131716.4 RegFile.scala 76:16:@131723.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@131722.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@131726.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@131720.4]
  assign regs_419_clock = clock; // @[:@131729.4]
  assign regs_419_reset = io_reset; // @[:@131730.4 RegFile.scala 76:16:@131737.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@131736.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@131740.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@131734.4]
  assign regs_420_clock = clock; // @[:@131743.4]
  assign regs_420_reset = io_reset; // @[:@131744.4 RegFile.scala 76:16:@131751.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@131750.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@131754.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@131748.4]
  assign regs_421_clock = clock; // @[:@131757.4]
  assign regs_421_reset = io_reset; // @[:@131758.4 RegFile.scala 76:16:@131765.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@131764.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@131768.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@131762.4]
  assign regs_422_clock = clock; // @[:@131771.4]
  assign regs_422_reset = io_reset; // @[:@131772.4 RegFile.scala 76:16:@131779.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@131778.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@131782.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@131776.4]
  assign regs_423_clock = clock; // @[:@131785.4]
  assign regs_423_reset = io_reset; // @[:@131786.4 RegFile.scala 76:16:@131793.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@131792.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@131796.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@131790.4]
  assign regs_424_clock = clock; // @[:@131799.4]
  assign regs_424_reset = io_reset; // @[:@131800.4 RegFile.scala 76:16:@131807.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@131806.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@131810.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@131804.4]
  assign regs_425_clock = clock; // @[:@131813.4]
  assign regs_425_reset = io_reset; // @[:@131814.4 RegFile.scala 76:16:@131821.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@131820.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@131824.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@131818.4]
  assign regs_426_clock = clock; // @[:@131827.4]
  assign regs_426_reset = io_reset; // @[:@131828.4 RegFile.scala 76:16:@131835.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@131834.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@131838.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@131832.4]
  assign regs_427_clock = clock; // @[:@131841.4]
  assign regs_427_reset = io_reset; // @[:@131842.4 RegFile.scala 76:16:@131849.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@131848.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@131852.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@131846.4]
  assign regs_428_clock = clock; // @[:@131855.4]
  assign regs_428_reset = io_reset; // @[:@131856.4 RegFile.scala 76:16:@131863.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@131862.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@131866.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@131860.4]
  assign regs_429_clock = clock; // @[:@131869.4]
  assign regs_429_reset = io_reset; // @[:@131870.4 RegFile.scala 76:16:@131877.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@131876.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@131880.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@131874.4]
  assign regs_430_clock = clock; // @[:@131883.4]
  assign regs_430_reset = io_reset; // @[:@131884.4 RegFile.scala 76:16:@131891.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@131890.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@131894.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@131888.4]
  assign regs_431_clock = clock; // @[:@131897.4]
  assign regs_431_reset = io_reset; // @[:@131898.4 RegFile.scala 76:16:@131905.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@131904.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@131908.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@131902.4]
  assign regs_432_clock = clock; // @[:@131911.4]
  assign regs_432_reset = io_reset; // @[:@131912.4 RegFile.scala 76:16:@131919.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@131918.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@131922.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@131916.4]
  assign regs_433_clock = clock; // @[:@131925.4]
  assign regs_433_reset = io_reset; // @[:@131926.4 RegFile.scala 76:16:@131933.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@131932.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@131936.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@131930.4]
  assign regs_434_clock = clock; // @[:@131939.4]
  assign regs_434_reset = io_reset; // @[:@131940.4 RegFile.scala 76:16:@131947.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@131946.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@131950.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@131944.4]
  assign regs_435_clock = clock; // @[:@131953.4]
  assign regs_435_reset = io_reset; // @[:@131954.4 RegFile.scala 76:16:@131961.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@131960.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@131964.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@131958.4]
  assign regs_436_clock = clock; // @[:@131967.4]
  assign regs_436_reset = io_reset; // @[:@131968.4 RegFile.scala 76:16:@131975.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@131974.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@131978.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@131972.4]
  assign regs_437_clock = clock; // @[:@131981.4]
  assign regs_437_reset = io_reset; // @[:@131982.4 RegFile.scala 76:16:@131989.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@131988.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@131992.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@131986.4]
  assign regs_438_clock = clock; // @[:@131995.4]
  assign regs_438_reset = io_reset; // @[:@131996.4 RegFile.scala 76:16:@132003.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@132002.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@132006.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@132000.4]
  assign regs_439_clock = clock; // @[:@132009.4]
  assign regs_439_reset = io_reset; // @[:@132010.4 RegFile.scala 76:16:@132017.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@132016.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@132020.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@132014.4]
  assign regs_440_clock = clock; // @[:@132023.4]
  assign regs_440_reset = io_reset; // @[:@132024.4 RegFile.scala 76:16:@132031.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@132030.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@132034.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@132028.4]
  assign regs_441_clock = clock; // @[:@132037.4]
  assign regs_441_reset = io_reset; // @[:@132038.4 RegFile.scala 76:16:@132045.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@132044.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@132048.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@132042.4]
  assign regs_442_clock = clock; // @[:@132051.4]
  assign regs_442_reset = io_reset; // @[:@132052.4 RegFile.scala 76:16:@132059.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@132058.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@132062.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@132056.4]
  assign regs_443_clock = clock; // @[:@132065.4]
  assign regs_443_reset = io_reset; // @[:@132066.4 RegFile.scala 76:16:@132073.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@132072.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@132076.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@132070.4]
  assign regs_444_clock = clock; // @[:@132079.4]
  assign regs_444_reset = io_reset; // @[:@132080.4 RegFile.scala 76:16:@132087.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@132086.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@132090.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@132084.4]
  assign regs_445_clock = clock; // @[:@132093.4]
  assign regs_445_reset = io_reset; // @[:@132094.4 RegFile.scala 76:16:@132101.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@132100.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@132104.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@132098.4]
  assign regs_446_clock = clock; // @[:@132107.4]
  assign regs_446_reset = io_reset; // @[:@132108.4 RegFile.scala 76:16:@132115.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@132114.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@132118.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@132112.4]
  assign regs_447_clock = clock; // @[:@132121.4]
  assign regs_447_reset = io_reset; // @[:@132122.4 RegFile.scala 76:16:@132129.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@132128.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@132132.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@132126.4]
  assign regs_448_clock = clock; // @[:@132135.4]
  assign regs_448_reset = io_reset; // @[:@132136.4 RegFile.scala 76:16:@132143.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@132142.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@132146.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@132140.4]
  assign regs_449_clock = clock; // @[:@132149.4]
  assign regs_449_reset = io_reset; // @[:@132150.4 RegFile.scala 76:16:@132157.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@132156.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@132160.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@132154.4]
  assign regs_450_clock = clock; // @[:@132163.4]
  assign regs_450_reset = io_reset; // @[:@132164.4 RegFile.scala 76:16:@132171.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@132170.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@132174.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@132168.4]
  assign regs_451_clock = clock; // @[:@132177.4]
  assign regs_451_reset = io_reset; // @[:@132178.4 RegFile.scala 76:16:@132185.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@132184.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@132188.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@132182.4]
  assign regs_452_clock = clock; // @[:@132191.4]
  assign regs_452_reset = io_reset; // @[:@132192.4 RegFile.scala 76:16:@132199.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@132198.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@132202.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@132196.4]
  assign regs_453_clock = clock; // @[:@132205.4]
  assign regs_453_reset = io_reset; // @[:@132206.4 RegFile.scala 76:16:@132213.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@132212.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@132216.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@132210.4]
  assign regs_454_clock = clock; // @[:@132219.4]
  assign regs_454_reset = io_reset; // @[:@132220.4 RegFile.scala 76:16:@132227.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@132226.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@132230.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@132224.4]
  assign regs_455_clock = clock; // @[:@132233.4]
  assign regs_455_reset = io_reset; // @[:@132234.4 RegFile.scala 76:16:@132241.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@132240.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@132244.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@132238.4]
  assign regs_456_clock = clock; // @[:@132247.4]
  assign regs_456_reset = io_reset; // @[:@132248.4 RegFile.scala 76:16:@132255.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@132254.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@132258.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@132252.4]
  assign regs_457_clock = clock; // @[:@132261.4]
  assign regs_457_reset = io_reset; // @[:@132262.4 RegFile.scala 76:16:@132269.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@132268.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@132272.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@132266.4]
  assign regs_458_clock = clock; // @[:@132275.4]
  assign regs_458_reset = io_reset; // @[:@132276.4 RegFile.scala 76:16:@132283.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@132282.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@132286.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@132280.4]
  assign regs_459_clock = clock; // @[:@132289.4]
  assign regs_459_reset = io_reset; // @[:@132290.4 RegFile.scala 76:16:@132297.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@132296.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@132300.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@132294.4]
  assign regs_460_clock = clock; // @[:@132303.4]
  assign regs_460_reset = io_reset; // @[:@132304.4 RegFile.scala 76:16:@132311.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@132310.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@132314.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@132308.4]
  assign regs_461_clock = clock; // @[:@132317.4]
  assign regs_461_reset = io_reset; // @[:@132318.4 RegFile.scala 76:16:@132325.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@132324.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@132328.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@132322.4]
  assign regs_462_clock = clock; // @[:@132331.4]
  assign regs_462_reset = io_reset; // @[:@132332.4 RegFile.scala 76:16:@132339.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@132338.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@132342.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@132336.4]
  assign regs_463_clock = clock; // @[:@132345.4]
  assign regs_463_reset = io_reset; // @[:@132346.4 RegFile.scala 76:16:@132353.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@132352.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@132356.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@132350.4]
  assign regs_464_clock = clock; // @[:@132359.4]
  assign regs_464_reset = io_reset; // @[:@132360.4 RegFile.scala 76:16:@132367.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@132366.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@132370.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@132364.4]
  assign regs_465_clock = clock; // @[:@132373.4]
  assign regs_465_reset = io_reset; // @[:@132374.4 RegFile.scala 76:16:@132381.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@132380.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@132384.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@132378.4]
  assign regs_466_clock = clock; // @[:@132387.4]
  assign regs_466_reset = io_reset; // @[:@132388.4 RegFile.scala 76:16:@132395.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@132394.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@132398.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@132392.4]
  assign regs_467_clock = clock; // @[:@132401.4]
  assign regs_467_reset = io_reset; // @[:@132402.4 RegFile.scala 76:16:@132409.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@132408.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@132412.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@132406.4]
  assign regs_468_clock = clock; // @[:@132415.4]
  assign regs_468_reset = io_reset; // @[:@132416.4 RegFile.scala 76:16:@132423.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@132422.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@132426.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@132420.4]
  assign regs_469_clock = clock; // @[:@132429.4]
  assign regs_469_reset = io_reset; // @[:@132430.4 RegFile.scala 76:16:@132437.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@132436.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@132440.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@132434.4]
  assign regs_470_clock = clock; // @[:@132443.4]
  assign regs_470_reset = io_reset; // @[:@132444.4 RegFile.scala 76:16:@132451.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@132450.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@132454.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@132448.4]
  assign regs_471_clock = clock; // @[:@132457.4]
  assign regs_471_reset = io_reset; // @[:@132458.4 RegFile.scala 76:16:@132465.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@132464.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@132468.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@132462.4]
  assign regs_472_clock = clock; // @[:@132471.4]
  assign regs_472_reset = io_reset; // @[:@132472.4 RegFile.scala 76:16:@132479.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@132478.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@132482.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@132476.4]
  assign regs_473_clock = clock; // @[:@132485.4]
  assign regs_473_reset = io_reset; // @[:@132486.4 RegFile.scala 76:16:@132493.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@132492.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@132496.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@132490.4]
  assign regs_474_clock = clock; // @[:@132499.4]
  assign regs_474_reset = io_reset; // @[:@132500.4 RegFile.scala 76:16:@132507.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@132506.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@132510.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@132504.4]
  assign regs_475_clock = clock; // @[:@132513.4]
  assign regs_475_reset = io_reset; // @[:@132514.4 RegFile.scala 76:16:@132521.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@132520.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@132524.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@132518.4]
  assign regs_476_clock = clock; // @[:@132527.4]
  assign regs_476_reset = io_reset; // @[:@132528.4 RegFile.scala 76:16:@132535.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@132534.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@132538.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@132532.4]
  assign regs_477_clock = clock; // @[:@132541.4]
  assign regs_477_reset = io_reset; // @[:@132542.4 RegFile.scala 76:16:@132549.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@132548.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@132552.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@132546.4]
  assign regs_478_clock = clock; // @[:@132555.4]
  assign regs_478_reset = io_reset; // @[:@132556.4 RegFile.scala 76:16:@132563.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@132562.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@132566.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@132560.4]
  assign regs_479_clock = clock; // @[:@132569.4]
  assign regs_479_reset = io_reset; // @[:@132570.4 RegFile.scala 76:16:@132577.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@132576.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@132580.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@132574.4]
  assign regs_480_clock = clock; // @[:@132583.4]
  assign regs_480_reset = io_reset; // @[:@132584.4 RegFile.scala 76:16:@132591.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@132590.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@132594.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@132588.4]
  assign regs_481_clock = clock; // @[:@132597.4]
  assign regs_481_reset = io_reset; // @[:@132598.4 RegFile.scala 76:16:@132605.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@132604.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@132608.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@132602.4]
  assign regs_482_clock = clock; // @[:@132611.4]
  assign regs_482_reset = io_reset; // @[:@132612.4 RegFile.scala 76:16:@132619.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@132618.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@132622.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@132616.4]
  assign regs_483_clock = clock; // @[:@132625.4]
  assign regs_483_reset = io_reset; // @[:@132626.4 RegFile.scala 76:16:@132633.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@132632.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@132636.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@132630.4]
  assign regs_484_clock = clock; // @[:@132639.4]
  assign regs_484_reset = io_reset; // @[:@132640.4 RegFile.scala 76:16:@132647.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@132646.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@132650.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@132644.4]
  assign regs_485_clock = clock; // @[:@132653.4]
  assign regs_485_reset = io_reset; // @[:@132654.4 RegFile.scala 76:16:@132661.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@132660.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@132664.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@132658.4]
  assign regs_486_clock = clock; // @[:@132667.4]
  assign regs_486_reset = io_reset; // @[:@132668.4 RegFile.scala 76:16:@132675.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@132674.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@132678.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@132672.4]
  assign regs_487_clock = clock; // @[:@132681.4]
  assign regs_487_reset = io_reset; // @[:@132682.4 RegFile.scala 76:16:@132689.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@132688.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@132692.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@132686.4]
  assign regs_488_clock = clock; // @[:@132695.4]
  assign regs_488_reset = io_reset; // @[:@132696.4 RegFile.scala 76:16:@132703.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@132702.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@132706.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@132700.4]
  assign regs_489_clock = clock; // @[:@132709.4]
  assign regs_489_reset = io_reset; // @[:@132710.4 RegFile.scala 76:16:@132717.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@132716.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@132720.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@132714.4]
  assign regs_490_clock = clock; // @[:@132723.4]
  assign regs_490_reset = io_reset; // @[:@132724.4 RegFile.scala 76:16:@132731.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@132730.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@132734.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@132728.4]
  assign regs_491_clock = clock; // @[:@132737.4]
  assign regs_491_reset = io_reset; // @[:@132738.4 RegFile.scala 76:16:@132745.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@132744.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@132748.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@132742.4]
  assign regs_492_clock = clock; // @[:@132751.4]
  assign regs_492_reset = io_reset; // @[:@132752.4 RegFile.scala 76:16:@132759.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@132758.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@132762.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@132756.4]
  assign regs_493_clock = clock; // @[:@132765.4]
  assign regs_493_reset = io_reset; // @[:@132766.4 RegFile.scala 76:16:@132773.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@132772.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@132776.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@132770.4]
  assign regs_494_clock = clock; // @[:@132779.4]
  assign regs_494_reset = io_reset; // @[:@132780.4 RegFile.scala 76:16:@132787.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@132786.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@132790.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@132784.4]
  assign regs_495_clock = clock; // @[:@132793.4]
  assign regs_495_reset = io_reset; // @[:@132794.4 RegFile.scala 76:16:@132801.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@132800.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@132804.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@132798.4]
  assign regs_496_clock = clock; // @[:@132807.4]
  assign regs_496_reset = io_reset; // @[:@132808.4 RegFile.scala 76:16:@132815.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@132814.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@132818.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@132812.4]
  assign regs_497_clock = clock; // @[:@132821.4]
  assign regs_497_reset = io_reset; // @[:@132822.4 RegFile.scala 76:16:@132829.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@132828.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@132832.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@132826.4]
  assign regs_498_clock = clock; // @[:@132835.4]
  assign regs_498_reset = io_reset; // @[:@132836.4 RegFile.scala 76:16:@132843.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@132842.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@132846.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@132840.4]
  assign regs_499_clock = clock; // @[:@132849.4]
  assign regs_499_reset = io_reset; // @[:@132850.4 RegFile.scala 76:16:@132857.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@132856.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@132860.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@132854.4]
  assign regs_500_clock = clock; // @[:@132863.4]
  assign regs_500_reset = io_reset; // @[:@132864.4 RegFile.scala 76:16:@132871.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@132870.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@132874.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@132868.4]
  assign regs_501_clock = clock; // @[:@132877.4]
  assign regs_501_reset = io_reset; // @[:@132878.4 RegFile.scala 76:16:@132885.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@132884.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@132888.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@132882.4]
  assign regs_502_clock = clock; // @[:@132891.4]
  assign regs_502_reset = io_reset; // @[:@132892.4 RegFile.scala 76:16:@132899.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@132898.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@132902.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@132896.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@133411.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@133412.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@133413.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@133414.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@133415.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@133416.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@133417.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@133418.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@133419.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@133420.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@133421.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@133422.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@133423.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@133424.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@133425.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@133426.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@133427.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@133428.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@133429.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@133430.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@133431.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@133432.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@133433.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@133434.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@133435.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@133436.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@133437.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@133438.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@133439.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@133440.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@133441.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@133442.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@133443.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@133444.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@133445.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@133446.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@133447.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@133448.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@133449.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@133450.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@133451.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@133452.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@133453.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@133454.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@133455.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@133456.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@133457.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@133458.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@133459.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@133460.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@133461.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@133462.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@133463.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@133464.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@133465.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@133466.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@133467.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@133468.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@133469.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@133470.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@133471.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@133472.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@133473.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@133474.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@133475.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@133476.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@133477.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@133478.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@133479.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@133480.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@133481.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@133482.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@133483.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@133484.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@133485.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@133486.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@133487.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@133488.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@133489.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@133490.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@133491.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@133492.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@133493.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@133494.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@133495.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@133496.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@133497.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@133498.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@133499.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@133500.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@133501.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@133502.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@133503.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@133504.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@133505.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@133506.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@133507.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@133508.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@133509.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@133510.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@133511.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@133512.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@133513.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@133514.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@133515.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@133516.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@133517.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@133518.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@133519.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@133520.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@133521.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@133522.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@133523.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@133524.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@133525.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@133526.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@133527.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@133528.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@133529.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@133530.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@133531.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@133532.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@133533.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@133534.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@133535.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@133536.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@133537.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@133538.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@133539.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@133540.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@133541.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@133542.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@133543.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@133544.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@133545.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@133546.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@133547.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@133548.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@133549.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@133550.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@133551.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@133552.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@133553.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@133554.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@133555.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@133556.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@133557.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@133558.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@133559.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@133560.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@133561.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@133562.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@133563.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@133564.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@133565.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@133566.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@133567.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@133568.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@133569.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@133570.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@133571.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@133572.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@133573.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@133574.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@133575.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@133576.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@133577.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@133578.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@133579.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@133580.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@133581.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@133582.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@133583.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@133584.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@133585.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@133586.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@133587.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@133588.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@133589.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@133590.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@133591.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@133592.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@133593.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@133594.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@133595.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@133596.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@133597.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@133598.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@133599.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@133600.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@133601.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@133602.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@133603.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@133604.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@133605.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@133606.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@133607.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@133608.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@133609.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@133610.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@133611.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@133612.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@133613.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@133614.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@133615.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@133616.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@133617.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@133618.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@133619.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@133620.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@133621.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@133622.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@133623.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@133624.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@133625.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@133626.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@133627.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@133628.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@133629.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@133630.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@133631.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@133632.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@133633.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@133634.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@133635.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@133636.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@133637.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@133638.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@133639.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@133640.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@133641.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@133642.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@133643.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@133644.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@133645.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@133646.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@133647.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@133648.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@133649.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@133650.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@133651.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@133652.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@133653.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@133654.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@133655.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@133656.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@133657.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@133658.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@133659.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@133660.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@133661.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@133662.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@133663.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@133664.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@133665.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@133666.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@133667.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@133668.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@133669.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@133670.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@133671.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@133672.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@133673.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@133674.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@133675.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@133676.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@133677.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@133678.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@133679.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@133680.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@133681.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@133682.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@133683.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@133684.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@133685.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@133686.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@133687.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@133688.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@133689.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@133690.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@133691.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@133692.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@133693.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@133694.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@133695.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@133696.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@133697.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@133698.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@133699.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@133700.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@133701.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@133702.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@133703.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@133704.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@133705.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@133706.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@133707.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@133708.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@133709.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@133710.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@133711.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@133712.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@133713.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@133714.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@133715.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@133716.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@133717.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@133718.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@133719.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@133720.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@133721.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@133722.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@133723.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@133724.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@133725.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@133726.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@133727.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@133728.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@133729.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@133730.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@133731.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@133732.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@133733.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@133734.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@133735.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@133736.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@133737.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@133738.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@133739.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@133740.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@133741.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@133742.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@133743.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@133744.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@133745.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@133746.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@133747.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@133748.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@133749.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@133750.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@133751.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@133752.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@133753.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@133754.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@133755.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@133756.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@133757.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@133758.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@133759.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@133760.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@133761.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@133762.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@133763.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@133764.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@133765.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@133766.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@133767.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@133768.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@133769.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@133770.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@133771.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@133772.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@133773.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@133774.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@133775.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@133776.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@133777.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@133778.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@133779.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@133780.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@133781.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@133782.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@133783.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@133784.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@133785.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@133786.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@133787.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@133788.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@133789.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@133790.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@133791.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@133792.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@133793.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@133794.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@133795.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@133796.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@133797.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@133798.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@133799.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@133800.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@133801.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@133802.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@133803.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@133804.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@133805.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@133806.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@133807.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@133808.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@133809.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@133810.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@133811.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@133812.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@133813.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@133814.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@133815.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@133816.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@133817.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@133818.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@133819.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@133820.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@133821.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@133822.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@133823.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@133824.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@133825.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@133826.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@133827.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@133828.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@133829.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@133830.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@133831.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@133832.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@133833.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@133834.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@133835.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@133836.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@133837.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@133838.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@133839.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@133840.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@133841.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@133842.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@133843.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@133844.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@133845.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@133846.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@133847.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@133848.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@133849.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@133850.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@133851.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@133852.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@133853.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@133854.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@133855.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@133856.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@133857.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@133858.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@133859.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@133860.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@133861.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@133862.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@133863.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@133864.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@133865.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@133866.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@133867.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@133868.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@133869.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@133870.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@133871.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@133872.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@133873.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@133874.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@133875.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@133876.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@133877.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@133878.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@133879.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@133880.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@133881.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@133882.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@133883.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@133884.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@133885.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@133886.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@133887.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@133888.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@133889.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@133890.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@133891.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@133892.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@133893.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@133894.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@133895.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@133896.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@133897.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@133898.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@133899.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@133900.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@133901.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@133902.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@133903.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@133904.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@133905.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@133906.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@133907.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@133908.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@133909.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@133910.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@133911.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@133912.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@133913.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@133914.4]
endmodule
module RetimeWrapper_838( // @[:@133938.2]
  input         clock, // @[:@133939.4]
  input         reset, // @[:@133940.4]
  input  [39:0] io_in, // @[:@133941.4]
  output [39:0] io_out // @[:@133941.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@133943.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@133943.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@133943.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@133943.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@133943.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@133943.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@133943.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@133956.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@133955.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@133954.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@133953.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@133952.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@133950.4]
endmodule
module FringeFF_503( // @[:@133958.2]
  input         clock, // @[:@133959.4]
  input         reset, // @[:@133960.4]
  input  [39:0] io_in, // @[:@133961.4]
  output [39:0] io_out, // @[:@133961.4]
  input         io_enable // @[:@133961.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@133964.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@133964.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@133964.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@133964.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@133969.4 package.scala 96:25:@133970.4]
  RetimeWrapper_838 RetimeWrapper ( // @[package.scala 93:22:@133964.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@133969.4 package.scala 96:25:@133970.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@133981.4]
  assign RetimeWrapper_clock = clock; // @[:@133965.4]
  assign RetimeWrapper_reset = reset; // @[:@133966.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@133967.4]
endmodule
module FringeCounter( // @[:@133983.2]
  input   clock, // @[:@133984.4]
  input   reset, // @[:@133985.4]
  input   io_enable, // @[:@133986.4]
  output  io_done // @[:@133986.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@133988.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@133988.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@133988.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@133988.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@133988.4]
  wire [40:0] count; // @[Cat.scala 30:58:@133995.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@133996.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@133997.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@133998.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@134000.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@133988.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@133995.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@133996.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@133997.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@133998.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@134000.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@134011.4]
  assign reg$_clock = clock; // @[:@133989.4]
  assign reg$_reset = reset; // @[:@133990.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@134002.6 FringeCounter.scala 37:15:@134005.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@133993.4]
endmodule
module FringeFF_504( // @[:@134045.2]
  input   clock, // @[:@134046.4]
  input   reset, // @[:@134047.4]
  input   io_in, // @[:@134048.4]
  input   io_reset, // @[:@134048.4]
  output  io_out, // @[:@134048.4]
  input   io_enable // @[:@134048.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@134051.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@134051.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@134051.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@134051.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@134051.4]
  wire  _T_18; // @[package.scala 96:25:@134056.4 package.scala 96:25:@134057.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@134062.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@134051.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@134056.4 package.scala 96:25:@134057.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@134062.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@134068.4]
  assign RetimeWrapper_clock = clock; // @[:@134052.4]
  assign RetimeWrapper_reset = reset; // @[:@134053.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@134055.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@134054.4]
endmodule
module Depulser( // @[:@134070.2]
  input   clock, // @[:@134071.4]
  input   reset, // @[:@134072.4]
  input   io_in, // @[:@134073.4]
  input   io_rst, // @[:@134073.4]
  output  io_out // @[:@134073.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@134075.4]
  wire  r_reset; // @[Depulser.scala 14:17:@134075.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@134075.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@134075.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@134075.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@134075.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@134075.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@134084.4]
  assign r_clock = clock; // @[:@134076.4]
  assign r_reset = reset; // @[:@134077.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@134079.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@134083.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@134082.4]
endmodule
module Fringe( // @[:@134086.2]
  input         clock, // @[:@134087.4]
  input         reset, // @[:@134088.4]
  input  [31:0] io_raddr, // @[:@134089.4]
  input         io_wen, // @[:@134089.4]
  input  [31:0] io_waddr, // @[:@134089.4]
  input  [63:0] io_wdata, // @[:@134089.4]
  output [63:0] io_rdata, // @[:@134089.4]
  output        io_enable, // @[:@134089.4]
  input         io_done, // @[:@134089.4]
  output        io_reset, // @[:@134089.4]
  output [63:0] io_argIns_0, // @[:@134089.4]
  output [63:0] io_argIns_1, // @[:@134089.4]
  input         io_argOuts_0_valid, // @[:@134089.4]
  input  [63:0] io_argOuts_0_bits, // @[:@134089.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@134089.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@134089.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@134089.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@134089.4]
  output        io_memStreams_stores_0_data_ready, // @[:@134089.4]
  input         io_memStreams_stores_0_data_valid, // @[:@134089.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@134089.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@134089.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@134089.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@134089.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@134089.4]
  input         io_dram_0_cmd_ready, // @[:@134089.4]
  output        io_dram_0_cmd_valid, // @[:@134089.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@134089.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@134089.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@134089.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@134089.4]
  input         io_dram_0_wdata_ready, // @[:@134089.4]
  output        io_dram_0_wdata_valid, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@134089.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@134089.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@134089.4]
  output        io_dram_0_rresp_ready, // @[:@134089.4]
  output        io_dram_0_wresp_ready, // @[:@134089.4]
  input         io_dram_0_wresp_valid, // @[:@134089.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@134089.4]
  input         io_dram_1_cmd_ready, // @[:@134089.4]
  output        io_dram_1_cmd_valid, // @[:@134089.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@134089.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@134089.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@134089.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@134089.4]
  input         io_dram_1_wdata_ready, // @[:@134089.4]
  output        io_dram_1_wdata_valid, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@134089.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@134089.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@134089.4]
  output        io_dram_1_rresp_ready, // @[:@134089.4]
  output        io_dram_1_wresp_ready, // @[:@134089.4]
  input         io_dram_1_wresp_valid, // @[:@134089.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@134089.4]
  input         io_dram_2_cmd_ready, // @[:@134089.4]
  output        io_dram_2_cmd_valid, // @[:@134089.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@134089.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@134089.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@134089.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@134089.4]
  input         io_dram_2_wdata_ready, // @[:@134089.4]
  output        io_dram_2_wdata_valid, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@134089.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@134089.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@134089.4]
  output        io_dram_2_rresp_ready, // @[:@134089.4]
  output        io_dram_2_wresp_ready, // @[:@134089.4]
  input         io_dram_2_wresp_valid, // @[:@134089.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@134089.4]
  input         io_dram_3_cmd_ready, // @[:@134089.4]
  output        io_dram_3_cmd_valid, // @[:@134089.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@134089.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@134089.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@134089.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@134089.4]
  input         io_dram_3_wdata_ready, // @[:@134089.4]
  output        io_dram_3_wdata_valid, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@134089.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@134089.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@134089.4]
  output        io_dram_3_rresp_ready, // @[:@134089.4]
  output        io_dram_3_wresp_ready, // @[:@134089.4]
  input         io_dram_3_wresp_valid, // @[:@134089.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@134089.4]
  input         io_heap_0_req_valid, // @[:@134089.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@134089.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@134089.4]
  output        io_heap_0_resp_valid, // @[:@134089.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@134089.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@134089.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@134095.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@134095.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@134095.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@134095.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@135088.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@135088.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@135088.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@136048.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@136048.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@136048.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@137008.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@137008.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@137008.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@137008.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@137968.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@137968.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@137968.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@137968.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@137968.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@137968.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@137977.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@137977.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@137977.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@137977.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@137977.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@137977.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@137977.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@137977.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@137977.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@140027.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@140027.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@140027.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@140027.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@140046.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@140046.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@140046.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@140046.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@140046.4]
  wire [63:0] _T_1020; // @[:@140004.4 :@140005.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@140006.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@140008.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@140010.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@140012.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@140014.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@140016.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@140018.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@140054.4]
  reg  _T_1047; // @[package.scala 152:20:@140057.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@140059.4]
  wire  _T_1049; // @[package.scala 153:8:@140060.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@140064.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@140065.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@140068.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@140069.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@140071.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@140072.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@140074.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@140077.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@140056.4 Fringe.scala 163:24:@140075.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@140056.4 Fringe.scala 162:28:@140073.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@140078.4]
  wire  alloc; // @[Fringe.scala 202:38:@141708.4]
  wire  dealloc; // @[Fringe.scala 203:40:@141709.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@141710.4]
  reg  _T_1572; // @[package.scala 152:20:@141711.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@141713.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@134095.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@135088.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@136048.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@137008.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@137968.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@137977.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@140027.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@140046.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@140004.4 :@140005.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@140006.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@140008.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@140010.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@140012.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@140014.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@140016.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@140018.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@140054.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@140059.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@140060.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@140064.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@140065.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@140068.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@140069.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@140071.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@140072.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@140074.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@140077.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@140056.4 Fringe.scala 163:24:@140075.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@140056.4 Fringe.scala 162:28:@140073.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@140078.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@141708.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@141709.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@141710.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@141713.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@140002.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@140022.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@140023.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@140044.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@140045.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@135014.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@135010.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@135005.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@135004.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@141206.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@141205.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@141204.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@141202.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@141201.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@141199.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@141183.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@141184.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@141185.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@141186.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@141187.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@141188.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@141189.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@141190.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@141191.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@141192.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@141193.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@141194.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@141195.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@141196.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@141197.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@141198.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@141119.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@141120.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@141121.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@141122.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@141123.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@141124.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@141125.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@141126.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@141127.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@141128.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@141129.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@141130.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@141131.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@141132.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@141133.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@141134.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@141135.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@141136.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@141137.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@141138.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@141139.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@141140.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@141141.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@141142.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@141143.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@141144.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@141145.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@141146.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@141147.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@141148.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@141149.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@141150.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@141151.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@141152.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@141153.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@141154.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@141155.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@141156.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@141157.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@141158.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@141159.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@141160.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@141161.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@141162.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@141163.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@141164.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@141165.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@141166.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@141167.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@141168.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@141169.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@141170.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@141171.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@141172.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@141173.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@141174.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@141175.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@141176.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@141177.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@141178.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@141179.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@141180.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@141181.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@141182.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@141118.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@141117.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@141098.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@141318.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@141317.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@141316.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@141314.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@141313.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@141311.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@141295.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@141296.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@141297.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@141298.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@141299.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@141300.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@141301.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@141302.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@141303.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@141304.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@141305.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@141306.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@141307.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@141308.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@141309.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@141310.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@141231.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@141232.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@141233.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@141234.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@141235.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@141236.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@141237.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@141238.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@141239.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@141240.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@141241.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@141242.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@141243.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@141244.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@141245.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@141246.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@141247.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@141248.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@141249.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@141250.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@141251.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@141252.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@141253.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@141254.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@141255.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@141256.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@141257.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@141258.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@141259.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@141260.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@141261.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@141262.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@141263.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@141264.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@141265.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@141266.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@141267.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@141268.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@141269.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@141270.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@141271.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@141272.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@141273.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@141274.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@141275.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@141276.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@141277.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@141278.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@141279.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@141280.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@141281.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@141282.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@141283.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@141284.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@141285.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@141286.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@141287.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@141288.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@141289.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@141290.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@141291.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@141292.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@141293.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@141294.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@141230.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@141229.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@141210.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@141430.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@141429.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@141428.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@141426.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@141425.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@141423.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@141407.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@141408.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@141409.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@141410.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@141411.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@141412.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@141413.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@141414.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@141415.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@141416.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@141417.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@141418.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@141419.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@141420.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@141421.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@141422.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@141343.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@141344.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@141345.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@141346.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@141347.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@141348.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@141349.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@141350.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@141351.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@141352.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@141353.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@141354.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@141355.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@141356.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@141357.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@141358.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@141359.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@141360.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@141361.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@141362.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@141363.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@141364.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@141365.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@141366.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@141367.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@141368.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@141369.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@141370.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@141371.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@141372.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@141373.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@141374.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@141375.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@141376.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@141377.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@141378.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@141379.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@141380.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@141381.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@141382.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@141383.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@141384.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@141385.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@141386.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@141387.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@141388.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@141389.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@141390.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@141391.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@141392.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@141393.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@141394.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@141395.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@141396.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@141397.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@141398.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@141399.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@141400.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@141401.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@141402.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@141403.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@141404.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@141405.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@141406.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@141342.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@141341.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@141322.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@141542.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@141541.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@141540.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@141538.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@141537.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@141535.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@141519.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@141520.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@141521.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@141522.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@141523.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@141524.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@141525.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@141526.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@141527.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@141528.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@141529.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@141530.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@141531.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@141532.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@141533.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@141534.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@141455.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@141456.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@141457.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@141458.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@141459.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@141460.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@141461.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@141462.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@141463.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@141464.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@141465.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@141466.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@141467.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@141468.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@141469.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@141470.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@141471.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@141472.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@141473.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@141474.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@141475.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@141476.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@141477.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@141478.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@141479.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@141480.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@141481.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@141482.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@141483.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@141484.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@141485.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@141486.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@141487.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@141488.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@141489.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@141490.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@141491.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@141492.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@141493.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@141494.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@141495.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@141496.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@141497.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@141498.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@141499.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@141500.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@141501.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@141502.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@141503.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@141504.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@141505.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@141506.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@141507.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@141508.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@141509.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@141510.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@141511.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@141512.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@141513.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@141514.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@141515.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@141516.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@141517.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@141518.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@141454.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@141453.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@141434.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@137973.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@137972.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@137971.4]
  assign dramArbs_0_clock = clock; // @[:@134096.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@134097.4 Fringe.scala 187:30:@141088.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@141092.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@135013.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@135012.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@135011.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@135009.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@135008.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@135007.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@135006.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@141207.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@141200.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@141097.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@141096.4]
  assign dramArbs_1_clock = clock; // @[:@135089.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@135090.4 Fringe.scala 187:30:@141089.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@141093.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@141319.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@141312.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@141209.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@141208.4]
  assign dramArbs_2_clock = clock; // @[:@136049.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@136050.4 Fringe.scala 187:30:@141090.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@141094.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@141431.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@141424.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@141321.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@141320.4]
  assign dramArbs_3_clock = clock; // @[:@137009.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@137010.4 Fringe.scala 187:30:@141091.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@141095.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@141543.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@141536.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@141433.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@141432.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@137976.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@137975.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@137974.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@141715.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@141716.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@141717.4]
  assign regs_clock = clock; // @[:@137978.4]
  assign regs_reset = reset; // @[:@137979.4 Fringe.scala 139:14:@140026.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@139998.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@140000.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@139999.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@140001.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@140024.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@140076.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@140080.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@140083.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@140082.4]
  assign timeoutCtr_clock = clock; // @[:@140028.4]
  assign timeoutCtr_reset = reset; // @[:@140029.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@140043.4]
  assign depulser_clock = clock; // @[:@140047.4]
  assign depulser_reset = reset; // @[:@140048.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@140053.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@140055.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@141732.2]
  input         clock, // @[:@141733.4]
  input         reset, // @[:@141734.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@141735.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@141735.4]
  input         io_S_AXI_AWVALID, // @[:@141735.4]
  output        io_S_AXI_AWREADY, // @[:@141735.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@141735.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@141735.4]
  input         io_S_AXI_ARVALID, // @[:@141735.4]
  output        io_S_AXI_ARREADY, // @[:@141735.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@141735.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@141735.4]
  input         io_S_AXI_WVALID, // @[:@141735.4]
  output        io_S_AXI_WREADY, // @[:@141735.4]
  output [31:0] io_S_AXI_RDATA, // @[:@141735.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@141735.4]
  output        io_S_AXI_RVALID, // @[:@141735.4]
  input         io_S_AXI_RREADY, // @[:@141735.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@141735.4]
  output        io_S_AXI_BVALID, // @[:@141735.4]
  input         io_S_AXI_BREADY, // @[:@141735.4]
  output [31:0] io_raddr, // @[:@141735.4]
  output        io_wen, // @[:@141735.4]
  output [31:0] io_waddr, // @[:@141735.4]
  output [31:0] io_wdata, // @[:@141735.4]
  input  [31:0] io_rdata // @[:@141735.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@141737.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@141761.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@141757.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@141753.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@141752.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@141751.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@141750.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@141748.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@141747.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@141769.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@141772.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@141770.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@141771.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@141773.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@141768.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@141765.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@141764.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@141763.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@141762.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@141760.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@141759.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@141758.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@141756.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@141755.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@141754.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@141749.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@141746.4]
endmodule
module MAGToAXI4Bridge( // @[:@141775.2]
  output         io_in_cmd_ready, // @[:@141778.4]
  input          io_in_cmd_valid, // @[:@141778.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@141778.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@141778.4]
  input          io_in_cmd_bits_isWr, // @[:@141778.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@141778.4]
  output         io_in_wdata_ready, // @[:@141778.4]
  input          io_in_wdata_valid, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@141778.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@141778.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@141778.4]
  input          io_in_wdata_bits_wlast, // @[:@141778.4]
  input          io_in_rresp_ready, // @[:@141778.4]
  input          io_in_wresp_ready, // @[:@141778.4]
  output         io_in_wresp_valid, // @[:@141778.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@141778.4]
  output [31:0]  io_M_AXI_AWID, // @[:@141778.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@141778.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@141778.4]
  output         io_M_AXI_AWVALID, // @[:@141778.4]
  input          io_M_AXI_AWREADY, // @[:@141778.4]
  output [31:0]  io_M_AXI_ARID, // @[:@141778.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@141778.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@141778.4]
  output         io_M_AXI_ARVALID, // @[:@141778.4]
  input          io_M_AXI_ARREADY, // @[:@141778.4]
  output [511:0] io_M_AXI_WDATA, // @[:@141778.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@141778.4]
  output         io_M_AXI_WLAST, // @[:@141778.4]
  output         io_M_AXI_WVALID, // @[:@141778.4]
  input          io_M_AXI_WREADY, // @[:@141778.4]
  output         io_M_AXI_RREADY, // @[:@141778.4]
  input  [31:0]  io_M_AXI_BID, // @[:@141778.4]
  input          io_M_AXI_BVALID, // @[:@141778.4]
  output         io_M_AXI_BREADY // @[:@141778.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@141935.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@141936.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@141937.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@141945.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@141972.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@141977.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@141988.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@141997.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@142006.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@142015.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@142024.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@142033.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@142041.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@141935.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@141936.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@141937.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@141945.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@141972.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@141977.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@141988.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@141997.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@142006.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@142015.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@142024.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@142033.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@142041.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@141949.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@142046.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@142099.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@142101.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@141950.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@141951.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@141955.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@141963.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@141933.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@141934.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@141938.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@141947.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@141979.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@142043.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@142044.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@142045.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@142096.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@142097.4]
endmodule
module FringeZynq( // @[:@143087.2]
  input          clock, // @[:@143088.4]
  input          reset, // @[:@143089.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@143090.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@143090.4]
  input          io_S_AXI_AWVALID, // @[:@143090.4]
  output         io_S_AXI_AWREADY, // @[:@143090.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@143090.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@143090.4]
  input          io_S_AXI_ARVALID, // @[:@143090.4]
  output         io_S_AXI_ARREADY, // @[:@143090.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@143090.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@143090.4]
  input          io_S_AXI_WVALID, // @[:@143090.4]
  output         io_S_AXI_WREADY, // @[:@143090.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@143090.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@143090.4]
  output         io_S_AXI_RVALID, // @[:@143090.4]
  input          io_S_AXI_RREADY, // @[:@143090.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@143090.4]
  output         io_S_AXI_BVALID, // @[:@143090.4]
  input          io_S_AXI_BREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@143090.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@143090.4]
  output         io_M_AXI_0_AWVALID, // @[:@143090.4]
  input          io_M_AXI_0_AWREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@143090.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@143090.4]
  output         io_M_AXI_0_ARVALID, // @[:@143090.4]
  input          io_M_AXI_0_ARREADY, // @[:@143090.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@143090.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@143090.4]
  output         io_M_AXI_0_WLAST, // @[:@143090.4]
  output         io_M_AXI_0_WVALID, // @[:@143090.4]
  input          io_M_AXI_0_WREADY, // @[:@143090.4]
  output         io_M_AXI_0_RREADY, // @[:@143090.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@143090.4]
  input          io_M_AXI_0_BVALID, // @[:@143090.4]
  output         io_M_AXI_0_BREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@143090.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@143090.4]
  output         io_M_AXI_1_AWVALID, // @[:@143090.4]
  input          io_M_AXI_1_AWREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@143090.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@143090.4]
  output         io_M_AXI_1_ARVALID, // @[:@143090.4]
  input          io_M_AXI_1_ARREADY, // @[:@143090.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@143090.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@143090.4]
  output         io_M_AXI_1_WLAST, // @[:@143090.4]
  output         io_M_AXI_1_WVALID, // @[:@143090.4]
  input          io_M_AXI_1_WREADY, // @[:@143090.4]
  output         io_M_AXI_1_RREADY, // @[:@143090.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@143090.4]
  input          io_M_AXI_1_BVALID, // @[:@143090.4]
  output         io_M_AXI_1_BREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@143090.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@143090.4]
  output         io_M_AXI_2_AWVALID, // @[:@143090.4]
  input          io_M_AXI_2_AWREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@143090.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@143090.4]
  output         io_M_AXI_2_ARVALID, // @[:@143090.4]
  input          io_M_AXI_2_ARREADY, // @[:@143090.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@143090.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@143090.4]
  output         io_M_AXI_2_WLAST, // @[:@143090.4]
  output         io_M_AXI_2_WVALID, // @[:@143090.4]
  input          io_M_AXI_2_WREADY, // @[:@143090.4]
  output         io_M_AXI_2_RREADY, // @[:@143090.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@143090.4]
  input          io_M_AXI_2_BVALID, // @[:@143090.4]
  output         io_M_AXI_2_BREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@143090.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@143090.4]
  output         io_M_AXI_3_AWVALID, // @[:@143090.4]
  input          io_M_AXI_3_AWREADY, // @[:@143090.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@143090.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@143090.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@143090.4]
  output         io_M_AXI_3_ARVALID, // @[:@143090.4]
  input          io_M_AXI_3_ARREADY, // @[:@143090.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@143090.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@143090.4]
  output         io_M_AXI_3_WLAST, // @[:@143090.4]
  output         io_M_AXI_3_WVALID, // @[:@143090.4]
  input          io_M_AXI_3_WREADY, // @[:@143090.4]
  output         io_M_AXI_3_RREADY, // @[:@143090.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@143090.4]
  input          io_M_AXI_3_BVALID, // @[:@143090.4]
  output         io_M_AXI_3_BREADY, // @[:@143090.4]
  output         io_enable, // @[:@143090.4]
  input          io_done, // @[:@143090.4]
  output         io_reset, // @[:@143090.4]
  output [63:0]  io_argIns_0, // @[:@143090.4]
  output [63:0]  io_argIns_1, // @[:@143090.4]
  input          io_argOuts_0_valid, // @[:@143090.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@143090.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@143090.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@143090.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@143090.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@143090.4]
  output         io_memStreams_stores_0_data_ready, // @[:@143090.4]
  input          io_memStreams_stores_0_data_valid, // @[:@143090.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@143090.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@143090.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@143090.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@143090.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@143090.4]
  input          io_heap_0_req_valid, // @[:@143090.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@143090.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@143090.4]
  output         io_heap_0_resp_valid, // @[:@143090.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@143090.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@143090.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@143561.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@143561.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@143561.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@144467.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@144467.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@144467.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@144467.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@144467.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@144467.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@144467.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@144467.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@144617.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@144617.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@144617.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@144617.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@144617.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@144617.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@144617.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@144773.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@144773.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@144773.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@144773.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@144773.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@144773.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@144773.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@144929.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@144929.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@144929.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@144929.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@144929.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@144929.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@144929.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145085.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145085.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145085.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145085.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145085.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145085.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145085.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145085.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@143561.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@144467.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@144617.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@144773.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@144929.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@145085.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@144485.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@144481.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@144477.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@144476.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@144475.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@144474.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@144472.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@144471.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@144772.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@144770.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@144769.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@144762.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@144760.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@144758.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@144757.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@144750.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@144748.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@144747.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@144746.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@144745.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@144737.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@144732.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@144928.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@144926.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@144925.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@144918.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@144916.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@144914.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@144913.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@144906.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@144904.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@144903.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@144902.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@144901.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@144893.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@144888.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@145084.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@145082.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@145081.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@145074.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@145072.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@145070.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@145069.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@145062.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@145060.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@145059.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@145058.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@145057.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@145049.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@145044.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@145240.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@145238.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@145237.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@145230.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@145228.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@145226.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@145225.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@145218.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@145216.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@145215.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@145214.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@145213.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@145205.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@145200.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@144495.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@144499.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@144500.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@144501.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@144588.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@144584.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@144579.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@144578.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@144613.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@144612.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@144611.4]
  assign fringeCommon_clock = clock; // @[:@143562.4]
  assign fringeCommon_reset = reset; // @[:@143563.4 FringeZynq.scala 117:22:@144498.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@144489.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@144490.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@144491.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@144492.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@144496.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@144503.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@144502.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@144587.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@144586.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@144585.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@144583.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@144582.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@144581.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@144580.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@144731.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@144724.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@144621.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@144620.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@144887.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@144880.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@144777.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@144776.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@145043.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@145036.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@144933.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@144932.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@145199.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@145192.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145089.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145088.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@144616.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@144615.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@144614.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@144468.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@144469.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@144488.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@144487.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@144486.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@144484.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@144483.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@144482.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@144480.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@144479.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@144478.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@144473.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@144470.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@144493.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@144730.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@144729.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@144728.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@144726.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@144725.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@144723.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@144707.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@144708.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@144709.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@144710.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@144711.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@144712.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@144713.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@144714.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@144715.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@144716.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@144717.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@144718.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@144719.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@144720.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@144721.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@144722.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@144643.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@144644.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@144645.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@144646.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@144647.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@144648.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@144649.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@144650.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@144651.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@144652.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@144653.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@144654.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@144655.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@144656.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@144657.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@144658.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@144659.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@144660.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@144661.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@144662.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@144663.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@144664.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@144665.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@144666.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@144667.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@144668.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@144669.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@144670.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@144671.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@144672.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@144673.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@144674.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@144675.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@144676.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@144677.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@144678.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@144679.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@144680.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@144681.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@144682.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@144683.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@144684.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@144685.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@144686.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@144687.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@144688.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@144689.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@144690.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@144691.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@144692.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@144693.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@144694.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@144695.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@144696.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@144697.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@144698.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@144699.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@144700.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@144701.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@144702.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@144703.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@144704.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@144705.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@144706.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@144642.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@144641.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@144622.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@144761.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@144749.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@144744.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@144736.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@144733.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@144886.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@144885.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@144884.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@144882.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@144881.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@144879.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@144863.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@144864.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@144865.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@144866.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@144867.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@144868.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@144869.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@144870.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@144871.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@144872.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@144873.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@144874.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@144875.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@144876.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@144877.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@144878.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@144799.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@144800.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@144801.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@144802.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@144803.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@144804.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@144805.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@144806.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@144807.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@144808.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@144809.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@144810.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@144811.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@144812.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@144813.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@144814.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@144815.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@144816.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@144817.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@144818.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@144819.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@144820.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@144821.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@144822.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@144823.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@144824.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@144825.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@144826.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@144827.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@144828.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@144829.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@144830.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@144831.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@144832.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@144833.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@144834.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@144835.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@144836.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@144837.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@144838.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@144839.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@144840.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@144841.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@144842.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@144843.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@144844.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@144845.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@144846.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@144847.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@144848.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@144849.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@144850.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@144851.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@144852.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@144853.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@144854.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@144855.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@144856.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@144857.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@144858.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@144859.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@144860.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@144861.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@144862.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@144798.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@144797.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@144778.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@144917.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@144905.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@144900.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@144892.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@144889.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@145042.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@145041.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@145040.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@145038.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@145037.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@145035.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@145019.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@145020.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@145021.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@145022.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@145023.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@145024.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@145025.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@145026.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@145027.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@145028.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@145029.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@145030.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@145031.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@145032.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@145033.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@145034.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@144955.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@144956.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@144957.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@144958.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@144959.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@144960.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@144961.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@144962.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@144963.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@144964.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@144965.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@144966.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@144967.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@144968.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@144969.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@144970.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@144971.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@144972.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@144973.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@144974.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@144975.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@144976.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@144977.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@144978.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@144979.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@144980.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@144981.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@144982.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@144983.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@144984.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@144985.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@144986.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@144987.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@144988.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@144989.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@144990.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@144991.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@144992.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@144993.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@144994.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@144995.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@144996.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@144997.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@144998.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@144999.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@145000.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@145001.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@145002.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@145003.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@145004.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@145005.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@145006.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@145007.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@145008.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@145009.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@145010.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@145011.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@145012.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@145013.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@145014.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@145015.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@145016.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@145017.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@145018.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@144954.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@144953.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@144934.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@145073.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@145061.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@145056.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@145048.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@145045.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@145198.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@145197.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@145196.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@145194.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@145193.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@145191.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@145175.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@145176.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@145177.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@145178.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@145179.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@145180.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@145181.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@145182.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@145183.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@145184.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@145185.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@145186.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@145187.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@145188.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@145189.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@145190.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@145111.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@145112.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@145113.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@145114.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@145115.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@145116.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@145117.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@145118.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@145119.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@145120.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@145121.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@145122.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@145123.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@145124.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@145125.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@145126.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@145127.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@145128.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@145129.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@145130.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@145131.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@145132.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@145133.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@145134.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@145135.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@145136.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@145137.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@145138.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@145139.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@145140.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@145141.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@145142.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@145143.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@145144.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@145145.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@145146.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@145147.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@145148.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@145149.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@145150.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@145151.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@145152.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@145153.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@145154.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@145155.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@145156.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@145157.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@145158.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@145159.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@145160.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@145161.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@145162.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@145163.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@145164.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@145165.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@145166.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@145167.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@145168.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@145169.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@145170.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@145171.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@145172.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@145173.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@145174.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@145110.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@145109.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@145090.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@145229.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@145217.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@145212.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@145204.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@145201.4]
endmodule
module SpatialIP( // @[:@145242.2]
  input          clock, // @[:@145243.4]
  input          reset, // @[:@145244.4]
  input          io_raddr, // @[:@145245.4]
  input          io_wen, // @[:@145245.4]
  input          io_waddr, // @[:@145245.4]
  input          io_wdata, // @[:@145245.4]
  output         io_rdata, // @[:@145245.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@145245.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@145245.4]
  input          io_S_AXI_AWVALID, // @[:@145245.4]
  output         io_S_AXI_AWREADY, // @[:@145245.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@145245.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@145245.4]
  input          io_S_AXI_ARVALID, // @[:@145245.4]
  output         io_S_AXI_ARREADY, // @[:@145245.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@145245.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@145245.4]
  input          io_S_AXI_WVALID, // @[:@145245.4]
  output         io_S_AXI_WREADY, // @[:@145245.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@145245.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@145245.4]
  output         io_S_AXI_RVALID, // @[:@145245.4]
  input          io_S_AXI_RREADY, // @[:@145245.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@145245.4]
  output         io_S_AXI_BVALID, // @[:@145245.4]
  input          io_S_AXI_BREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@145245.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@145245.4]
  output         io_M_AXI_0_AWLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@145245.4]
  output         io_M_AXI_0_AWVALID, // @[:@145245.4]
  input          io_M_AXI_0_AWREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@145245.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@145245.4]
  output         io_M_AXI_0_ARLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@145245.4]
  output         io_M_AXI_0_ARVALID, // @[:@145245.4]
  input          io_M_AXI_0_ARREADY, // @[:@145245.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@145245.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@145245.4]
  output         io_M_AXI_0_WLAST, // @[:@145245.4]
  output         io_M_AXI_0_WVALID, // @[:@145245.4]
  input          io_M_AXI_0_WREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@145245.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@145245.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@145245.4]
  input          io_M_AXI_0_RLAST, // @[:@145245.4]
  input          io_M_AXI_0_RVALID, // @[:@145245.4]
  output         io_M_AXI_0_RREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@145245.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@145245.4]
  input          io_M_AXI_0_BVALID, // @[:@145245.4]
  output         io_M_AXI_0_BREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@145245.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@145245.4]
  output         io_M_AXI_1_AWLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@145245.4]
  output         io_M_AXI_1_AWVALID, // @[:@145245.4]
  input          io_M_AXI_1_AWREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@145245.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@145245.4]
  output         io_M_AXI_1_ARLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@145245.4]
  output         io_M_AXI_1_ARVALID, // @[:@145245.4]
  input          io_M_AXI_1_ARREADY, // @[:@145245.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@145245.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@145245.4]
  output         io_M_AXI_1_WLAST, // @[:@145245.4]
  output         io_M_AXI_1_WVALID, // @[:@145245.4]
  input          io_M_AXI_1_WREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@145245.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@145245.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@145245.4]
  input          io_M_AXI_1_RLAST, // @[:@145245.4]
  input          io_M_AXI_1_RVALID, // @[:@145245.4]
  output         io_M_AXI_1_RREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@145245.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@145245.4]
  input          io_M_AXI_1_BVALID, // @[:@145245.4]
  output         io_M_AXI_1_BREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@145245.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@145245.4]
  output         io_M_AXI_2_AWLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@145245.4]
  output         io_M_AXI_2_AWVALID, // @[:@145245.4]
  input          io_M_AXI_2_AWREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@145245.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@145245.4]
  output         io_M_AXI_2_ARLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@145245.4]
  output         io_M_AXI_2_ARVALID, // @[:@145245.4]
  input          io_M_AXI_2_ARREADY, // @[:@145245.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@145245.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@145245.4]
  output         io_M_AXI_2_WLAST, // @[:@145245.4]
  output         io_M_AXI_2_WVALID, // @[:@145245.4]
  input          io_M_AXI_2_WREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@145245.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@145245.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@145245.4]
  input          io_M_AXI_2_RLAST, // @[:@145245.4]
  input          io_M_AXI_2_RVALID, // @[:@145245.4]
  output         io_M_AXI_2_RREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@145245.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@145245.4]
  input          io_M_AXI_2_BVALID, // @[:@145245.4]
  output         io_M_AXI_2_BREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@145245.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@145245.4]
  output         io_M_AXI_3_AWLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@145245.4]
  output         io_M_AXI_3_AWVALID, // @[:@145245.4]
  input          io_M_AXI_3_AWREADY, // @[:@145245.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@145245.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@145245.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@145245.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@145245.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@145245.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@145245.4]
  output         io_M_AXI_3_ARLOCK, // @[:@145245.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@145245.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@145245.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@145245.4]
  output         io_M_AXI_3_ARVALID, // @[:@145245.4]
  input          io_M_AXI_3_ARREADY, // @[:@145245.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@145245.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@145245.4]
  output         io_M_AXI_3_WLAST, // @[:@145245.4]
  output         io_M_AXI_3_WVALID, // @[:@145245.4]
  input          io_M_AXI_3_WREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@145245.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@145245.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@145245.4]
  input          io_M_AXI_3_RLAST, // @[:@145245.4]
  input          io_M_AXI_3_RVALID, // @[:@145245.4]
  output         io_M_AXI_3_RREADY, // @[:@145245.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@145245.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@145245.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@145245.4]
  input          io_M_AXI_3_BVALID, // @[:@145245.4]
  output         io_M_AXI_3_BREADY, // @[:@145245.4]
  input          io_TOP_AXI_AWID, // @[:@145245.4]
  input          io_TOP_AXI_AWUSER, // @[:@145245.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@145245.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@145245.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@145245.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@145245.4]
  input          io_TOP_AXI_AWLOCK, // @[:@145245.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@145245.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@145245.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@145245.4]
  input          io_TOP_AXI_AWVALID, // @[:@145245.4]
  input          io_TOP_AXI_AWREADY, // @[:@145245.4]
  input          io_TOP_AXI_ARID, // @[:@145245.4]
  input          io_TOP_AXI_ARUSER, // @[:@145245.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@145245.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@145245.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@145245.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@145245.4]
  input          io_TOP_AXI_ARLOCK, // @[:@145245.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@145245.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@145245.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@145245.4]
  input          io_TOP_AXI_ARVALID, // @[:@145245.4]
  input          io_TOP_AXI_ARREADY, // @[:@145245.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@145245.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@145245.4]
  input          io_TOP_AXI_WLAST, // @[:@145245.4]
  input          io_TOP_AXI_WVALID, // @[:@145245.4]
  input          io_TOP_AXI_WREADY, // @[:@145245.4]
  input          io_TOP_AXI_RID, // @[:@145245.4]
  input          io_TOP_AXI_RUSER, // @[:@145245.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@145245.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@145245.4]
  input          io_TOP_AXI_RLAST, // @[:@145245.4]
  input          io_TOP_AXI_RVALID, // @[:@145245.4]
  input          io_TOP_AXI_RREADY, // @[:@145245.4]
  input          io_TOP_AXI_BID, // @[:@145245.4]
  input          io_TOP_AXI_BUSER, // @[:@145245.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@145245.4]
  input          io_TOP_AXI_BVALID, // @[:@145245.4]
  input          io_TOP_AXI_BREADY, // @[:@145245.4]
  input          io_DWIDTH_AXI_AWID, // @[:@145245.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@145245.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@145245.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@145245.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@145245.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@145245.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@145245.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@145245.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@145245.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@145245.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@145245.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@145245.4]
  input          io_DWIDTH_AXI_ARID, // @[:@145245.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@145245.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@145245.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@145245.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@145245.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@145245.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@145245.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@145245.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@145245.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@145245.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@145245.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@145245.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@145245.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@145245.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@145245.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@145245.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@145245.4]
  input          io_DWIDTH_AXI_RID, // @[:@145245.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@145245.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@145245.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@145245.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@145245.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@145245.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@145245.4]
  input          io_DWIDTH_AXI_BID, // @[:@145245.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@145245.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@145245.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@145245.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@145245.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@145245.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@145245.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@145245.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@145245.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@145245.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@145245.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@145245.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@145245.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@145245.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@145245.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@145245.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@145245.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@145245.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@145245.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@145245.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@145245.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@145245.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@145245.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@145245.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@145245.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@145245.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@145245.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@145245.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@145245.4]
  input          io_PROTOCOL_AXI_RID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@145245.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@145245.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@145245.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@145245.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@145245.4]
  input          io_PROTOCOL_AXI_BID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@145245.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@145245.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@145245.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@145245.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@145245.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@145245.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@145245.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@145245.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@145245.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@145245.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@145245.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@145245.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@145245.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@145245.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@145245.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@145245.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@145245.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@145245.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@145245.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@145245.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@145245.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@145245.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@145245.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@145245.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@145247.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@145247.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@145247.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@145247.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@145247.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@145247.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@145247.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@145247.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@145247.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@145247.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@145389.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@145389.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@145389.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@145389.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@145389.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@145389.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@145389.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@145247.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@145389.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@145407.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@145403.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@145399.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@145398.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@145397.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@145396.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@145394.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@145393.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@145451.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@145450.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@145449.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@145448.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@145447.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@145446.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@145445.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@145444.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@145443.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@145442.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@145441.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@145439.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@145438.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@145437.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@145436.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@145435.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@145434.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@145433.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@145432.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@145431.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@145430.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@145429.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@145427.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@145426.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@145425.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@145424.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@145416.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@145411.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@145492.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@145491.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@145490.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@145489.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@145488.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@145487.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@145486.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@145485.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@145484.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@145483.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@145482.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@145480.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@145479.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@145478.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@145477.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@145476.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@145475.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@145474.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@145473.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@145472.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@145471.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@145470.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@145468.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@145467.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@145466.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@145465.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@145457.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@145452.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@145533.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@145532.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@145531.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@145530.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@145529.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@145528.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@145527.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@145526.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@145525.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@145524.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@145523.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@145521.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@145520.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@145519.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@145518.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@145517.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@145516.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@145515.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@145514.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@145513.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@145512.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@145511.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@145509.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@145508.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@145507.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@145506.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@145498.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@145493.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@145574.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@145573.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@145572.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@145571.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@145570.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@145569.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@145568.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@145567.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@145566.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@145565.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@145564.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@145562.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@145561.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@145560.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@145559.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@145558.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@145557.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@145556.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@145555.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@145554.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@145553.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@145552.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@145550.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@145549.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@145548.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@145547.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@145539.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@145534.4]
  assign accel_clock = clock; // @[:@145248.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@145249.4 Zynq.scala 54:17:@145863.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@145858.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@145851.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@145846.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@145830.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@145831.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@145832.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@145833.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@145834.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@145835.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@145836.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@145837.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@145838.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@145839.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@145840.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@145841.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@145842.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@145843.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@145844.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@145845.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@145829.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@145825.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@145820.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@145819.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@145818.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@145799.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@145783.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@145784.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@145785.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@145786.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@145787.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@145788.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@145789.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@145790.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@145791.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@145792.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@145793.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@145794.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@145795.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@145796.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@145797.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@145798.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@145782.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@145747.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@145746.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@145854.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@145853.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@145852.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@145740.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@145741.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@145744.4]
  assign FringeZynq_clock = clock; // @[:@145390.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@145391.4 Zynq.scala 53:18:@145862.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@145410.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@145409.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@145408.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@145406.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@145405.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@145404.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@145402.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@145401.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@145400.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@145395.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@145392.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@145440.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@145428.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@145423.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@145415.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@145412.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@145481.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@145469.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@145464.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@145456.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@145453.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@145522.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@145510.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@145505.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@145497.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@145494.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@145563.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@145551.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@145546.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@145538.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@145535.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@145859.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@145743.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@145742.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@145828.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@145827.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@145826.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@145824.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@145823.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@145822.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@145821.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@145857.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@145856.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@145855.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




