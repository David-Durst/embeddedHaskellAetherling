module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module atomTupleCreator_t0Int_t1Int (input [7:0] I0/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O__0/*verilator public*/, output [7:0] O__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O__0 = I0;
assign O__1 = I1;
assign valid_down = valid_up;
endmodule

module coreir_term #(parameter width = 1) (input [width-1:0] in/*verilator public*/);

endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out/*verilator public*/);
  assign out = value;
endmodule

module coreir_add #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 + in1;
endmodule

module lutN #(parameter N = 1, parameter init = 1) (input [N-1:0] in/*verilator public*/, output out/*verilator public*/);
  assign out = init[in];
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit840 (input [319:0] in/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/, output [7:0] out_10/*verilator public*/, output [7:0] out_11/*verilator public*/, output [7:0] out_12/*verilator public*/, output [7:0] out_13/*verilator public*/, output [7:0] out_14/*verilator public*/, output [7:0] out_15/*verilator public*/, output [7:0] out_16/*verilator public*/, output [7:0] out_17/*verilator public*/, output [7:0] out_18/*verilator public*/, output [7:0] out_19/*verilator public*/, output [7:0] out_2/*verilator public*/, output [7:0] out_20/*verilator public*/, output [7:0] out_21/*verilator public*/, output [7:0] out_22/*verilator public*/, output [7:0] out_23/*verilator public*/, output [7:0] out_24/*verilator public*/, output [7:0] out_25/*verilator public*/, output [7:0] out_26/*verilator public*/, output [7:0] out_27/*verilator public*/, output [7:0] out_28/*verilator public*/, output [7:0] out_29/*verilator public*/, output [7:0] out_3/*verilator public*/, output [7:0] out_30/*verilator public*/, output [7:0] out_31/*verilator public*/, output [7:0] out_32/*verilator public*/, output [7:0] out_33/*verilator public*/, output [7:0] out_34/*verilator public*/, output [7:0] out_35/*verilator public*/, output [7:0] out_36/*verilator public*/, output [7:0] out_37/*verilator public*/, output [7:0] out_38/*verilator public*/, output [7:0] out_39/*verilator public*/, output [7:0] out_4/*verilator public*/, output [7:0] out_5/*verilator public*/, output [7:0] out_6/*verilator public*/, output [7:0] out_7/*verilator public*/, output [7:0] out_8/*verilator public*/, output [7:0] out_9/*verilator public*/);
assign out_0 = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
assign out_1 = {in[15],in[14],in[13],in[12],in[11],in[10],in[9],in[8]};
assign out_10 = {in[87],in[86],in[85],in[84],in[83],in[82],in[81],in[80]};
assign out_11 = {in[95],in[94],in[93],in[92],in[91],in[90],in[89],in[88]};
assign out_12 = {in[103],in[102],in[101],in[100],in[99],in[98],in[97],in[96]};
assign out_13 = {in[111],in[110],in[109],in[108],in[107],in[106],in[105],in[104]};
assign out_14 = {in[119],in[118],in[117],in[116],in[115],in[114],in[113],in[112]};
assign out_15 = {in[127],in[126],in[125],in[124],in[123],in[122],in[121],in[120]};
assign out_16 = {in[135],in[134],in[133],in[132],in[131],in[130],in[129],in[128]};
assign out_17 = {in[143],in[142],in[141],in[140],in[139],in[138],in[137],in[136]};
assign out_18 = {in[151],in[150],in[149],in[148],in[147],in[146],in[145],in[144]};
assign out_19 = {in[159],in[158],in[157],in[156],in[155],in[154],in[153],in[152]};
assign out_2 = {in[23],in[22],in[21],in[20],in[19],in[18],in[17],in[16]};
assign out_20 = {in[167],in[166],in[165],in[164],in[163],in[162],in[161],in[160]};
assign out_21 = {in[175],in[174],in[173],in[172],in[171],in[170],in[169],in[168]};
assign out_22 = {in[183],in[182],in[181],in[180],in[179],in[178],in[177],in[176]};
assign out_23 = {in[191],in[190],in[189],in[188],in[187],in[186],in[185],in[184]};
assign out_24 = {in[199],in[198],in[197],in[196],in[195],in[194],in[193],in[192]};
assign out_25 = {in[207],in[206],in[205],in[204],in[203],in[202],in[201],in[200]};
assign out_26 = {in[215],in[214],in[213],in[212],in[211],in[210],in[209],in[208]};
assign out_27 = {in[223],in[222],in[221],in[220],in[219],in[218],in[217],in[216]};
assign out_28 = {in[231],in[230],in[229],in[228],in[227],in[226],in[225],in[224]};
assign out_29 = {in[239],in[238],in[237],in[236],in[235],in[234],in[233],in[232]};
assign out_3 = {in[31],in[30],in[29],in[28],in[27],in[26],in[25],in[24]};
assign out_30 = {in[247],in[246],in[245],in[244],in[243],in[242],in[241],in[240]};
assign out_31 = {in[255],in[254],in[253],in[252],in[251],in[250],in[249],in[248]};
assign out_32 = {in[263],in[262],in[261],in[260],in[259],in[258],in[257],in[256]};
assign out_33 = {in[271],in[270],in[269],in[268],in[267],in[266],in[265],in[264]};
assign out_34 = {in[279],in[278],in[277],in[276],in[275],in[274],in[273],in[272]};
assign out_35 = {in[287],in[286],in[285],in[284],in[283],in[282],in[281],in[280]};
assign out_36 = {in[295],in[294],in[293],in[292],in[291],in[290],in[289],in[288]};
assign out_37 = {in[303],in[302],in[301],in[300],in[299],in[298],in[297],in[296]};
assign out_38 = {in[311],in[310],in[309],in[308],in[307],in[306],in[305],in[304]};
assign out_39 = {in[319],in[318],in[317],in[316],in[315],in[314],in[313],in[312]};
assign out_4 = {in[39],in[38],in[37],in[36],in[35],in[34],in[33],in[32]};
assign out_5 = {in[47],in[46],in[45],in[44],in[43],in[42],in[41],in[40]};
assign out_6 = {in[55],in[54],in[53],in[52],in[51],in[50],in[49],in[48]};
assign out_7 = {in[63],in[62],in[61],in[60],in[59],in[58],in[57],in[56]};
assign out_8 = {in[71],in[70],in[69],in[68],in[67],in[66],in[65],in[64]};
assign out_9 = {in[79],in[78],in[77],in[76],in[75],in[74],in[73],in[72]};
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit8 (input [7:0] in/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit (input [0:0] in/*verilator public*/, output out/*verilator public*/);
assign out = in[0];
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit840 (input [7:0] in_0/*verilator public*/, input [7:0] in_1/*verilator public*/, input [7:0] in_10/*verilator public*/, input [7:0] in_11/*verilator public*/, input [7:0] in_12/*verilator public*/, input [7:0] in_13/*verilator public*/, input [7:0] in_14/*verilator public*/, input [7:0] in_15/*verilator public*/, input [7:0] in_16/*verilator public*/, input [7:0] in_17/*verilator public*/, input [7:0] in_18/*verilator public*/, input [7:0] in_19/*verilator public*/, input [7:0] in_2/*verilator public*/, input [7:0] in_20/*verilator public*/, input [7:0] in_21/*verilator public*/, input [7:0] in_22/*verilator public*/, input [7:0] in_23/*verilator public*/, input [7:0] in_24/*verilator public*/, input [7:0] in_25/*verilator public*/, input [7:0] in_26/*verilator public*/, input [7:0] in_27/*verilator public*/, input [7:0] in_28/*verilator public*/, input [7:0] in_29/*verilator public*/, input [7:0] in_3/*verilator public*/, input [7:0] in_30/*verilator public*/, input [7:0] in_31/*verilator public*/, input [7:0] in_32/*verilator public*/, input [7:0] in_33/*verilator public*/, input [7:0] in_34/*verilator public*/, input [7:0] in_35/*verilator public*/, input [7:0] in_36/*verilator public*/, input [7:0] in_37/*verilator public*/, input [7:0] in_38/*verilator public*/, input [7:0] in_39/*verilator public*/, input [7:0] in_4/*verilator public*/, input [7:0] in_5/*verilator public*/, input [7:0] in_6/*verilator public*/, input [7:0] in_7/*verilator public*/, input [7:0] in_8/*verilator public*/, input [7:0] in_9/*verilator public*/, output [319:0] out/*verilator public*/);
assign out = {in_39[7],in_39[6],in_39[5],in_39[4],in_39[3],in_39[2],in_39[1],in_39[0],in_38[7],in_38[6],in_38[5],in_38[4],in_38[3],in_38[2],in_38[1],in_38[0],in_37[7],in_37[6],in_37[5],in_37[4],in_37[3],in_37[2],in_37[1],in_37[0],in_36[7],in_36[6],in_36[5],in_36[4],in_36[3],in_36[2],in_36[1],in_36[0],in_35[7],in_35[6],in_35[5],in_35[4],in_35[3],in_35[2],in_35[1],in_35[0],in_34[7],in_34[6],in_34[5],in_34[4],in_34[3],in_34[2],in_34[1],in_34[0],in_33[7],in_33[6],in_33[5],in_33[4],in_33[3],in_33[2],in_33[1],in_33[0],in_32[7],in_32[6],in_32[5],in_32[4],in_32[3],in_32[2],in_32[1],in_32[0],in_31[7],in_31[6],in_31[5],in_31[4],in_31[3],in_31[2],in_31[1],in_31[0],in_30[7],in_30[6],in_30[5],in_30[4],in_30[3],in_30[2],in_30[1],in_30[0],in_29[7],in_29[6],in_29[5],in_29[4],in_29[3],in_29[2],in_29[1],in_29[0],in_28[7],in_28[6],in_28[5],in_28[4],in_28[3],in_28[2],in_28[1],in_28[0],in_27[7],in_27[6],in_27[5],in_27[4],in_27[3],in_27[2],in_27[1],in_27[0],in_26[7],in_26[6],in_26[5],in_26[4],in_26[3],in_26[2],in_26[1],in_26[0],in_25[7],in_25[6],in_25[5],in_25[4],in_25[3],in_25[2],in_25[1],in_25[0],in_24[7],in_24[6],in_24[5],in_24[4],in_24[3],in_24[2],in_24[1],in_24[0],in_23[7],in_23[6],in_23[5],in_23[4],in_23[3],in_23[2],in_23[1],in_23[0],in_22[7],in_22[6],in_22[5],in_22[4],in_22[3],in_22[2],in_22[1],in_22[0],in_21[7],in_21[6],in_21[5],in_21[4],in_21[3],in_21[2],in_21[1],in_21[0],in_20[7],in_20[6],in_20[5],in_20[4],in_20[3],in_20[2],in_20[1],in_20[0],in_19[7],in_19[6],in_19[5],in_19[4],in_19[3],in_19[2],in_19[1],in_19[0],in_18[7],in_18[6],in_18[5],in_18[4],in_18[3],in_18[2],in_18[1],in_18[0],in_17[7],in_17[6],in_17[5],in_17[4],in_17[3],in_17[2],in_17[1],in_17[0],in_16[7],in_16[6],in_16[5],in_16[4],in_16[3],in_16[2],in_16[1],in_16[0],in_15[7],in_15[6],in_15[5],in_15[4],in_15[3],in_15[2],in_15[1],in_15[0],in_14[7],in_14[6],in_14[5],in_14[4],in_14[3],in_14[2],in_14[1],in_14[0],in_13[7],in_13[6],in_13[5],in_13[4],in_13[3],in_13[2],in_13[1],in_13[0],in_12[7],in_12[6],in_12[5],in_12[4],in_12[3],in_12[2],in_12[1],in_12[0],in_11[7],in_11[6],in_11[5],in_11[4],in_11[3],in_11[2],in_11[1],in_11[0],in_10[7],in_10[6],in_10[5],in_10[4],in_10[3],in_10[2],in_10[1],in_10[0],in_9[7],in_9[6],in_9[5],in_9[4],in_9[3],in_9[2],in_9[1],in_9[0],in_8[7],in_8[6],in_8[5],in_8[4],in_8[3],in_8[2],in_8[1],in_8[0],in_7[7],in_7[6],in_7[5],in_7[4],in_7[3],in_7[2],in_7[1],in_7[0],in_6[7],in_6[6],in_6[5],in_6[4],in_6[3],in_6[2],in_6[1],in_6[0],in_5[7],in_5[6],in_5[5],in_5[4],in_5[3],in_5[2],in_5[1],in_5[0],in_4[7],in_4[6],in_4[5],in_4[4],in_4[3],in_4[2],in_4[1],in_4[0],in_3[7],in_3[6],in_3[5],in_3[4],in_3[3],in_3[2],in_3[1],in_3[0],in_2[7],in_2[6],in_2[5],in_2[4],in_2[3],in_2[2],in_2[1],in_2[0],in_1[7],in_1[6],in_1[5],in_1[4],in_1[3],in_1[2],in_1[1],in_1[0],in_0[7],in_0[6],in_0[5],in_0[4],in_0[3],in_0[2],in_0[1],in_0[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit8 (input [7:0] in/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit (input in/*verilator public*/, output [0:0] out/*verilator public*/);
assign out = in;
endmodule

module Term_Bitt (input I/*verilator public*/);
wire [0:0] dehydrate_tBit_inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBit_inst0_out));
endmodule

module SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] const_0_1_out;
Term_Bitt Term_Bitt_inst0(.I(CE));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
assign O = const_0_1_out;
endmodule

module LUT1_1 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h1), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_0 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h0), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT_Array_8_Bit_t_1n (input CLK/*verilator public*/, input [0:0] addr/*verilator public*/, output [7:0] data/*verilator public*/);
wire LUT1_0_inst0_O;
wire LUT1_0_inst1_O;
wire LUT1_0_inst2_O;
wire LUT1_0_inst3_O;
wire LUT1_0_inst4_O;
wire LUT1_0_inst5_O;
wire LUT1_1_inst0_O;
wire LUT1_1_inst1_O;
wire [7:0] hydrate_tArray_8_Bit__inst0_out;
LUT1_0 LUT1_0_inst0(.I0(addr[0]), .O(LUT1_0_inst0_O));
LUT1_0 LUT1_0_inst1(.I0(addr[0]), .O(LUT1_0_inst1_O));
LUT1_0 LUT1_0_inst2(.I0(addr[0]), .O(LUT1_0_inst2_O));
LUT1_0 LUT1_0_inst3(.I0(addr[0]), .O(LUT1_0_inst3_O));
LUT1_0 LUT1_0_inst4(.I0(addr[0]), .O(LUT1_0_inst4_O));
LUT1_0 LUT1_0_inst5(.I0(addr[0]), .O(LUT1_0_inst5_O));
LUT1_1 LUT1_1_inst0(.I0(addr[0]), .O(LUT1_1_inst0_O));
LUT1_1 LUT1_1_inst1(.I0(addr[0]), .O(LUT1_1_inst1_O));
\aetherlinglib_hydrate__hydratedTypeBit8 hydrate_tArray_8_Bit__inst0(.in({LUT1_0_inst5_O,LUT1_0_inst4_O,LUT1_0_inst3_O,LUT1_0_inst2_O,LUT1_0_inst1_O,LUT1_1_inst1_O,LUT1_0_inst0_O,LUT1_1_inst0_O}), .out(hydrate_tArray_8_Bit__inst0_out));
assign data = hydrate_tArray_8_Bit__inst0_out;
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Bit_t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8_inst0_O;
wire [7:0] dehydrate_tArray_8_Bit__inst0_out;
wire [7:0] hydrate_tArray_8_Bit__inst0_out;
Register8 Register8_inst0(.CLK(CLK), .I(dehydrate_tArray_8_Bit__inst0_out), .O(Register8_inst0_O));
\aetherlinglib_dehydrate__hydratedTypeBit8 dehydrate_tArray_8_Bit__inst0(.in(I), .out(dehydrate_tArray_8_Bit__inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit8 hydrate_tArray_8_Bit__inst0(.in(Register8_inst0_O), .out(hydrate_tArray_8_Bit__inst0_out));
assign O = hydrate_tArray_8_Bit__inst0_out;
endmodule

module Register320 (input CLK/*verilator public*/, input [319:0] I/*verilator public*/, output [319:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10(.CLK(CLK), .I(I[10]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100(.CLK(CLK), .I(I[100]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101(.CLK(CLK), .I(I[101]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102(.CLK(CLK), .I(I[102]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103(.CLK(CLK), .I(I[103]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104(.CLK(CLK), .I(I[104]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105(.CLK(CLK), .I(I[105]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106(.CLK(CLK), .I(I[106]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107(.CLK(CLK), .I(I[107]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108(.CLK(CLK), .I(I[108]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109(.CLK(CLK), .I(I[109]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11(.CLK(CLK), .I(I[11]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110(.CLK(CLK), .I(I[110]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111(.CLK(CLK), .I(I[111]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112(.CLK(CLK), .I(I[112]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113(.CLK(CLK), .I(I[113]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114(.CLK(CLK), .I(I[114]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115(.CLK(CLK), .I(I[115]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116(.CLK(CLK), .I(I[116]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117(.CLK(CLK), .I(I[117]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118(.CLK(CLK), .I(I[118]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119(.CLK(CLK), .I(I[119]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12(.CLK(CLK), .I(I[12]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120(.CLK(CLK), .I(I[120]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121(.CLK(CLK), .I(I[121]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122(.CLK(CLK), .I(I[122]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123(.CLK(CLK), .I(I[123]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124(.CLK(CLK), .I(I[124]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125(.CLK(CLK), .I(I[125]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126(.CLK(CLK), .I(I[126]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127(.CLK(CLK), .I(I[127]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128(.CLK(CLK), .I(I[128]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129(.CLK(CLK), .I(I[129]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13(.CLK(CLK), .I(I[13]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130(.CLK(CLK), .I(I[130]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131(.CLK(CLK), .I(I[131]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132(.CLK(CLK), .I(I[132]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133(.CLK(CLK), .I(I[133]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134(.CLK(CLK), .I(I[134]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135(.CLK(CLK), .I(I[135]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136(.CLK(CLK), .I(I[136]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137(.CLK(CLK), .I(I[137]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138(.CLK(CLK), .I(I[138]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139(.CLK(CLK), .I(I[139]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14(.CLK(CLK), .I(I[14]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140(.CLK(CLK), .I(I[140]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141(.CLK(CLK), .I(I[141]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142(.CLK(CLK), .I(I[142]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143(.CLK(CLK), .I(I[143]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144(.CLK(CLK), .I(I[144]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145(.CLK(CLK), .I(I[145]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146(.CLK(CLK), .I(I[146]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147(.CLK(CLK), .I(I[147]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148(.CLK(CLK), .I(I[148]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149(.CLK(CLK), .I(I[149]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15(.CLK(CLK), .I(I[15]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150(.CLK(CLK), .I(I[150]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151(.CLK(CLK), .I(I[151]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152(.CLK(CLK), .I(I[152]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153(.CLK(CLK), .I(I[153]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154(.CLK(CLK), .I(I[154]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155(.CLK(CLK), .I(I[155]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156(.CLK(CLK), .I(I[156]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157(.CLK(CLK), .I(I[157]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158(.CLK(CLK), .I(I[158]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159(.CLK(CLK), .I(I[159]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16(.CLK(CLK), .I(I[16]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160(.CLK(CLK), .I(I[160]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161(.CLK(CLK), .I(I[161]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162(.CLK(CLK), .I(I[162]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163(.CLK(CLK), .I(I[163]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164(.CLK(CLK), .I(I[164]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165(.CLK(CLK), .I(I[165]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166(.CLK(CLK), .I(I[166]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167(.CLK(CLK), .I(I[167]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168(.CLK(CLK), .I(I[168]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169(.CLK(CLK), .I(I[169]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17(.CLK(CLK), .I(I[17]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170(.CLK(CLK), .I(I[170]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171(.CLK(CLK), .I(I[171]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172(.CLK(CLK), .I(I[172]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173(.CLK(CLK), .I(I[173]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174(.CLK(CLK), .I(I[174]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175(.CLK(CLK), .I(I[175]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176(.CLK(CLK), .I(I[176]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177(.CLK(CLK), .I(I[177]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178(.CLK(CLK), .I(I[178]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179(.CLK(CLK), .I(I[179]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18(.CLK(CLK), .I(I[18]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180(.CLK(CLK), .I(I[180]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181(.CLK(CLK), .I(I[181]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182(.CLK(CLK), .I(I[182]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183(.CLK(CLK), .I(I[183]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184(.CLK(CLK), .I(I[184]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185(.CLK(CLK), .I(I[185]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186(.CLK(CLK), .I(I[186]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187(.CLK(CLK), .I(I[187]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188(.CLK(CLK), .I(I[188]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189(.CLK(CLK), .I(I[189]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19(.CLK(CLK), .I(I[19]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190(.CLK(CLK), .I(I[190]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191(.CLK(CLK), .I(I[191]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192(.CLK(CLK), .I(I[192]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193(.CLK(CLK), .I(I[193]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194(.CLK(CLK), .I(I[194]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195(.CLK(CLK), .I(I[195]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196(.CLK(CLK), .I(I[196]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197(.CLK(CLK), .I(I[197]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198(.CLK(CLK), .I(I[198]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199(.CLK(CLK), .I(I[199]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20(.CLK(CLK), .I(I[20]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200(.CLK(CLK), .I(I[200]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201(.CLK(CLK), .I(I[201]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202(.CLK(CLK), .I(I[202]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203(.CLK(CLK), .I(I[203]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204(.CLK(CLK), .I(I[204]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205(.CLK(CLK), .I(I[205]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206(.CLK(CLK), .I(I[206]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207(.CLK(CLK), .I(I[207]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208(.CLK(CLK), .I(I[208]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209(.CLK(CLK), .I(I[209]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21(.CLK(CLK), .I(I[21]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210(.CLK(CLK), .I(I[210]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211(.CLK(CLK), .I(I[211]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212(.CLK(CLK), .I(I[212]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213(.CLK(CLK), .I(I[213]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214(.CLK(CLK), .I(I[214]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215(.CLK(CLK), .I(I[215]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216(.CLK(CLK), .I(I[216]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217(.CLK(CLK), .I(I[217]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218(.CLK(CLK), .I(I[218]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219(.CLK(CLK), .I(I[219]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22(.CLK(CLK), .I(I[22]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220(.CLK(CLK), .I(I[220]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221(.CLK(CLK), .I(I[221]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222(.CLK(CLK), .I(I[222]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223(.CLK(CLK), .I(I[223]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224(.CLK(CLK), .I(I[224]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225(.CLK(CLK), .I(I[225]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226(.CLK(CLK), .I(I[226]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227(.CLK(CLK), .I(I[227]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228(.CLK(CLK), .I(I[228]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229(.CLK(CLK), .I(I[229]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23(.CLK(CLK), .I(I[23]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230(.CLK(CLK), .I(I[230]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231(.CLK(CLK), .I(I[231]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232(.CLK(CLK), .I(I[232]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233(.CLK(CLK), .I(I[233]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234(.CLK(CLK), .I(I[234]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235(.CLK(CLK), .I(I[235]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236(.CLK(CLK), .I(I[236]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237(.CLK(CLK), .I(I[237]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238(.CLK(CLK), .I(I[238]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239(.CLK(CLK), .I(I[239]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24(.CLK(CLK), .I(I[24]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240(.CLK(CLK), .I(I[240]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241(.CLK(CLK), .I(I[241]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242(.CLK(CLK), .I(I[242]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243(.CLK(CLK), .I(I[243]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244(.CLK(CLK), .I(I[244]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245(.CLK(CLK), .I(I[245]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246(.CLK(CLK), .I(I[246]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247(.CLK(CLK), .I(I[247]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248(.CLK(CLK), .I(I[248]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249(.CLK(CLK), .I(I[249]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25(.CLK(CLK), .I(I[25]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250(.CLK(CLK), .I(I[250]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251(.CLK(CLK), .I(I[251]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252(.CLK(CLK), .I(I[252]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253(.CLK(CLK), .I(I[253]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254(.CLK(CLK), .I(I[254]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255(.CLK(CLK), .I(I[255]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256(.CLK(CLK), .I(I[256]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257(.CLK(CLK), .I(I[257]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258(.CLK(CLK), .I(I[258]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259(.CLK(CLK), .I(I[259]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26(.CLK(CLK), .I(I[26]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260(.CLK(CLK), .I(I[260]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261(.CLK(CLK), .I(I[261]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262(.CLK(CLK), .I(I[262]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263(.CLK(CLK), .I(I[263]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264(.CLK(CLK), .I(I[264]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265(.CLK(CLK), .I(I[265]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266(.CLK(CLK), .I(I[266]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267(.CLK(CLK), .I(I[267]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268(.CLK(CLK), .I(I[268]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269(.CLK(CLK), .I(I[269]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27(.CLK(CLK), .I(I[27]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270(.CLK(CLK), .I(I[270]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271(.CLK(CLK), .I(I[271]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272(.CLK(CLK), .I(I[272]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273(.CLK(CLK), .I(I[273]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274(.CLK(CLK), .I(I[274]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275(.CLK(CLK), .I(I[275]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276(.CLK(CLK), .I(I[276]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277(.CLK(CLK), .I(I[277]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278(.CLK(CLK), .I(I[278]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279(.CLK(CLK), .I(I[279]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28(.CLK(CLK), .I(I[28]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280(.CLK(CLK), .I(I[280]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281(.CLK(CLK), .I(I[281]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282(.CLK(CLK), .I(I[282]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283(.CLK(CLK), .I(I[283]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284(.CLK(CLK), .I(I[284]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285(.CLK(CLK), .I(I[285]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286(.CLK(CLK), .I(I[286]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287(.CLK(CLK), .I(I[287]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288(.CLK(CLK), .I(I[288]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289(.CLK(CLK), .I(I[289]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29(.CLK(CLK), .I(I[29]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290(.CLK(CLK), .I(I[290]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291(.CLK(CLK), .I(I[291]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292(.CLK(CLK), .I(I[292]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293(.CLK(CLK), .I(I[293]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294(.CLK(CLK), .I(I[294]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295(.CLK(CLK), .I(I[295]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296(.CLK(CLK), .I(I[296]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297(.CLK(CLK), .I(I[297]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298(.CLK(CLK), .I(I[298]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299(.CLK(CLK), .I(I[299]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30(.CLK(CLK), .I(I[30]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300(.CLK(CLK), .I(I[300]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301(.CLK(CLK), .I(I[301]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302(.CLK(CLK), .I(I[302]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303(.CLK(CLK), .I(I[303]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304(.CLK(CLK), .I(I[304]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305(.CLK(CLK), .I(I[305]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306(.CLK(CLK), .I(I[306]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307(.CLK(CLK), .I(I[307]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308(.CLK(CLK), .I(I[308]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309(.CLK(CLK), .I(I[309]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31(.CLK(CLK), .I(I[31]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310(.CLK(CLK), .I(I[310]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311(.CLK(CLK), .I(I[311]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312(.CLK(CLK), .I(I[312]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313(.CLK(CLK), .I(I[313]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314(.CLK(CLK), .I(I[314]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315(.CLK(CLK), .I(I[315]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316(.CLK(CLK), .I(I[316]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317(.CLK(CLK), .I(I[317]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318(.CLK(CLK), .I(I[318]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319(.CLK(CLK), .I(I[319]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32(.CLK(CLK), .I(I[32]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33(.CLK(CLK), .I(I[33]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34(.CLK(CLK), .I(I[34]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35(.CLK(CLK), .I(I[35]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36(.CLK(CLK), .I(I[36]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37(.CLK(CLK), .I(I[37]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38(.CLK(CLK), .I(I[38]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39(.CLK(CLK), .I(I[39]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40(.CLK(CLK), .I(I[40]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41(.CLK(CLK), .I(I[41]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42(.CLK(CLK), .I(I[42]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43(.CLK(CLK), .I(I[43]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44(.CLK(CLK), .I(I[44]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45(.CLK(CLK), .I(I[45]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46(.CLK(CLK), .I(I[46]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47(.CLK(CLK), .I(I[47]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48(.CLK(CLK), .I(I[48]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49(.CLK(CLK), .I(I[49]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50(.CLK(CLK), .I(I[50]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51(.CLK(CLK), .I(I[51]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52(.CLK(CLK), .I(I[52]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53(.CLK(CLK), .I(I[53]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54(.CLK(CLK), .I(I[54]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55(.CLK(CLK), .I(I[55]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56(.CLK(CLK), .I(I[56]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57(.CLK(CLK), .I(I[57]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58(.CLK(CLK), .I(I[58]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59(.CLK(CLK), .I(I[59]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60(.CLK(CLK), .I(I[60]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61(.CLK(CLK), .I(I[61]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62(.CLK(CLK), .I(I[62]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63(.CLK(CLK), .I(I[63]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64(.CLK(CLK), .I(I[64]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65(.CLK(CLK), .I(I[65]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66(.CLK(CLK), .I(I[66]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67(.CLK(CLK), .I(I[67]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68(.CLK(CLK), .I(I[68]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69(.CLK(CLK), .I(I[69]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70(.CLK(CLK), .I(I[70]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71(.CLK(CLK), .I(I[71]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72(.CLK(CLK), .I(I[72]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73(.CLK(CLK), .I(I[73]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74(.CLK(CLK), .I(I[74]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75(.CLK(CLK), .I(I[75]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76(.CLK(CLK), .I(I[76]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77(.CLK(CLK), .I(I[77]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78(.CLK(CLK), .I(I[78]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79(.CLK(CLK), .I(I[79]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8(.CLK(CLK), .I(I[8]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80(.CLK(CLK), .I(I[80]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81(.CLK(CLK), .I(I[81]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82(.CLK(CLK), .I(I[82]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83(.CLK(CLK), .I(I[83]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84(.CLK(CLK), .I(I[84]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85(.CLK(CLK), .I(I[85]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86(.CLK(CLK), .I(I[86]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87(.CLK(CLK), .I(I[87]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88(.CLK(CLK), .I(I[88]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89(.CLK(CLK), .I(I[89]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9(.CLK(CLK), .I(I[9]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90(.CLK(CLK), .I(I[90]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91(.CLK(CLK), .I(I[91]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92(.CLK(CLK), .I(I[92]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93(.CLK(CLK), .I(I[93]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94(.CLK(CLK), .I(I[94]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95(.CLK(CLK), .I(I[95]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96(.CLK(CLK), .I(I[96]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97(.CLK(CLK), .I(I[97]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98(.CLK(CLK), .I(I[98]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99(.CLK(CLK), .I(I[99]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/);
wire [319:0] Register320_inst0_O;
wire [319:0] dehydrate_tArray_40_Array_8_Bit___inst0_out;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_0;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_1;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_10;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_11;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_12;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_13;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_14;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_15;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_16;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_17;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_18;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_19;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_2;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_20;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_21;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_22;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_23;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_24;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_25;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_26;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_27;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_28;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_29;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_3;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_30;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_31;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_32;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_33;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_34;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_35;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_36;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_37;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_38;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_39;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_4;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_5;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_6;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_7;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_8;
wire [7:0] hydrate_tArray_40_Array_8_Bit___inst0_out_9;
Register320 Register320_inst0(.CLK(CLK), .I(dehydrate_tArray_40_Array_8_Bit___inst0_out), .O(Register320_inst0_O));
\aetherlinglib_dehydrate__hydratedTypeBit840 dehydrate_tArray_40_Array_8_Bit___inst0(.in_0(I_0), .in_1(I_1), .in_10(I_10), .in_11(I_11), .in_12(I_12), .in_13(I_13), .in_14(I_14), .in_15(I_15), .in_16(I_16), .in_17(I_17), .in_18(I_18), .in_19(I_19), .in_2(I_2), .in_20(I_20), .in_21(I_21), .in_22(I_22), .in_23(I_23), .in_24(I_24), .in_25(I_25), .in_26(I_26), .in_27(I_27), .in_28(I_28), .in_29(I_29), .in_3(I_3), .in_30(I_30), .in_31(I_31), .in_32(I_32), .in_33(I_33), .in_34(I_34), .in_35(I_35), .in_36(I_36), .in_37(I_37), .in_38(I_38), .in_39(I_39), .in_4(I_4), .in_5(I_5), .in_6(I_6), .in_7(I_7), .in_8(I_8), .in_9(I_9), .out(dehydrate_tArray_40_Array_8_Bit___inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit840 hydrate_tArray_40_Array_8_Bit___inst0(.in(Register320_inst0_O), .out_0(hydrate_tArray_40_Array_8_Bit___inst0_out_0), .out_1(hydrate_tArray_40_Array_8_Bit___inst0_out_1), .out_10(hydrate_tArray_40_Array_8_Bit___inst0_out_10), .out_11(hydrate_tArray_40_Array_8_Bit___inst0_out_11), .out_12(hydrate_tArray_40_Array_8_Bit___inst0_out_12), .out_13(hydrate_tArray_40_Array_8_Bit___inst0_out_13), .out_14(hydrate_tArray_40_Array_8_Bit___inst0_out_14), .out_15(hydrate_tArray_40_Array_8_Bit___inst0_out_15), .out_16(hydrate_tArray_40_Array_8_Bit___inst0_out_16), .out_17(hydrate_tArray_40_Array_8_Bit___inst0_out_17), .out_18(hydrate_tArray_40_Array_8_Bit___inst0_out_18), .out_19(hydrate_tArray_40_Array_8_Bit___inst0_out_19), .out_2(hydrate_tArray_40_Array_8_Bit___inst0_out_2), .out_20(hydrate_tArray_40_Array_8_Bit___inst0_out_20), .out_21(hydrate_tArray_40_Array_8_Bit___inst0_out_21), .out_22(hydrate_tArray_40_Array_8_Bit___inst0_out_22), .out_23(hydrate_tArray_40_Array_8_Bit___inst0_out_23), .out_24(hydrate_tArray_40_Array_8_Bit___inst0_out_24), .out_25(hydrate_tArray_40_Array_8_Bit___inst0_out_25), .out_26(hydrate_tArray_40_Array_8_Bit___inst0_out_26), .out_27(hydrate_tArray_40_Array_8_Bit___inst0_out_27), .out_28(hydrate_tArray_40_Array_8_Bit___inst0_out_28), .out_29(hydrate_tArray_40_Array_8_Bit___inst0_out_29), .out_3(hydrate_tArray_40_Array_8_Bit___inst0_out_3), .out_30(hydrate_tArray_40_Array_8_Bit___inst0_out_30), .out_31(hydrate_tArray_40_Array_8_Bit___inst0_out_31), .out_32(hydrate_tArray_40_Array_8_Bit___inst0_out_32), .out_33(hydrate_tArray_40_Array_8_Bit___inst0_out_33), .out_34(hydrate_tArray_40_Array_8_Bit___inst0_out_34), .out_35(hydrate_tArray_40_Array_8_Bit___inst0_out_35), .out_36(hydrate_tArray_40_Array_8_Bit___inst0_out_36), .out_37(hydrate_tArray_40_Array_8_Bit___inst0_out_37), .out_38(hydrate_tArray_40_Array_8_Bit___inst0_out_38), .out_39(hydrate_tArray_40_Array_8_Bit___inst0_out_39), .out_4(hydrate_tArray_40_Array_8_Bit___inst0_out_4), .out_5(hydrate_tArray_40_Array_8_Bit___inst0_out_5), .out_6(hydrate_tArray_40_Array_8_Bit___inst0_out_6), .out_7(hydrate_tArray_40_Array_8_Bit___inst0_out_7), .out_8(hydrate_tArray_40_Array_8_Bit___inst0_out_8), .out_9(hydrate_tArray_40_Array_8_Bit___inst0_out_9));
assign O_0 = hydrate_tArray_40_Array_8_Bit___inst0_out_0;
assign O_1 = hydrate_tArray_40_Array_8_Bit___inst0_out_1;
assign O_10 = hydrate_tArray_40_Array_8_Bit___inst0_out_10;
assign O_11 = hydrate_tArray_40_Array_8_Bit___inst0_out_11;
assign O_12 = hydrate_tArray_40_Array_8_Bit___inst0_out_12;
assign O_13 = hydrate_tArray_40_Array_8_Bit___inst0_out_13;
assign O_14 = hydrate_tArray_40_Array_8_Bit___inst0_out_14;
assign O_15 = hydrate_tArray_40_Array_8_Bit___inst0_out_15;
assign O_16 = hydrate_tArray_40_Array_8_Bit___inst0_out_16;
assign O_17 = hydrate_tArray_40_Array_8_Bit___inst0_out_17;
assign O_18 = hydrate_tArray_40_Array_8_Bit___inst0_out_18;
assign O_19 = hydrate_tArray_40_Array_8_Bit___inst0_out_19;
assign O_2 = hydrate_tArray_40_Array_8_Bit___inst0_out_2;
assign O_20 = hydrate_tArray_40_Array_8_Bit___inst0_out_20;
assign O_21 = hydrate_tArray_40_Array_8_Bit___inst0_out_21;
assign O_22 = hydrate_tArray_40_Array_8_Bit___inst0_out_22;
assign O_23 = hydrate_tArray_40_Array_8_Bit___inst0_out_23;
assign O_24 = hydrate_tArray_40_Array_8_Bit___inst0_out_24;
assign O_25 = hydrate_tArray_40_Array_8_Bit___inst0_out_25;
assign O_26 = hydrate_tArray_40_Array_8_Bit___inst0_out_26;
assign O_27 = hydrate_tArray_40_Array_8_Bit___inst0_out_27;
assign O_28 = hydrate_tArray_40_Array_8_Bit___inst0_out_28;
assign O_29 = hydrate_tArray_40_Array_8_Bit___inst0_out_29;
assign O_3 = hydrate_tArray_40_Array_8_Bit___inst0_out_3;
assign O_30 = hydrate_tArray_40_Array_8_Bit___inst0_out_30;
assign O_31 = hydrate_tArray_40_Array_8_Bit___inst0_out_31;
assign O_32 = hydrate_tArray_40_Array_8_Bit___inst0_out_32;
assign O_33 = hydrate_tArray_40_Array_8_Bit___inst0_out_33;
assign O_34 = hydrate_tArray_40_Array_8_Bit___inst0_out_34;
assign O_35 = hydrate_tArray_40_Array_8_Bit___inst0_out_35;
assign O_36 = hydrate_tArray_40_Array_8_Bit___inst0_out_36;
assign O_37 = hydrate_tArray_40_Array_8_Bit___inst0_out_37;
assign O_38 = hydrate_tArray_40_Array_8_Bit___inst0_out_38;
assign O_39 = hydrate_tArray_40_Array_8_Bit___inst0_out_39;
assign O_4 = hydrate_tArray_40_Array_8_Bit___inst0_out_4;
assign O_5 = hydrate_tArray_40_Array_8_Bit___inst0_out_5;
assign O_6 = hydrate_tArray_40_Array_8_Bit___inst0_out_6;
assign O_7 = hydrate_tArray_40_Array_8_Bit___inst0_out_7;
assign O_8 = hydrate_tArray_40_Array_8_Bit___inst0_out_8;
assign O_9 = hydrate_tArray_40_Array_8_Bit___inst0_out_9;
endmodule

module Register1 (input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
assign O = DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
endmodule

module Register_Bitt_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] Register1_inst0_O;
wire [0:0] dehydrate_tBit_inst0_out;
wire hydrate_tBit_inst0_out;
Register1 Register1_inst0(.CLK(CLK), .I(dehydrate_tBit_inst0_out), .O(Register1_inst0_O));
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit hydrate_tBit_inst0(.in(Register1_inst0_O), .out(hydrate_tBit_inst0_out));
assign O = hydrate_tBit_inst0_out;
endmodule

module FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
wire [7:0] Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_11(I_11), .I_12(I_12), .I_13(I_13), .I_14(I_14), .I_15(I_15), .I_16(I_16), .I_17(I_17), .I_18(I_18), .I_19(I_19), .I_2(I_2), .I_20(I_20), .I_21(I_21), .I_22(I_22), .I_23(I_23), .I_24(I_24), .I_25(I_25), .I_26(I_26), .I_27(I_27), .I_28(I_28), .I_29(I_29), .I_3(I_3), .I_30(I_30), .I_31(I_31), .I_32(I_32), .I_33(I_33), .I_34(I_34), .I_35(I_35), .I_36(I_36), .I_37(I_37), .I_38(I_38), .I_39(I_39), .I_4(I_4), .I_5(I_5), .I_6(I_6), .I_7(I_7), .I_8(I_8), .I_9(I_9), .O_0(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0), .O_1(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1), .O_10(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10), .O_11(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11), .O_12(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12), .O_13(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13), .O_14(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14), .O_15(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15), .O_16(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16), .O_17(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17), .O_18(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18), .O_19(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19), .O_2(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2), .O_20(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20), .O_21(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21), .O_22(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22), .O_23(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23), .O_24(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24), .O_25(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25), .O_26(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26), .O_27(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27), .O_28(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28), .O_29(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29), .O_3(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3), .O_30(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30), .O_31(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31), .O_32(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32), .O_33(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33), .O_34(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34), .O_35(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35), .O_36(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36), .O_37(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37), .O_38(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38), .O_39(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39), .O_4(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4), .O_5(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5), .O_6(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6), .O_7(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7), .O_8(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8), .O_9(Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_1 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
assign O_10 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
assign O_11 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
assign O_12 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
assign O_13 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
assign O_14 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
assign O_15 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
assign O_16 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
assign O_17 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
assign O_18 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
assign O_19 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
assign O_2 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
assign O_20 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20;
assign O_21 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21;
assign O_22 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22;
assign O_23 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23;
assign O_24 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24;
assign O_25 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25;
assign O_26 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26;
assign O_27 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27;
assign O_28 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28;
assign O_29 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29;
assign O_3 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
assign O_30 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30;
assign O_31 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31;
assign O_32 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32;
assign O_33 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33;
assign O_34 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34;
assign O_35 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35;
assign O_36 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36;
assign O_37 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37;
assign O_38 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38;
assign O_39 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39;
assign O_4 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
assign O_5 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
assign O_6 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
assign O_7 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
assign O_8 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
assign O_9 = Register_Array_40_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] LUT_Array_8_Bit_t_1n_inst0_data;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
LUT_Array_8_Bit_t_1n LUT_Array_8_Bit_t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data(LUT_Array_8_Bit_t_1n_inst0_data));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O = LUT_Array_8_Bit_t_1n_inst0_data;
assign valid_down = coreir_const11_inst0_out[0];
endmodule

module Add_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] coreir_add8_inst0_out;
coreir_add #(.width(8)) coreir_add8_inst0(.in0(I__0), .in1(I__1), .out(coreir_add8_inst0_out));
assign O = coreir_add8_inst0_out;
assign valid_down = valid_up;
endmodule

module Module_0 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Add_Atom_inst0_O;
wire Add_Atom_inst0_valid_down;
wire [7:0] Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O;
wire Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O;
wire FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire and_inst0_out;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
Add_Atom Add_Atom_inst0(.I__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .I__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .O(Add_Atom_inst0_O), .valid_down(Add_Atom_inst0_valid_down), .valid_up(atomTupleCreator_t0Int_t1Int_inst0_valid_down));
Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .valid_down(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .O(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .valid_down(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
corebit_and and_inst0(.in0(valid_up), .in1(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I), .I1(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(and_inst0_out));
assign O = Add_Atom_inst0_O;
assign valid_down = Add_Atom_inst0_valid_down;
endmodule

module NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Module_0_inst0_O;
wire Module_0_inst0_valid_down;
wire [7:0] Module_0_inst1_O;
wire Module_0_inst1_valid_down;
wire [7:0] Module_0_inst10_O;
wire Module_0_inst10_valid_down;
wire [7:0] Module_0_inst11_O;
wire Module_0_inst11_valid_down;
wire [7:0] Module_0_inst12_O;
wire Module_0_inst12_valid_down;
wire [7:0] Module_0_inst13_O;
wire Module_0_inst13_valid_down;
wire [7:0] Module_0_inst14_O;
wire Module_0_inst14_valid_down;
wire [7:0] Module_0_inst15_O;
wire Module_0_inst15_valid_down;
wire [7:0] Module_0_inst16_O;
wire Module_0_inst16_valid_down;
wire [7:0] Module_0_inst17_O;
wire Module_0_inst17_valid_down;
wire [7:0] Module_0_inst18_O;
wire Module_0_inst18_valid_down;
wire [7:0] Module_0_inst19_O;
wire Module_0_inst19_valid_down;
wire [7:0] Module_0_inst2_O;
wire Module_0_inst2_valid_down;
wire [7:0] Module_0_inst20_O;
wire Module_0_inst20_valid_down;
wire [7:0] Module_0_inst21_O;
wire Module_0_inst21_valid_down;
wire [7:0] Module_0_inst22_O;
wire Module_0_inst22_valid_down;
wire [7:0] Module_0_inst23_O;
wire Module_0_inst23_valid_down;
wire [7:0] Module_0_inst24_O;
wire Module_0_inst24_valid_down;
wire [7:0] Module_0_inst25_O;
wire Module_0_inst25_valid_down;
wire [7:0] Module_0_inst26_O;
wire Module_0_inst26_valid_down;
wire [7:0] Module_0_inst27_O;
wire Module_0_inst27_valid_down;
wire [7:0] Module_0_inst28_O;
wire Module_0_inst28_valid_down;
wire [7:0] Module_0_inst29_O;
wire Module_0_inst29_valid_down;
wire [7:0] Module_0_inst3_O;
wire Module_0_inst3_valid_down;
wire [7:0] Module_0_inst30_O;
wire Module_0_inst30_valid_down;
wire [7:0] Module_0_inst31_O;
wire Module_0_inst31_valid_down;
wire [7:0] Module_0_inst32_O;
wire Module_0_inst32_valid_down;
wire [7:0] Module_0_inst33_O;
wire Module_0_inst33_valid_down;
wire [7:0] Module_0_inst34_O;
wire Module_0_inst34_valid_down;
wire [7:0] Module_0_inst35_O;
wire Module_0_inst35_valid_down;
wire [7:0] Module_0_inst36_O;
wire Module_0_inst36_valid_down;
wire [7:0] Module_0_inst37_O;
wire Module_0_inst37_valid_down;
wire [7:0] Module_0_inst38_O;
wire Module_0_inst38_valid_down;
wire [7:0] Module_0_inst39_O;
wire Module_0_inst39_valid_down;
wire [7:0] Module_0_inst4_O;
wire Module_0_inst4_valid_down;
wire [7:0] Module_0_inst5_O;
wire Module_0_inst5_valid_down;
wire [7:0] Module_0_inst6_O;
wire Module_0_inst6_valid_down;
wire [7:0] Module_0_inst7_O;
wire Module_0_inst7_valid_down;
wire [7:0] Module_0_inst8_O;
wire Module_0_inst8_valid_down;
wire [7:0] Module_0_inst9_O;
wire Module_0_inst9_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst11_out;
wire and_inst12_out;
wire and_inst13_out;
wire and_inst14_out;
wire and_inst15_out;
wire and_inst16_out;
wire and_inst17_out;
wire and_inst18_out;
wire and_inst19_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst26_out;
wire and_inst27_out;
wire and_inst28_out;
wire and_inst29_out;
wire and_inst3_out;
wire and_inst30_out;
wire and_inst31_out;
wire and_inst32_out;
wire and_inst33_out;
wire and_inst34_out;
wire and_inst35_out;
wire and_inst36_out;
wire and_inst37_out;
wire and_inst38_out;
wire and_inst4_out;
wire and_inst5_out;
wire and_inst6_out;
wire and_inst7_out;
wire and_inst8_out;
wire and_inst9_out;
Module_0 Module_0_inst0(.CLK(CLK), .I(I_0), .O(Module_0_inst0_O), .valid_down(Module_0_inst0_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst1(.CLK(CLK), .I(I_1), .O(Module_0_inst1_O), .valid_down(Module_0_inst1_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst10(.CLK(CLK), .I(I_10), .O(Module_0_inst10_O), .valid_down(Module_0_inst10_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst11(.CLK(CLK), .I(I_11), .O(Module_0_inst11_O), .valid_down(Module_0_inst11_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst12(.CLK(CLK), .I(I_12), .O(Module_0_inst12_O), .valid_down(Module_0_inst12_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst13(.CLK(CLK), .I(I_13), .O(Module_0_inst13_O), .valid_down(Module_0_inst13_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst14(.CLK(CLK), .I(I_14), .O(Module_0_inst14_O), .valid_down(Module_0_inst14_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst15(.CLK(CLK), .I(I_15), .O(Module_0_inst15_O), .valid_down(Module_0_inst15_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst16(.CLK(CLK), .I(I_16), .O(Module_0_inst16_O), .valid_down(Module_0_inst16_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst17(.CLK(CLK), .I(I_17), .O(Module_0_inst17_O), .valid_down(Module_0_inst17_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst18(.CLK(CLK), .I(I_18), .O(Module_0_inst18_O), .valid_down(Module_0_inst18_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst19(.CLK(CLK), .I(I_19), .O(Module_0_inst19_O), .valid_down(Module_0_inst19_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst2(.CLK(CLK), .I(I_2), .O(Module_0_inst2_O), .valid_down(Module_0_inst2_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst20(.CLK(CLK), .I(I_20), .O(Module_0_inst20_O), .valid_down(Module_0_inst20_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst21(.CLK(CLK), .I(I_21), .O(Module_0_inst21_O), .valid_down(Module_0_inst21_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst22(.CLK(CLK), .I(I_22), .O(Module_0_inst22_O), .valid_down(Module_0_inst22_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst23(.CLK(CLK), .I(I_23), .O(Module_0_inst23_O), .valid_down(Module_0_inst23_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst24(.CLK(CLK), .I(I_24), .O(Module_0_inst24_O), .valid_down(Module_0_inst24_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst25(.CLK(CLK), .I(I_25), .O(Module_0_inst25_O), .valid_down(Module_0_inst25_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst26(.CLK(CLK), .I(I_26), .O(Module_0_inst26_O), .valid_down(Module_0_inst26_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst27(.CLK(CLK), .I(I_27), .O(Module_0_inst27_O), .valid_down(Module_0_inst27_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst28(.CLK(CLK), .I(I_28), .O(Module_0_inst28_O), .valid_down(Module_0_inst28_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst29(.CLK(CLK), .I(I_29), .O(Module_0_inst29_O), .valid_down(Module_0_inst29_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst3(.CLK(CLK), .I(I_3), .O(Module_0_inst3_O), .valid_down(Module_0_inst3_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst30(.CLK(CLK), .I(I_30), .O(Module_0_inst30_O), .valid_down(Module_0_inst30_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst31(.CLK(CLK), .I(I_31), .O(Module_0_inst31_O), .valid_down(Module_0_inst31_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst32(.CLK(CLK), .I(I_32), .O(Module_0_inst32_O), .valid_down(Module_0_inst32_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst33(.CLK(CLK), .I(I_33), .O(Module_0_inst33_O), .valid_down(Module_0_inst33_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst34(.CLK(CLK), .I(I_34), .O(Module_0_inst34_O), .valid_down(Module_0_inst34_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst35(.CLK(CLK), .I(I_35), .O(Module_0_inst35_O), .valid_down(Module_0_inst35_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst36(.CLK(CLK), .I(I_36), .O(Module_0_inst36_O), .valid_down(Module_0_inst36_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst37(.CLK(CLK), .I(I_37), .O(Module_0_inst37_O), .valid_down(Module_0_inst37_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst38(.CLK(CLK), .I(I_38), .O(Module_0_inst38_O), .valid_down(Module_0_inst38_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst39(.CLK(CLK), .I(I_39), .O(Module_0_inst39_O), .valid_down(Module_0_inst39_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst4(.CLK(CLK), .I(I_4), .O(Module_0_inst4_O), .valid_down(Module_0_inst4_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst5(.CLK(CLK), .I(I_5), .O(Module_0_inst5_O), .valid_down(Module_0_inst5_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst6(.CLK(CLK), .I(I_6), .O(Module_0_inst6_O), .valid_down(Module_0_inst6_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst7(.CLK(CLK), .I(I_7), .O(Module_0_inst7_O), .valid_down(Module_0_inst7_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst8(.CLK(CLK), .I(I_8), .O(Module_0_inst8_O), .valid_down(Module_0_inst8_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst9(.CLK(CLK), .I(I_9), .O(Module_0_inst9_O), .valid_down(Module_0_inst9_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Module_0_inst0_valid_down), .in1(Module_0_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Module_0_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(Module_0_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(Module_0_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(Module_0_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(Module_0_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(Module_0_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(Module_0_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(Module_0_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(Module_0_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(Module_0_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(Module_0_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Module_0_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(Module_0_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(Module_0_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(Module_0_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(Module_0_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(Module_0_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(Module_0_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst26(.in0(and_inst25_out), .in1(Module_0_inst27_valid_down), .out(and_inst26_out));
corebit_and and_inst27(.in0(and_inst26_out), .in1(Module_0_inst28_valid_down), .out(and_inst27_out));
corebit_and and_inst28(.in0(and_inst27_out), .in1(Module_0_inst29_valid_down), .out(and_inst28_out));
corebit_and and_inst29(.in0(and_inst28_out), .in1(Module_0_inst30_valid_down), .out(and_inst29_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Module_0_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst30(.in0(and_inst29_out), .in1(Module_0_inst31_valid_down), .out(and_inst30_out));
corebit_and and_inst31(.in0(and_inst30_out), .in1(Module_0_inst32_valid_down), .out(and_inst31_out));
corebit_and and_inst32(.in0(and_inst31_out), .in1(Module_0_inst33_valid_down), .out(and_inst32_out));
corebit_and and_inst33(.in0(and_inst32_out), .in1(Module_0_inst34_valid_down), .out(and_inst33_out));
corebit_and and_inst34(.in0(and_inst33_out), .in1(Module_0_inst35_valid_down), .out(and_inst34_out));
corebit_and and_inst35(.in0(and_inst34_out), .in1(Module_0_inst36_valid_down), .out(and_inst35_out));
corebit_and and_inst36(.in0(and_inst35_out), .in1(Module_0_inst37_valid_down), .out(and_inst36_out));
corebit_and and_inst37(.in0(and_inst36_out), .in1(Module_0_inst38_valid_down), .out(and_inst37_out));
corebit_and and_inst38(.in0(and_inst37_out), .in1(Module_0_inst39_valid_down), .out(and_inst38_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Module_0_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Module_0_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Module_0_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Module_0_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(Module_0_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(Module_0_inst10_valid_down), .out(and_inst9_out));
assign O_0 = Module_0_inst0_O;
assign O_1 = Module_0_inst1_O;
assign O_10 = Module_0_inst10_O;
assign O_11 = Module_0_inst11_O;
assign O_12 = Module_0_inst12_O;
assign O_13 = Module_0_inst13_O;
assign O_14 = Module_0_inst14_O;
assign O_15 = Module_0_inst15_O;
assign O_16 = Module_0_inst16_O;
assign O_17 = Module_0_inst17_O;
assign O_18 = Module_0_inst18_O;
assign O_19 = Module_0_inst19_O;
assign O_2 = Module_0_inst2_O;
assign O_20 = Module_0_inst20_O;
assign O_21 = Module_0_inst21_O;
assign O_22 = Module_0_inst22_O;
assign O_23 = Module_0_inst23_O;
assign O_24 = Module_0_inst24_O;
assign O_25 = Module_0_inst25_O;
assign O_26 = Module_0_inst26_O;
assign O_27 = Module_0_inst27_O;
assign O_28 = Module_0_inst28_O;
assign O_29 = Module_0_inst29_O;
assign O_3 = Module_0_inst3_O;
assign O_30 = Module_0_inst30_O;
assign O_31 = Module_0_inst31_O;
assign O_32 = Module_0_inst32_O;
assign O_33 = Module_0_inst33_O;
assign O_34 = Module_0_inst34_O;
assign O_35 = Module_0_inst35_O;
assign O_36 = Module_0_inst36_O;
assign O_37 = Module_0_inst37_O;
assign O_38 = Module_0_inst38_O;
assign O_39 = Module_0_inst39_O;
assign O_4 = Module_0_inst4_O;
assign O_5 = Module_0_inst5_O;
assign O_6 = Module_0_inst6_O;
assign O_7 = Module_0_inst7_O;
assign O_8 = Module_0_inst8_O;
assign O_9 = Module_0_inst9_O;
assign valid_down = and_inst38_out;
endmodule

module Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_9/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
wire [7:0] NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
wire NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_11(I_11), .I_12(I_12), .I_13(I_13), .I_14(I_14), .I_15(I_15), .I_16(I_16), .I_17(I_17), .I_18(I_18), .I_19(I_19), .I_2(I_2), .I_20(I_20), .I_21(I_21), .I_22(I_22), .I_23(I_23), .I_24(I_24), .I_25(I_25), .I_26(I_26), .I_27(I_27), .I_28(I_28), .I_29(I_29), .I_3(I_3), .I_30(I_30), .I_31(I_31), .I_32(I_32), .I_33(I_33), .I_34(I_34), .I_35(I_35), .I_36(I_36), .I_37(I_37), .I_38(I_38), .I_39(I_39), .I_4(I_4), .I_5(I_5), .I_6(I_6), .I_7(I_7), .I_8(I_8), .I_9(I_9), .O_0(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_10(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .O_11(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .O_12(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .O_13(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .O_14(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .O_15(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .O_16(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .O_17(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .O_18(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .O_19(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .O_2(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .O_20(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .O_21(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .O_22(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .O_23(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .O_24(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .O_25(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .O_26(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .O_27(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .O_28(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .O_29(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .O_3(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .O_30(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .O_31(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .O_32(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .O_33(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .O_34(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .O_35(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .O_36(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .O_37(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .O_38(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .O_39(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .O_4(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .O_5(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .O_6(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .O_7(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .O_8(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .O_9(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .valid_down(NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(valid_up));
assign O_0 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
assign O_1 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
assign O_10 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
assign O_11 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
assign O_12 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
assign O_13 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
assign O_14 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
assign O_15 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
assign O_16 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
assign O_17 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
assign O_18 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
assign O_19 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
assign O_2 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
assign O_20 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20;
assign O_21 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21;
assign O_22 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22;
assign O_23 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23;
assign O_24 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24;
assign O_25 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25;
assign O_26 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26;
assign O_27 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27;
assign O_28 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28;
assign O_29 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29;
assign O_3 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
assign O_30 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30;
assign O_31 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31;
assign O_32 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32;
assign O_33 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33;
assign O_34 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34;
assign O_35 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35;
assign O_36 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36;
assign O_37 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37;
assign O_38 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38;
assign O_39 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39;
assign O_4 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
assign O_5 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
assign O_6 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
assign O_7 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
assign O_8 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
assign O_9 = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
assign valid_down = NativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
endmodule

module top (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_9/*verilator public*/, input [7:0] hi_0/*verilator public*/, input [7:0] hi_1/*verilator public*/, input [7:0] hi_10/*verilator public*/, input [7:0] hi_11/*verilator public*/, input [7:0] hi_12/*verilator public*/, input [7:0] hi_13/*verilator public*/, input [7:0] hi_14/*verilator public*/, input [7:0] hi_15/*verilator public*/, input [7:0] hi_16/*verilator public*/, input [7:0] hi_17/*verilator public*/, input [7:0] hi_18/*verilator public*/, input [7:0] hi_19/*verilator public*/, input [7:0] hi_2/*verilator public*/, input [7:0] hi_20/*verilator public*/, input [7:0] hi_21/*verilator public*/, input [7:0] hi_22/*verilator public*/, input [7:0] hi_23/*verilator public*/, input [7:0] hi_24/*verilator public*/, input [7:0] hi_25/*verilator public*/, input [7:0] hi_26/*verilator public*/, input [7:0] hi_27/*verilator public*/, input [7:0] hi_28/*verilator public*/, input [7:0] hi_29/*verilator public*/, input [7:0] hi_3/*verilator public*/, input [7:0] hi_30/*verilator public*/, input [7:0] hi_31/*verilator public*/, input [7:0] hi_32/*verilator public*/, input [7:0] hi_33/*verilator public*/, input [7:0] hi_34/*verilator public*/, input [7:0] hi_35/*verilator public*/, input [7:0] hi_36/*verilator public*/, input [7:0] hi_37/*verilator public*/, input [7:0] hi_38/*verilator public*/, input [7:0] hi_39/*verilator public*/, input [7:0] hi_4/*verilator public*/, input [7:0] hi_5/*verilator public*/, input [7:0] hi_6/*verilator public*/, input [7:0] hi_7/*verilator public*/, input [7:0] hi_8/*verilator public*/, input [7:0] hi_9/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9;
wire FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9;
wire FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9;
wire FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_20;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_21;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_22;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_23;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_24;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_25;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_26;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_27;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_28;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_29;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_30;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_31;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_32;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_33;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_34;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_35;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_36;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_37;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_38;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_39;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8;
wire [7:0] FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9;
wire FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
wire [7:0] Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
wire Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(hi_0), .I_1(hi_1), .I_10(hi_10), .I_11(hi_11), .I_12(hi_12), .I_13(hi_13), .I_14(hi_14), .I_15(hi_15), .I_16(hi_16), .I_17(hi_17), .I_18(hi_18), .I_19(hi_19), .I_2(hi_2), .I_20(hi_20), .I_21(hi_21), .I_22(hi_22), .I_23(hi_23), .I_24(hi_24), .I_25(hi_25), .I_26(hi_26), .I_27(hi_27), .I_28(hi_28), .I_29(hi_29), .I_3(hi_3), .I_30(hi_30), .I_31(hi_31), .I_32(hi_32), .I_33(hi_33), .I_34(hi_34), .I_35(hi_35), .I_36(hi_36), .I_37(hi_37), .I_38(hi_38), .I_39(hi_39), .I_4(hi_4), .I_5(hi_5), .I_6(hi_6), .I_7(hi_7), .I_8(hi_8), .I_9(hi_9), .O_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .O_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .O_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .O_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .O_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .O_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .O_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .O_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .O_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .O_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .O_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20), .O_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21), .O_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22), .O_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23), .O_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24), .O_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25), .O_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26), .O_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27), .O_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28), .O_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29), .O_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .O_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30), .O_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31), .O_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32), .O_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33), .O_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34), .O_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35), .O_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36), .O_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37), .O_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38), .O_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39), .O_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .O_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .O_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .O_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .O_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .O_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .valid_down(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .I_1(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .I_10(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .I_11(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .I_12(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .I_13(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .I_14(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .I_15(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .I_16(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .I_17(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .I_18(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .I_19(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .I_2(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .I_20(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .I_21(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .I_22(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .I_23(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .I_24(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .I_25(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .I_26(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .I_27(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .I_28(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .I_29(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .I_3(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .I_30(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .I_31(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .I_32(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .I_33(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .I_34(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .I_35(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .I_36(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .I_37(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .I_38(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .I_39(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .I_4(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .I_5(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .I_6(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .I_7(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .I_8(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .I_9(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .O_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .O_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .O_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .O_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .O_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .O_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .O_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .O_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .O_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .O_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .O_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .O_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .O_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20), .O_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21), .O_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22), .O_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23), .O_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24), .O_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25), .O_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26), .O_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27), .O_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28), .O_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29), .O_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .O_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30), .O_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31), .O_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32), .O_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33), .O_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34), .O_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35), .O_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36), .O_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37), .O_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38), .O_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39), .O_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .O_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .O_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .O_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .O_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .O_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .valid_down(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down));
FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .I_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .I_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .I_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .I_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .I_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .I_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .I_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .I_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .I_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .I_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .I_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .I_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .I_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20), .I_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21), .I_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22), .I_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23), .I_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24), .I_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25), .I_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26), .I_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27), .I_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28), .I_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29), .I_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .I_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30), .I_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31), .I_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32), .I_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33), .I_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34), .I_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35), .I_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36), .I_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37), .I_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38), .I_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39), .I_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .I_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .I_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .I_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .I_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .I_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .O_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .O_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .O_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .O_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .O_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .O_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .O_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .O_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .O_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .O_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .O_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .O_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .O_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20), .O_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21), .O_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22), .O_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23), .O_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24), .O_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25), .O_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26), .O_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27), .O_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28), .O_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29), .O_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .O_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30), .O_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31), .O_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32), .O_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33), .O_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34), .O_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35), .O_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36), .O_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37), .O_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38), .O_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39), .O_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .O_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .O_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .O_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .O_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .O_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .valid_down(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3(.CLK(CLK), .I_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .I_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .I_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .I_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .I_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .I_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .I_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .I_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .I_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .I_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .I_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .I_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .I_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .I_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20), .I_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21), .I_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22), .I_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23), .I_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24), .I_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25), .I_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26), .I_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27), .I_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28), .I_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29), .I_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .I_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30), .I_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31), .I_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32), .I_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33), .I_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34), .I_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35), .I_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36), .I_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37), .I_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38), .I_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39), .I_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .I_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .I_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .I_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .I_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .I_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .O_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .O_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1), .O_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10), .O_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11), .O_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12), .O_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13), .O_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14), .O_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15), .O_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16), .O_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17), .O_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18), .O_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19), .O_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2), .O_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_20), .O_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_21), .O_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_22), .O_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_23), .O_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_24), .O_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_25), .O_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_26), .O_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_27), .O_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_28), .O_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_29), .O_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3), .O_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_30), .O_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_31), .O_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_32), .O_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_33), .O_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_34), .O_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_35), .O_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_36), .O_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_37), .O_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_38), .O_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_39), .O_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4), .O_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5), .O_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6), .O_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7), .O_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8), .O_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9), .valid_down(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .valid_up(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down));
Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0(.CLK(CLK), .I_0(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I_1(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I_10(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .I_11(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .I_12(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .I_13(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .I_14(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .I_15(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .I_16(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .I_17(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .I_18(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .I_19(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .I_2(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .I_20(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20), .I_21(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21), .I_22(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22), .I_23(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23), .I_24(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24), .I_25(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25), .I_26(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26), .I_27(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27), .I_28(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28), .I_29(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29), .I_3(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .I_30(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30), .I_31(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31), .I_32(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32), .I_33(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33), .I_34(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34), .I_35(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35), .I_36(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36), .I_37(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37), .I_38(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38), .I_39(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39), .I_4(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .I_5(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .I_6(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .I_7(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .I_8(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .I_9(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .O_0(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_10(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .O_11(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .O_12(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .O_13(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .O_14(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .O_15(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .O_16(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .O_17(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .O_18(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .O_19(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .O_2(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .O_20(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .O_21(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .O_22(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .O_23(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .O_24(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .O_25(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .O_26(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .O_27(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .O_28(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .O_29(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .O_3(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .O_30(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .O_31(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .O_32(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .O_33(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .O_34(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .O_35(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .O_36(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .O_37(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .O_38(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .O_39(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .O_4(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .O_5(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .O_6(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .O_7(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .O_8(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .O_9(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .valid_down(Map_T_n5_i0_opNativeMapParallel_n40_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___I_Array_40_Array_8_In_Bit____O_Array_40_Array_8_Out_Bit____CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
assign O_0 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
assign O_1 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1;
assign O_10 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10;
assign O_11 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11;
assign O_12 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12;
assign O_13 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13;
assign O_14 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14;
assign O_15 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15;
assign O_16 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16;
assign O_17 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17;
assign O_18 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18;
assign O_19 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19;
assign O_2 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2;
assign O_20 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_20;
assign O_21 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_21;
assign O_22 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_22;
assign O_23 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_23;
assign O_24 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_24;
assign O_25 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_25;
assign O_26 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_26;
assign O_27 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_27;
assign O_28 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_28;
assign O_29 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_29;
assign O_3 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3;
assign O_30 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_30;
assign O_31 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_31;
assign O_32 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_32;
assign O_33 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_33;
assign O_34 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_34;
assign O_35 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_35;
assign O_36 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_36;
assign O_37 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_37;
assign O_38 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_38;
assign O_39 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_39;
assign O_4 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4;
assign O_5 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5;
assign O_6 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6;
assign O_7 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7;
assign O_8 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8;
assign O_9 = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9;
assign valid_down = FIFO_tTSeq_5_0_SSeq_40_Int___delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
endmodule

