// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I_0_0_0/*verilator public*/, 
  output [7:0] O_0_0_0/*verilator public*/, 
  input [7:0] I_1_0_0/*verilator public*/, 
  output [7:0] O_1_0_0/*verilator public*/, 
  input [7:0] I_2_0_0/*verilator public*/, 
  output [7:0] O_2_0_0/*verilator public*/, 
  input [7:0] I_3_0_0/*verilator public*/, 
  output [7:0] O_3_0_0/*verilator public*/, 
  input [7:0] I_4_0_0/*verilator public*/, 
  output [7:0] O_4_0_0/*verilator public*/, 
  input [7:0] I_5_0_0/*verilator public*/, 
  output [7:0] O_5_0_0/*verilator public*/, 
  input [7:0] I_6_0_0/*verilator public*/, 
  output [7:0] O_6_0_0/*verilator public*/, 
  input [7:0] I_7_0_0/*verilator public*/, 
  output [7:0] O_7_0_0/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x526_TREADY(dontcare), // @[:@1298.4]
    .io_in_x526_TDATA({I_0_0_0,I_1_0_0,I_2_0_0,I_3_0_0,I_4_0_0,I_5_0_0,I_6_0_0,I_7_0_0}), // @[:@1298.4]
    .io_in_x526_TID(8'h0),
    .io_in_x526_TDEST(8'h0),
    .io_in_x527_TVALID(valid_down), // @[:@1298.4]
    .io_in_x527_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0,O_4_0_0,O_5_0_0,O_6_0_0,O_7_0_0}), // @[:@1298.4]
    .io_in_x527_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x534_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule



module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh1a); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh1a); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x981_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh2); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x534_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x980_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  input   io_ins_3, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2, // @[:@4931.4]
  output  io_outs_3 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4935.4]
  wire  _T_23; // @[StickySelects.scala 24:52:@4936.4]
  wire  _T_24; // @[StickySelects.scala 24:21:@4937.4]
  reg  _T_27; // @[StickySelects.scala 21:22:@4939.4]
  reg [31:0] _RAND_1;
  wire  _T_28; // @[StickySelects.scala 22:54:@4940.4]
  wire  _T_29; // @[StickySelects.scala 22:54:@4941.4]
  wire  _T_31; // @[StickySelects.scala 24:52:@4942.4]
  wire  _T_32; // @[StickySelects.scala 24:21:@4943.4]
  reg  _T_35; // @[StickySelects.scala 21:22:@4945.4]
  reg [31:0] _RAND_2;
  wire  _T_36; // @[StickySelects.scala 22:54:@4946.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@4947.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@4948.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@4949.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@4951.4]
  reg [31:0] _RAND_3;
  wire  _T_45; // @[StickySelects.scala 22:54:@4953.4]
  wire  _T_47; // @[StickySelects.scala 24:52:@4954.4]
  wire  _T_48; // @[StickySelects.scala 24:21:@4955.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4935.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4936.4]
  assign _T_24 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 24:21:@4937.4]
  assign _T_28 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4940.4]
  assign _T_29 = _T_28 | io_ins_3; // @[StickySelects.scala 22:54:@4941.4]
  assign _T_31 = io_ins_1 | _T_27; // @[StickySelects.scala 24:52:@4942.4]
  assign _T_32 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 24:21:@4943.4]
  assign _T_36 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4946.4]
  assign _T_37 = _T_36 | io_ins_3; // @[StickySelects.scala 22:54:@4947.4]
  assign _T_39 = io_ins_2 | _T_35; // @[StickySelects.scala 24:52:@4948.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@4949.4]
  assign _T_45 = _T_36 | io_ins_2; // @[StickySelects.scala 22:54:@4953.4]
  assign _T_47 = io_ins_3 | _T_43; // @[StickySelects.scala 24:52:@4954.4]
  assign _T_48 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 24:21:@4955.4]
  assign io_outs_0 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 28:52:@4957.4]
  assign io_outs_1 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 28:52:@4958.4]
  assign io_outs_2 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@4959.4]
  assign io_outs_3 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 28:52:@4960.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_27 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_35 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_43 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_21) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_29) begin
        _T_27 <= 1'h0;
      end else begin
        _T_27 <= _T_31;
      end
    end
    if (reset) begin
      _T_35 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_35 <= 1'h0;
      end else begin
        _T_35 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_45) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_47;
      end
    end
  end
endmodule
module StickySelects_2( // @[:@4996.2]
  input   clock, // @[:@4997.4]
  input   reset, // @[:@4998.4]
  input   io_ins_0, // @[:@4999.4]
  input   io_ins_1, // @[:@4999.4]
  input   io_ins_2, // @[:@4999.4]
  input   io_ins_3, // @[:@4999.4]
  input   io_ins_4, // @[:@4999.4]
  input   io_ins_5, // @[:@4999.4]
  input   io_ins_6, // @[:@4999.4]
  input   io_ins_7, // @[:@4999.4]
  output  io_outs_0, // @[:@4999.4]
  output  io_outs_1, // @[:@4999.4]
  output  io_outs_2, // @[:@4999.4]
  output  io_outs_3, // @[:@4999.4]
  output  io_outs_4, // @[:@4999.4]
  output  io_outs_5, // @[:@4999.4]
  output  io_outs_6, // @[:@4999.4]
  output  io_outs_7 // @[:@4999.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@5001.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@5002.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@5003.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@5004.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@5005.4]
  wire  _T_24; // @[StickySelects.scala 22:54:@5006.4]
  wire  _T_25; // @[StickySelects.scala 22:54:@5007.4]
  wire  _T_27; // @[StickySelects.scala 24:52:@5008.4]
  wire  _T_28; // @[StickySelects.scala 24:21:@5009.4]
  reg  _T_31; // @[StickySelects.scala 21:22:@5011.4]
  reg [31:0] _RAND_1;
  wire  _T_32; // @[StickySelects.scala 22:54:@5012.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@5013.4]
  wire  _T_34; // @[StickySelects.scala 22:54:@5014.4]
  wire  _T_35; // @[StickySelects.scala 22:54:@5015.4]
  wire  _T_36; // @[StickySelects.scala 22:54:@5016.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@5017.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@5018.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@5019.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@5021.4]
  reg [31:0] _RAND_2;
  wire  _T_44; // @[StickySelects.scala 22:54:@5022.4]
  wire  _T_45; // @[StickySelects.scala 22:54:@5023.4]
  wire  _T_46; // @[StickySelects.scala 22:54:@5024.4]
  wire  _T_47; // @[StickySelects.scala 22:54:@5025.4]
  wire  _T_48; // @[StickySelects.scala 22:54:@5026.4]
  wire  _T_49; // @[StickySelects.scala 22:54:@5027.4]
  wire  _T_51; // @[StickySelects.scala 24:52:@5028.4]
  wire  _T_52; // @[StickySelects.scala 24:21:@5029.4]
  reg  _T_55; // @[StickySelects.scala 21:22:@5031.4]
  reg [31:0] _RAND_3;
  wire  _T_57; // @[StickySelects.scala 22:54:@5033.4]
  wire  _T_58; // @[StickySelects.scala 22:54:@5034.4]
  wire  _T_59; // @[StickySelects.scala 22:54:@5035.4]
  wire  _T_60; // @[StickySelects.scala 22:54:@5036.4]
  wire  _T_61; // @[StickySelects.scala 22:54:@5037.4]
  wire  _T_63; // @[StickySelects.scala 24:52:@5038.4]
  wire  _T_64; // @[StickySelects.scala 24:21:@5039.4]
  reg  _T_67; // @[StickySelects.scala 21:22:@5041.4]
  reg [31:0] _RAND_4;
  wire  _T_70; // @[StickySelects.scala 22:54:@5044.4]
  wire  _T_71; // @[StickySelects.scala 22:54:@5045.4]
  wire  _T_72; // @[StickySelects.scala 22:54:@5046.4]
  wire  _T_73; // @[StickySelects.scala 22:54:@5047.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@5048.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@5049.4]
  reg  _T_79; // @[StickySelects.scala 21:22:@5051.4]
  reg [31:0] _RAND_5;
  wire  _T_83; // @[StickySelects.scala 22:54:@5055.4]
  wire  _T_84; // @[StickySelects.scala 22:54:@5056.4]
  wire  _T_85; // @[StickySelects.scala 22:54:@5057.4]
  wire  _T_87; // @[StickySelects.scala 24:52:@5058.4]
  wire  _T_88; // @[StickySelects.scala 24:21:@5059.4]
  reg  _T_91; // @[StickySelects.scala 21:22:@5061.4]
  reg [31:0] _RAND_6;
  wire  _T_96; // @[StickySelects.scala 22:54:@5066.4]
  wire  _T_97; // @[StickySelects.scala 22:54:@5067.4]
  wire  _T_99; // @[StickySelects.scala 24:52:@5068.4]
  wire  _T_100; // @[StickySelects.scala 24:21:@5069.4]
  reg  _T_103; // @[StickySelects.scala 21:22:@5071.4]
  reg [31:0] _RAND_7;
  wire  _T_109; // @[StickySelects.scala 22:54:@5077.4]
  wire  _T_111; // @[StickySelects.scala 24:52:@5078.4]
  wire  _T_112; // @[StickySelects.scala 24:21:@5079.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@5002.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@5003.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@5004.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@5005.4]
  assign _T_24 = _T_23 | io_ins_6; // @[StickySelects.scala 22:54:@5006.4]
  assign _T_25 = _T_24 | io_ins_7; // @[StickySelects.scala 22:54:@5007.4]
  assign _T_27 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@5008.4]
  assign _T_28 = _T_25 ? 1'h0 : _T_27; // @[StickySelects.scala 24:21:@5009.4]
  assign _T_32 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@5012.4]
  assign _T_33 = _T_32 | io_ins_3; // @[StickySelects.scala 22:54:@5013.4]
  assign _T_34 = _T_33 | io_ins_4; // @[StickySelects.scala 22:54:@5014.4]
  assign _T_35 = _T_34 | io_ins_5; // @[StickySelects.scala 22:54:@5015.4]
  assign _T_36 = _T_35 | io_ins_6; // @[StickySelects.scala 22:54:@5016.4]
  assign _T_37 = _T_36 | io_ins_7; // @[StickySelects.scala 22:54:@5017.4]
  assign _T_39 = io_ins_1 | _T_31; // @[StickySelects.scala 24:52:@5018.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@5019.4]
  assign _T_44 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@5022.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 22:54:@5023.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 22:54:@5024.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 22:54:@5025.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 22:54:@5026.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 22:54:@5027.4]
  assign _T_51 = io_ins_2 | _T_43; // @[StickySelects.scala 24:52:@5028.4]
  assign _T_52 = _T_49 ? 1'h0 : _T_51; // @[StickySelects.scala 24:21:@5029.4]
  assign _T_57 = _T_44 | io_ins_2; // @[StickySelects.scala 22:54:@5033.4]
  assign _T_58 = _T_57 | io_ins_4; // @[StickySelects.scala 22:54:@5034.4]
  assign _T_59 = _T_58 | io_ins_5; // @[StickySelects.scala 22:54:@5035.4]
  assign _T_60 = _T_59 | io_ins_6; // @[StickySelects.scala 22:54:@5036.4]
  assign _T_61 = _T_60 | io_ins_7; // @[StickySelects.scala 22:54:@5037.4]
  assign _T_63 = io_ins_3 | _T_55; // @[StickySelects.scala 24:52:@5038.4]
  assign _T_64 = _T_61 ? 1'h0 : _T_63; // @[StickySelects.scala 24:21:@5039.4]
  assign _T_70 = _T_57 | io_ins_3; // @[StickySelects.scala 22:54:@5044.4]
  assign _T_71 = _T_70 | io_ins_5; // @[StickySelects.scala 22:54:@5045.4]
  assign _T_72 = _T_71 | io_ins_6; // @[StickySelects.scala 22:54:@5046.4]
  assign _T_73 = _T_72 | io_ins_7; // @[StickySelects.scala 22:54:@5047.4]
  assign _T_75 = io_ins_4 | _T_67; // @[StickySelects.scala 24:52:@5048.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@5049.4]
  assign _T_83 = _T_70 | io_ins_4; // @[StickySelects.scala 22:54:@5055.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 22:54:@5056.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 22:54:@5057.4]
  assign _T_87 = io_ins_5 | _T_79; // @[StickySelects.scala 24:52:@5058.4]
  assign _T_88 = _T_85 ? 1'h0 : _T_87; // @[StickySelects.scala 24:21:@5059.4]
  assign _T_96 = _T_83 | io_ins_5; // @[StickySelects.scala 22:54:@5066.4]
  assign _T_97 = _T_96 | io_ins_7; // @[StickySelects.scala 22:54:@5067.4]
  assign _T_99 = io_ins_6 | _T_91; // @[StickySelects.scala 24:52:@5068.4]
  assign _T_100 = _T_97 ? 1'h0 : _T_99; // @[StickySelects.scala 24:21:@5069.4]
  assign _T_109 = _T_96 | io_ins_6; // @[StickySelects.scala 22:54:@5077.4]
  assign _T_111 = io_ins_7 | _T_103; // @[StickySelects.scala 24:52:@5078.4]
  assign _T_112 = _T_109 ? 1'h0 : _T_111; // @[StickySelects.scala 24:21:@5079.4]
  assign io_outs_0 = _T_25 ? 1'h0 : _T_27; // @[StickySelects.scala 28:52:@5081.4]
  assign io_outs_1 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@5082.4]
  assign io_outs_2 = _T_49 ? 1'h0 : _T_51; // @[StickySelects.scala 28:52:@5083.4]
  assign io_outs_3 = _T_61 ? 1'h0 : _T_63; // @[StickySelects.scala 28:52:@5084.4]
  assign io_outs_4 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@5085.4]
  assign io_outs_5 = _T_85 ? 1'h0 : _T_87; // @[StickySelects.scala 28:52:@5086.4]
  assign io_outs_6 = _T_97 ? 1'h0 : _T_99; // @[StickySelects.scala 28:52:@5087.4]
  assign io_outs_7 = _T_109 ? 1'h0 : _T_111; // @[StickySelects.scala 28:52:@5088.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_31 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_43 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_55 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_67 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_79 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_91 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_103 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_25) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_27;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_31 <= 1'h0;
      end else begin
        _T_31 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_49) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_51;
      end
    end
    if (reset) begin
      _T_55 <= 1'h0;
    end else begin
      if (_T_61) begin
        _T_55 <= 1'h0;
      end else begin
        _T_55 <= _T_63;
      end
    end
    if (reset) begin
      _T_67 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_67 <= 1'h0;
      end else begin
        _T_67 <= _T_75;
      end
    end
    if (reset) begin
      _T_79 <= 1'h0;
    end else begin
      if (_T_85) begin
        _T_79 <= 1'h0;
      end else begin
        _T_79 <= _T_87;
      end
    end
    if (reset) begin
      _T_91 <= 1'h0;
    end else begin
      if (_T_97) begin
        _T_91 <= 1'h0;
      end else begin
        _T_91 <= _T_99;
      end
    end
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      if (_T_109) begin
        _T_103 <= 1'h0;
      end else begin
        _T_103 <= _T_111;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5964.2]
  input   clock, // @[:@5965.4]
  input   reset, // @[:@5966.4]
  input   io_flow, // @[:@5967.4]
  input   io_in, // @[:@5967.4]
  output  io_out // @[:@5967.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5969.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5969.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5982.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5981.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5980.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5979.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5978.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5976.4]
endmodule
module x539_lb_0( // @[:@9024.2]
  input        clock, // @[:@9025.4]
  input        reset, // @[:@9026.4]
  input  [2:0] io_rPort_23_banks_0, // @[:@9027.4]
  input        io_rPort_23_ofs_0, // @[:@9027.4]
  input        io_rPort_23_en_0, // @[:@9027.4]
  input        io_rPort_23_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_23_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_22_banks_0, // @[:@9027.4]
  input        io_rPort_22_ofs_0, // @[:@9027.4]
  input        io_rPort_22_en_0, // @[:@9027.4]
  input        io_rPort_22_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_22_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_21_banks_0, // @[:@9027.4]
  input        io_rPort_21_ofs_0, // @[:@9027.4]
  input        io_rPort_21_en_0, // @[:@9027.4]
  input        io_rPort_21_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_21_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_20_banks_0, // @[:@9027.4]
  input        io_rPort_20_ofs_0, // @[:@9027.4]
  input        io_rPort_20_en_0, // @[:@9027.4]
  input        io_rPort_20_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_20_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_19_banks_0, // @[:@9027.4]
  input        io_rPort_19_ofs_0, // @[:@9027.4]
  input        io_rPort_19_en_0, // @[:@9027.4]
  input        io_rPort_19_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_19_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_18_banks_0, // @[:@9027.4]
  input        io_rPort_18_ofs_0, // @[:@9027.4]
  input        io_rPort_18_en_0, // @[:@9027.4]
  input        io_rPort_18_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_18_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@9027.4]
  input        io_rPort_17_ofs_0, // @[:@9027.4]
  input        io_rPort_17_en_0, // @[:@9027.4]
  input        io_rPort_17_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_17_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@9027.4]
  input        io_rPort_16_ofs_0, // @[:@9027.4]
  input        io_rPort_16_en_0, // @[:@9027.4]
  input        io_rPort_16_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_16_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@9027.4]
  input        io_rPort_15_ofs_0, // @[:@9027.4]
  input        io_rPort_15_en_0, // @[:@9027.4]
  input        io_rPort_15_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_15_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@9027.4]
  input        io_rPort_14_ofs_0, // @[:@9027.4]
  input        io_rPort_14_en_0, // @[:@9027.4]
  input        io_rPort_14_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_14_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@9027.4]
  input        io_rPort_13_ofs_0, // @[:@9027.4]
  input        io_rPort_13_en_0, // @[:@9027.4]
  input        io_rPort_13_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_13_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@9027.4]
  input        io_rPort_12_ofs_0, // @[:@9027.4]
  input        io_rPort_12_en_0, // @[:@9027.4]
  input        io_rPort_12_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_12_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@9027.4]
  input        io_rPort_11_ofs_0, // @[:@9027.4]
  input        io_rPort_11_en_0, // @[:@9027.4]
  input        io_rPort_11_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_11_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@9027.4]
  input        io_rPort_10_ofs_0, // @[:@9027.4]
  input        io_rPort_10_en_0, // @[:@9027.4]
  input        io_rPort_10_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_10_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@9027.4]
  input        io_rPort_9_ofs_0, // @[:@9027.4]
  input        io_rPort_9_en_0, // @[:@9027.4]
  input        io_rPort_9_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_9_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@9027.4]
  input        io_rPort_8_ofs_0, // @[:@9027.4]
  input        io_rPort_8_en_0, // @[:@9027.4]
  input        io_rPort_8_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_8_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@9027.4]
  input        io_rPort_7_ofs_0, // @[:@9027.4]
  input        io_rPort_7_en_0, // @[:@9027.4]
  input        io_rPort_7_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_7_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@9027.4]
  input        io_rPort_6_ofs_0, // @[:@9027.4]
  input        io_rPort_6_en_0, // @[:@9027.4]
  input        io_rPort_6_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_6_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@9027.4]
  input        io_rPort_5_ofs_0, // @[:@9027.4]
  input        io_rPort_5_en_0, // @[:@9027.4]
  input        io_rPort_5_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_5_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@9027.4]
  input        io_rPort_4_ofs_0, // @[:@9027.4]
  input        io_rPort_4_en_0, // @[:@9027.4]
  input        io_rPort_4_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_4_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@9027.4]
  input        io_rPort_3_ofs_0, // @[:@9027.4]
  input        io_rPort_3_en_0, // @[:@9027.4]
  input        io_rPort_3_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_3_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@9027.4]
  input        io_rPort_2_ofs_0, // @[:@9027.4]
  input        io_rPort_2_en_0, // @[:@9027.4]
  input        io_rPort_2_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_2_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@9027.4]
  input        io_rPort_1_ofs_0, // @[:@9027.4]
  input        io_rPort_1_en_0, // @[:@9027.4]
  input        io_rPort_1_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_1_output_0, // @[:@9027.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@9027.4]
  input        io_rPort_0_ofs_0, // @[:@9027.4]
  input        io_rPort_0_en_0, // @[:@9027.4]
  input        io_rPort_0_backpressure, // @[:@9027.4]
  output [7:0] io_rPort_0_output_0, // @[:@9027.4]
  input  [2:0] io_wPort_7_banks_0, // @[:@9027.4]
  input        io_wPort_7_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_7_data_0, // @[:@9027.4]
  input        io_wPort_7_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_6_banks_0, // @[:@9027.4]
  input        io_wPort_6_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_6_data_0, // @[:@9027.4]
  input        io_wPort_6_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_5_banks_0, // @[:@9027.4]
  input        io_wPort_5_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_5_data_0, // @[:@9027.4]
  input        io_wPort_5_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_4_banks_0, // @[:@9027.4]
  input        io_wPort_4_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_4_data_0, // @[:@9027.4]
  input        io_wPort_4_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@9027.4]
  input        io_wPort_3_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_3_data_0, // @[:@9027.4]
  input        io_wPort_3_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@9027.4]
  input        io_wPort_2_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_2_data_0, // @[:@9027.4]
  input        io_wPort_2_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@9027.4]
  input        io_wPort_1_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_1_data_0, // @[:@9027.4]
  input        io_wPort_1_en_0, // @[:@9027.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@9027.4]
  input        io_wPort_0_ofs_0, // @[:@9027.4]
  input  [7:0] io_wPort_0_data_0, // @[:@9027.4]
  input        io_wPort_0_en_0 // @[:@9027.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@9238.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@9238.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@9254.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@9254.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@9270.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@9270.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@9286.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@9286.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@9302.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@9302.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@9318.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@9318.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@9334.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@9334.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@9350.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@9350.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@9366.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@9366.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@9382.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@9382.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@9398.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@9398.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@9414.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@9414.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@9430.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@9430.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@9446.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@9446.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@9462.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@9462.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@9478.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@9478.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@9778.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@9818.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@9870.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@9942.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@10002.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@10042.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@10094.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@10166.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@10226.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@10266.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@10318.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@10390.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@10450.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@10490.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 121:29:@10542.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 121:29:@10614.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@10675.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@10683.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@10691.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@10699.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@10723.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@10731.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@10739.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@10747.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@10771.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@10779.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@10787.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@10795.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@10819.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@10827.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@10835.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@10843.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@10867.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@10875.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@10883.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@10891.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@10915.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@10923.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@10931.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@10939.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@10963.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@10971.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@10979.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@10987.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@11011.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@11019.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@11027.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@11035.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@11059.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@11067.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@11075.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@11083.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@11107.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@11115.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@11123.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@11131.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@11155.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@11163.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@11171.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@11179.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@11203.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@11211.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@11219.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@11227.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@11251.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@11259.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@11267.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@11275.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@11299.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@11307.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@11315.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@11323.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@11347.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@11355.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@11363.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@11371.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@11395.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@11403.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@11411.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@11419.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@11443.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@11451.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@11459.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@11467.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@11491.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@11499.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@11507.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@11515.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@11539.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@11547.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@11555.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@11563.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@11587.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@11595.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@11603.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@11611.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@11635.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@11643.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@11651.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@11659.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@11683.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@11691.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@11699.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@11707.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@11731.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@11739.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@11747.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@11755.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@11779.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@11787.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@11795.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@11803.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@11803.4]
  wire  _T_1032; // @[MemPrimitives.scala 82:210:@9494.4]
  wire  _T_1035; // @[MemPrimitives.scala 83:102:@9496.4]
  wire  _T_1037; // @[MemPrimitives.scala 82:210:@9497.4]
  wire  _T_1040; // @[MemPrimitives.scala 83:102:@9499.4]
  wire [9:0] _T_1042; // @[Cat.scala 30:58:@9501.4]
  wire [9:0] _T_1044; // @[Cat.scala 30:58:@9503.4]
  wire [9:0] _T_1045; // @[Mux.scala 31:69:@9504.4]
  wire  _T_1050; // @[MemPrimitives.scala 82:210:@9511.4]
  wire  _T_1053; // @[MemPrimitives.scala 83:102:@9513.4]
  wire  _T_1055; // @[MemPrimitives.scala 82:210:@9514.4]
  wire  _T_1058; // @[MemPrimitives.scala 83:102:@9516.4]
  wire [9:0] _T_1060; // @[Cat.scala 30:58:@9518.4]
  wire [9:0] _T_1062; // @[Cat.scala 30:58:@9520.4]
  wire [9:0] _T_1063; // @[Mux.scala 31:69:@9521.4]
  wire  _T_1068; // @[MemPrimitives.scala 82:210:@9528.4]
  wire  _T_1071; // @[MemPrimitives.scala 83:102:@9530.4]
  wire  _T_1073; // @[MemPrimitives.scala 82:210:@9531.4]
  wire  _T_1076; // @[MemPrimitives.scala 83:102:@9533.4]
  wire [9:0] _T_1078; // @[Cat.scala 30:58:@9535.4]
  wire [9:0] _T_1080; // @[Cat.scala 30:58:@9537.4]
  wire [9:0] _T_1081; // @[Mux.scala 31:69:@9538.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@9545.4]
  wire  _T_1089; // @[MemPrimitives.scala 83:102:@9547.4]
  wire  _T_1091; // @[MemPrimitives.scala 82:210:@9548.4]
  wire  _T_1094; // @[MemPrimitives.scala 83:102:@9550.4]
  wire [9:0] _T_1096; // @[Cat.scala 30:58:@9552.4]
  wire [9:0] _T_1098; // @[Cat.scala 30:58:@9554.4]
  wire [9:0] _T_1099; // @[Mux.scala 31:69:@9555.4]
  wire  _T_1104; // @[MemPrimitives.scala 82:210:@9562.4]
  wire  _T_1107; // @[MemPrimitives.scala 83:102:@9564.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:210:@9565.4]
  wire  _T_1112; // @[MemPrimitives.scala 83:102:@9567.4]
  wire [9:0] _T_1114; // @[Cat.scala 30:58:@9569.4]
  wire [9:0] _T_1116; // @[Cat.scala 30:58:@9571.4]
  wire [9:0] _T_1117; // @[Mux.scala 31:69:@9572.4]
  wire  _T_1122; // @[MemPrimitives.scala 82:210:@9579.4]
  wire  _T_1125; // @[MemPrimitives.scala 83:102:@9581.4]
  wire  _T_1127; // @[MemPrimitives.scala 82:210:@9582.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@9584.4]
  wire [9:0] _T_1132; // @[Cat.scala 30:58:@9586.4]
  wire [9:0] _T_1134; // @[Cat.scala 30:58:@9588.4]
  wire [9:0] _T_1135; // @[Mux.scala 31:69:@9589.4]
  wire  _T_1140; // @[MemPrimitives.scala 82:210:@9596.4]
  wire  _T_1143; // @[MemPrimitives.scala 83:102:@9598.4]
  wire  _T_1145; // @[MemPrimitives.scala 82:210:@9599.4]
  wire  _T_1148; // @[MemPrimitives.scala 83:102:@9601.4]
  wire [9:0] _T_1150; // @[Cat.scala 30:58:@9603.4]
  wire [9:0] _T_1152; // @[Cat.scala 30:58:@9605.4]
  wire [9:0] _T_1153; // @[Mux.scala 31:69:@9606.4]
  wire  _T_1158; // @[MemPrimitives.scala 82:210:@9613.4]
  wire  _T_1161; // @[MemPrimitives.scala 83:102:@9615.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:210:@9616.4]
  wire  _T_1166; // @[MemPrimitives.scala 83:102:@9618.4]
  wire [9:0] _T_1168; // @[Cat.scala 30:58:@9620.4]
  wire [9:0] _T_1170; // @[Cat.scala 30:58:@9622.4]
  wire [9:0] _T_1171; // @[Mux.scala 31:69:@9623.4]
  wire  _T_1176; // @[MemPrimitives.scala 82:210:@9630.4]
  wire  _T_1179; // @[MemPrimitives.scala 83:102:@9632.4]
  wire  _T_1181; // @[MemPrimitives.scala 82:210:@9633.4]
  wire  _T_1184; // @[MemPrimitives.scala 83:102:@9635.4]
  wire [9:0] _T_1186; // @[Cat.scala 30:58:@9637.4]
  wire [9:0] _T_1188; // @[Cat.scala 30:58:@9639.4]
  wire [9:0] _T_1189; // @[Mux.scala 31:69:@9640.4]
  wire  _T_1194; // @[MemPrimitives.scala 82:210:@9647.4]
  wire  _T_1197; // @[MemPrimitives.scala 83:102:@9649.4]
  wire  _T_1199; // @[MemPrimitives.scala 82:210:@9650.4]
  wire  _T_1202; // @[MemPrimitives.scala 83:102:@9652.4]
  wire [9:0] _T_1204; // @[Cat.scala 30:58:@9654.4]
  wire [9:0] _T_1206; // @[Cat.scala 30:58:@9656.4]
  wire [9:0] _T_1207; // @[Mux.scala 31:69:@9657.4]
  wire  _T_1212; // @[MemPrimitives.scala 82:210:@9664.4]
  wire  _T_1215; // @[MemPrimitives.scala 83:102:@9666.4]
  wire  _T_1217; // @[MemPrimitives.scala 82:210:@9667.4]
  wire  _T_1220; // @[MemPrimitives.scala 83:102:@9669.4]
  wire [9:0] _T_1222; // @[Cat.scala 30:58:@9671.4]
  wire [9:0] _T_1224; // @[Cat.scala 30:58:@9673.4]
  wire [9:0] _T_1225; // @[Mux.scala 31:69:@9674.4]
  wire  _T_1230; // @[MemPrimitives.scala 82:210:@9681.4]
  wire  _T_1233; // @[MemPrimitives.scala 83:102:@9683.4]
  wire  _T_1235; // @[MemPrimitives.scala 82:210:@9684.4]
  wire  _T_1238; // @[MemPrimitives.scala 83:102:@9686.4]
  wire [9:0] _T_1240; // @[Cat.scala 30:58:@9688.4]
  wire [9:0] _T_1242; // @[Cat.scala 30:58:@9690.4]
  wire [9:0] _T_1243; // @[Mux.scala 31:69:@9691.4]
  wire  _T_1248; // @[MemPrimitives.scala 82:210:@9698.4]
  wire  _T_1251; // @[MemPrimitives.scala 83:102:@9700.4]
  wire  _T_1253; // @[MemPrimitives.scala 82:210:@9701.4]
  wire  _T_1256; // @[MemPrimitives.scala 83:102:@9703.4]
  wire [9:0] _T_1258; // @[Cat.scala 30:58:@9705.4]
  wire [9:0] _T_1260; // @[Cat.scala 30:58:@9707.4]
  wire [9:0] _T_1261; // @[Mux.scala 31:69:@9708.4]
  wire  _T_1266; // @[MemPrimitives.scala 82:210:@9715.4]
  wire  _T_1269; // @[MemPrimitives.scala 83:102:@9717.4]
  wire  _T_1271; // @[MemPrimitives.scala 82:210:@9718.4]
  wire  _T_1274; // @[MemPrimitives.scala 83:102:@9720.4]
  wire [9:0] _T_1276; // @[Cat.scala 30:58:@9722.4]
  wire [9:0] _T_1278; // @[Cat.scala 30:58:@9724.4]
  wire [9:0] _T_1279; // @[Mux.scala 31:69:@9725.4]
  wire  _T_1284; // @[MemPrimitives.scala 82:210:@9732.4]
  wire  _T_1287; // @[MemPrimitives.scala 83:102:@9734.4]
  wire  _T_1289; // @[MemPrimitives.scala 82:210:@9735.4]
  wire  _T_1292; // @[MemPrimitives.scala 83:102:@9737.4]
  wire [9:0] _T_1294; // @[Cat.scala 30:58:@9739.4]
  wire [9:0] _T_1296; // @[Cat.scala 30:58:@9741.4]
  wire [9:0] _T_1297; // @[Mux.scala 31:69:@9742.4]
  wire  _T_1302; // @[MemPrimitives.scala 82:210:@9749.4]
  wire  _T_1305; // @[MemPrimitives.scala 83:102:@9751.4]
  wire  _T_1307; // @[MemPrimitives.scala 82:210:@9752.4]
  wire  _T_1310; // @[MemPrimitives.scala 83:102:@9754.4]
  wire [9:0] _T_1312; // @[Cat.scala 30:58:@9756.4]
  wire [9:0] _T_1314; // @[Cat.scala 30:58:@9758.4]
  wire [9:0] _T_1315; // @[Mux.scala 31:69:@9759.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@9766.4]
  wire  _T_1325; // @[MemPrimitives.scala 110:210:@9769.4]
  wire  _T_1330; // @[MemPrimitives.scala 110:210:@9772.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:210:@9775.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@9785.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@9786.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@9787.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@9788.4]
  wire [2:0] _T_1344; // @[Cat.scala 30:58:@9790.4]
  wire [2:0] _T_1346; // @[Cat.scala 30:58:@9792.4]
  wire [2:0] _T_1348; // @[Cat.scala 30:58:@9794.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@9796.4]
  wire [2:0] _T_1351; // @[Mux.scala 31:69:@9797.4]
  wire [2:0] _T_1352; // @[Mux.scala 31:69:@9798.4]
  wire [2:0] _T_1353; // @[Mux.scala 31:69:@9799.4]
  wire  _T_1358; // @[MemPrimitives.scala 110:210:@9806.4]
  wire  _T_1363; // @[MemPrimitives.scala 110:210:@9809.4]
  wire  _T_1368; // @[MemPrimitives.scala 110:210:@9812.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:210:@9815.4]
  wire  _T_1377; // @[MemPrimitives.scala 123:41:@9825.4]
  wire  _T_1378; // @[MemPrimitives.scala 123:41:@9826.4]
  wire  _T_1379; // @[MemPrimitives.scala 123:41:@9827.4]
  wire  _T_1380; // @[MemPrimitives.scala 123:41:@9828.4]
  wire [2:0] _T_1382; // @[Cat.scala 30:58:@9830.4]
  wire [2:0] _T_1384; // @[Cat.scala 30:58:@9832.4]
  wire [2:0] _T_1386; // @[Cat.scala 30:58:@9834.4]
  wire [2:0] _T_1388; // @[Cat.scala 30:58:@9836.4]
  wire [2:0] _T_1389; // @[Mux.scala 31:69:@9837.4]
  wire [2:0] _T_1390; // @[Mux.scala 31:69:@9838.4]
  wire [2:0] _T_1391; // @[Mux.scala 31:69:@9839.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@9846.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:210:@9849.4]
  wire  _T_1406; // @[MemPrimitives.scala 110:210:@9852.4]
  wire  _T_1411; // @[MemPrimitives.scala 110:210:@9855.4]
  wire  _T_1416; // @[MemPrimitives.scala 110:210:@9858.4]
  wire  _T_1421; // @[MemPrimitives.scala 110:210:@9861.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@9864.4]
  wire  _T_1431; // @[MemPrimitives.scala 110:210:@9867.4]
  wire  _T_1435; // @[MemPrimitives.scala 123:41:@9881.4]
  wire  _T_1436; // @[MemPrimitives.scala 123:41:@9882.4]
  wire  _T_1437; // @[MemPrimitives.scala 123:41:@9883.4]
  wire  _T_1438; // @[MemPrimitives.scala 123:41:@9884.4]
  wire  _T_1439; // @[MemPrimitives.scala 123:41:@9885.4]
  wire  _T_1440; // @[MemPrimitives.scala 123:41:@9886.4]
  wire  _T_1441; // @[MemPrimitives.scala 123:41:@9887.4]
  wire  _T_1442; // @[MemPrimitives.scala 123:41:@9888.4]
  wire [2:0] _T_1444; // @[Cat.scala 30:58:@9890.4]
  wire [2:0] _T_1446; // @[Cat.scala 30:58:@9892.4]
  wire [2:0] _T_1448; // @[Cat.scala 30:58:@9894.4]
  wire [2:0] _T_1450; // @[Cat.scala 30:58:@9896.4]
  wire [2:0] _T_1452; // @[Cat.scala 30:58:@9898.4]
  wire [2:0] _T_1454; // @[Cat.scala 30:58:@9900.4]
  wire [2:0] _T_1456; // @[Cat.scala 30:58:@9902.4]
  wire [2:0] _T_1458; // @[Cat.scala 30:58:@9904.4]
  wire [2:0] _T_1459; // @[Mux.scala 31:69:@9905.4]
  wire [2:0] _T_1460; // @[Mux.scala 31:69:@9906.4]
  wire [2:0] _T_1461; // @[Mux.scala 31:69:@9907.4]
  wire [2:0] _T_1462; // @[Mux.scala 31:69:@9908.4]
  wire [2:0] _T_1463; // @[Mux.scala 31:69:@9909.4]
  wire [2:0] _T_1464; // @[Mux.scala 31:69:@9910.4]
  wire [2:0] _T_1465; // @[Mux.scala 31:69:@9911.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@9918.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:210:@9921.4]
  wire  _T_1480; // @[MemPrimitives.scala 110:210:@9924.4]
  wire  _T_1485; // @[MemPrimitives.scala 110:210:@9927.4]
  wire  _T_1490; // @[MemPrimitives.scala 110:210:@9930.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:210:@9933.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@9936.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:210:@9939.4]
  wire  _T_1509; // @[MemPrimitives.scala 123:41:@9953.4]
  wire  _T_1510; // @[MemPrimitives.scala 123:41:@9954.4]
  wire  _T_1511; // @[MemPrimitives.scala 123:41:@9955.4]
  wire  _T_1512; // @[MemPrimitives.scala 123:41:@9956.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@9957.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@9958.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@9959.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@9960.4]
  wire [2:0] _T_1518; // @[Cat.scala 30:58:@9962.4]
  wire [2:0] _T_1520; // @[Cat.scala 30:58:@9964.4]
  wire [2:0] _T_1522; // @[Cat.scala 30:58:@9966.4]
  wire [2:0] _T_1524; // @[Cat.scala 30:58:@9968.4]
  wire [2:0] _T_1526; // @[Cat.scala 30:58:@9970.4]
  wire [2:0] _T_1528; // @[Cat.scala 30:58:@9972.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@9974.4]
  wire [2:0] _T_1532; // @[Cat.scala 30:58:@9976.4]
  wire [2:0] _T_1533; // @[Mux.scala 31:69:@9977.4]
  wire [2:0] _T_1534; // @[Mux.scala 31:69:@9978.4]
  wire [2:0] _T_1535; // @[Mux.scala 31:69:@9979.4]
  wire [2:0] _T_1536; // @[Mux.scala 31:69:@9980.4]
  wire [2:0] _T_1537; // @[Mux.scala 31:69:@9981.4]
  wire [2:0] _T_1538; // @[Mux.scala 31:69:@9982.4]
  wire [2:0] _T_1539; // @[Mux.scala 31:69:@9983.4]
  wire  _T_1544; // @[MemPrimitives.scala 110:210:@9990.4]
  wire  _T_1549; // @[MemPrimitives.scala 110:210:@9993.4]
  wire  _T_1554; // @[MemPrimitives.scala 110:210:@9996.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:210:@9999.4]
  wire  _T_1563; // @[MemPrimitives.scala 123:41:@10009.4]
  wire  _T_1564; // @[MemPrimitives.scala 123:41:@10010.4]
  wire  _T_1565; // @[MemPrimitives.scala 123:41:@10011.4]
  wire  _T_1566; // @[MemPrimitives.scala 123:41:@10012.4]
  wire [2:0] _T_1568; // @[Cat.scala 30:58:@10014.4]
  wire [2:0] _T_1570; // @[Cat.scala 30:58:@10016.4]
  wire [2:0] _T_1572; // @[Cat.scala 30:58:@10018.4]
  wire [2:0] _T_1574; // @[Cat.scala 30:58:@10020.4]
  wire [2:0] _T_1575; // @[Mux.scala 31:69:@10021.4]
  wire [2:0] _T_1576; // @[Mux.scala 31:69:@10022.4]
  wire [2:0] _T_1577; // @[Mux.scala 31:69:@10023.4]
  wire  _T_1582; // @[MemPrimitives.scala 110:210:@10030.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:210:@10033.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@10036.4]
  wire  _T_1597; // @[MemPrimitives.scala 110:210:@10039.4]
  wire  _T_1601; // @[MemPrimitives.scala 123:41:@10049.4]
  wire  _T_1602; // @[MemPrimitives.scala 123:41:@10050.4]
  wire  _T_1603; // @[MemPrimitives.scala 123:41:@10051.4]
  wire  _T_1604; // @[MemPrimitives.scala 123:41:@10052.4]
  wire [2:0] _T_1606; // @[Cat.scala 30:58:@10054.4]
  wire [2:0] _T_1608; // @[Cat.scala 30:58:@10056.4]
  wire [2:0] _T_1610; // @[Cat.scala 30:58:@10058.4]
  wire [2:0] _T_1612; // @[Cat.scala 30:58:@10060.4]
  wire [2:0] _T_1613; // @[Mux.scala 31:69:@10061.4]
  wire [2:0] _T_1614; // @[Mux.scala 31:69:@10062.4]
  wire [2:0] _T_1615; // @[Mux.scala 31:69:@10063.4]
  wire  _T_1620; // @[MemPrimitives.scala 110:210:@10070.4]
  wire  _T_1625; // @[MemPrimitives.scala 110:210:@10073.4]
  wire  _T_1630; // @[MemPrimitives.scala 110:210:@10076.4]
  wire  _T_1635; // @[MemPrimitives.scala 110:210:@10079.4]
  wire  _T_1640; // @[MemPrimitives.scala 110:210:@10082.4]
  wire  _T_1645; // @[MemPrimitives.scala 110:210:@10085.4]
  wire  _T_1650; // @[MemPrimitives.scala 110:210:@10088.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:210:@10091.4]
  wire  _T_1659; // @[MemPrimitives.scala 123:41:@10105.4]
  wire  _T_1660; // @[MemPrimitives.scala 123:41:@10106.4]
  wire  _T_1661; // @[MemPrimitives.scala 123:41:@10107.4]
  wire  _T_1662; // @[MemPrimitives.scala 123:41:@10108.4]
  wire  _T_1663; // @[MemPrimitives.scala 123:41:@10109.4]
  wire  _T_1664; // @[MemPrimitives.scala 123:41:@10110.4]
  wire  _T_1665; // @[MemPrimitives.scala 123:41:@10111.4]
  wire  _T_1666; // @[MemPrimitives.scala 123:41:@10112.4]
  wire [2:0] _T_1668; // @[Cat.scala 30:58:@10114.4]
  wire [2:0] _T_1670; // @[Cat.scala 30:58:@10116.4]
  wire [2:0] _T_1672; // @[Cat.scala 30:58:@10118.4]
  wire [2:0] _T_1674; // @[Cat.scala 30:58:@10120.4]
  wire [2:0] _T_1676; // @[Cat.scala 30:58:@10122.4]
  wire [2:0] _T_1678; // @[Cat.scala 30:58:@10124.4]
  wire [2:0] _T_1680; // @[Cat.scala 30:58:@10126.4]
  wire [2:0] _T_1682; // @[Cat.scala 30:58:@10128.4]
  wire [2:0] _T_1683; // @[Mux.scala 31:69:@10129.4]
  wire [2:0] _T_1684; // @[Mux.scala 31:69:@10130.4]
  wire [2:0] _T_1685; // @[Mux.scala 31:69:@10131.4]
  wire [2:0] _T_1686; // @[Mux.scala 31:69:@10132.4]
  wire [2:0] _T_1687; // @[Mux.scala 31:69:@10133.4]
  wire [2:0] _T_1688; // @[Mux.scala 31:69:@10134.4]
  wire [2:0] _T_1689; // @[Mux.scala 31:69:@10135.4]
  wire  _T_1694; // @[MemPrimitives.scala 110:210:@10142.4]
  wire  _T_1699; // @[MemPrimitives.scala 110:210:@10145.4]
  wire  _T_1704; // @[MemPrimitives.scala 110:210:@10148.4]
  wire  _T_1709; // @[MemPrimitives.scala 110:210:@10151.4]
  wire  _T_1714; // @[MemPrimitives.scala 110:210:@10154.4]
  wire  _T_1719; // @[MemPrimitives.scala 110:210:@10157.4]
  wire  _T_1724; // @[MemPrimitives.scala 110:210:@10160.4]
  wire  _T_1729; // @[MemPrimitives.scala 110:210:@10163.4]
  wire  _T_1733; // @[MemPrimitives.scala 123:41:@10177.4]
  wire  _T_1734; // @[MemPrimitives.scala 123:41:@10178.4]
  wire  _T_1735; // @[MemPrimitives.scala 123:41:@10179.4]
  wire  _T_1736; // @[MemPrimitives.scala 123:41:@10180.4]
  wire  _T_1737; // @[MemPrimitives.scala 123:41:@10181.4]
  wire  _T_1738; // @[MemPrimitives.scala 123:41:@10182.4]
  wire  _T_1739; // @[MemPrimitives.scala 123:41:@10183.4]
  wire  _T_1740; // @[MemPrimitives.scala 123:41:@10184.4]
  wire [2:0] _T_1742; // @[Cat.scala 30:58:@10186.4]
  wire [2:0] _T_1744; // @[Cat.scala 30:58:@10188.4]
  wire [2:0] _T_1746; // @[Cat.scala 30:58:@10190.4]
  wire [2:0] _T_1748; // @[Cat.scala 30:58:@10192.4]
  wire [2:0] _T_1750; // @[Cat.scala 30:58:@10194.4]
  wire [2:0] _T_1752; // @[Cat.scala 30:58:@10196.4]
  wire [2:0] _T_1754; // @[Cat.scala 30:58:@10198.4]
  wire [2:0] _T_1756; // @[Cat.scala 30:58:@10200.4]
  wire [2:0] _T_1757; // @[Mux.scala 31:69:@10201.4]
  wire [2:0] _T_1758; // @[Mux.scala 31:69:@10202.4]
  wire [2:0] _T_1759; // @[Mux.scala 31:69:@10203.4]
  wire [2:0] _T_1760; // @[Mux.scala 31:69:@10204.4]
  wire [2:0] _T_1761; // @[Mux.scala 31:69:@10205.4]
  wire [2:0] _T_1762; // @[Mux.scala 31:69:@10206.4]
  wire [2:0] _T_1763; // @[Mux.scala 31:69:@10207.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@10214.4]
  wire  _T_1773; // @[MemPrimitives.scala 110:210:@10217.4]
  wire  _T_1778; // @[MemPrimitives.scala 110:210:@10220.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:210:@10223.4]
  wire  _T_1787; // @[MemPrimitives.scala 123:41:@10233.4]
  wire  _T_1788; // @[MemPrimitives.scala 123:41:@10234.4]
  wire  _T_1789; // @[MemPrimitives.scala 123:41:@10235.4]
  wire  _T_1790; // @[MemPrimitives.scala 123:41:@10236.4]
  wire [2:0] _T_1792; // @[Cat.scala 30:58:@10238.4]
  wire [2:0] _T_1794; // @[Cat.scala 30:58:@10240.4]
  wire [2:0] _T_1796; // @[Cat.scala 30:58:@10242.4]
  wire [2:0] _T_1798; // @[Cat.scala 30:58:@10244.4]
  wire [2:0] _T_1799; // @[Mux.scala 31:69:@10245.4]
  wire [2:0] _T_1800; // @[Mux.scala 31:69:@10246.4]
  wire [2:0] _T_1801; // @[Mux.scala 31:69:@10247.4]
  wire  _T_1806; // @[MemPrimitives.scala 110:210:@10254.4]
  wire  _T_1811; // @[MemPrimitives.scala 110:210:@10257.4]
  wire  _T_1816; // @[MemPrimitives.scala 110:210:@10260.4]
  wire  _T_1821; // @[MemPrimitives.scala 110:210:@10263.4]
  wire  _T_1825; // @[MemPrimitives.scala 123:41:@10273.4]
  wire  _T_1826; // @[MemPrimitives.scala 123:41:@10274.4]
  wire  _T_1827; // @[MemPrimitives.scala 123:41:@10275.4]
  wire  _T_1828; // @[MemPrimitives.scala 123:41:@10276.4]
  wire [2:0] _T_1830; // @[Cat.scala 30:58:@10278.4]
  wire [2:0] _T_1832; // @[Cat.scala 30:58:@10280.4]
  wire [2:0] _T_1834; // @[Cat.scala 30:58:@10282.4]
  wire [2:0] _T_1836; // @[Cat.scala 30:58:@10284.4]
  wire [2:0] _T_1837; // @[Mux.scala 31:69:@10285.4]
  wire [2:0] _T_1838; // @[Mux.scala 31:69:@10286.4]
  wire [2:0] _T_1839; // @[Mux.scala 31:69:@10287.4]
  wire  _T_1844; // @[MemPrimitives.scala 110:210:@10294.4]
  wire  _T_1849; // @[MemPrimitives.scala 110:210:@10297.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@10300.4]
  wire  _T_1859; // @[MemPrimitives.scala 110:210:@10303.4]
  wire  _T_1864; // @[MemPrimitives.scala 110:210:@10306.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:210:@10309.4]
  wire  _T_1874; // @[MemPrimitives.scala 110:210:@10312.4]
  wire  _T_1879; // @[MemPrimitives.scala 110:210:@10315.4]
  wire  _T_1883; // @[MemPrimitives.scala 123:41:@10329.4]
  wire  _T_1884; // @[MemPrimitives.scala 123:41:@10330.4]
  wire  _T_1885; // @[MemPrimitives.scala 123:41:@10331.4]
  wire  _T_1886; // @[MemPrimitives.scala 123:41:@10332.4]
  wire  _T_1887; // @[MemPrimitives.scala 123:41:@10333.4]
  wire  _T_1888; // @[MemPrimitives.scala 123:41:@10334.4]
  wire  _T_1889; // @[MemPrimitives.scala 123:41:@10335.4]
  wire  _T_1890; // @[MemPrimitives.scala 123:41:@10336.4]
  wire [2:0] _T_1892; // @[Cat.scala 30:58:@10338.4]
  wire [2:0] _T_1894; // @[Cat.scala 30:58:@10340.4]
  wire [2:0] _T_1896; // @[Cat.scala 30:58:@10342.4]
  wire [2:0] _T_1898; // @[Cat.scala 30:58:@10344.4]
  wire [2:0] _T_1900; // @[Cat.scala 30:58:@10346.4]
  wire [2:0] _T_1902; // @[Cat.scala 30:58:@10348.4]
  wire [2:0] _T_1904; // @[Cat.scala 30:58:@10350.4]
  wire [2:0] _T_1906; // @[Cat.scala 30:58:@10352.4]
  wire [2:0] _T_1907; // @[Mux.scala 31:69:@10353.4]
  wire [2:0] _T_1908; // @[Mux.scala 31:69:@10354.4]
  wire [2:0] _T_1909; // @[Mux.scala 31:69:@10355.4]
  wire [2:0] _T_1910; // @[Mux.scala 31:69:@10356.4]
  wire [2:0] _T_1911; // @[Mux.scala 31:69:@10357.4]
  wire [2:0] _T_1912; // @[Mux.scala 31:69:@10358.4]
  wire [2:0] _T_1913; // @[Mux.scala 31:69:@10359.4]
  wire  _T_1918; // @[MemPrimitives.scala 110:210:@10366.4]
  wire  _T_1923; // @[MemPrimitives.scala 110:210:@10369.4]
  wire  _T_1928; // @[MemPrimitives.scala 110:210:@10372.4]
  wire  _T_1933; // @[MemPrimitives.scala 110:210:@10375.4]
  wire  _T_1938; // @[MemPrimitives.scala 110:210:@10378.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:210:@10381.4]
  wire  _T_1948; // @[MemPrimitives.scala 110:210:@10384.4]
  wire  _T_1953; // @[MemPrimitives.scala 110:210:@10387.4]
  wire  _T_1957; // @[MemPrimitives.scala 123:41:@10401.4]
  wire  _T_1958; // @[MemPrimitives.scala 123:41:@10402.4]
  wire  _T_1959; // @[MemPrimitives.scala 123:41:@10403.4]
  wire  _T_1960; // @[MemPrimitives.scala 123:41:@10404.4]
  wire  _T_1961; // @[MemPrimitives.scala 123:41:@10405.4]
  wire  _T_1962; // @[MemPrimitives.scala 123:41:@10406.4]
  wire  _T_1963; // @[MemPrimitives.scala 123:41:@10407.4]
  wire  _T_1964; // @[MemPrimitives.scala 123:41:@10408.4]
  wire [2:0] _T_1966; // @[Cat.scala 30:58:@10410.4]
  wire [2:0] _T_1968; // @[Cat.scala 30:58:@10412.4]
  wire [2:0] _T_1970; // @[Cat.scala 30:58:@10414.4]
  wire [2:0] _T_1972; // @[Cat.scala 30:58:@10416.4]
  wire [2:0] _T_1974; // @[Cat.scala 30:58:@10418.4]
  wire [2:0] _T_1976; // @[Cat.scala 30:58:@10420.4]
  wire [2:0] _T_1978; // @[Cat.scala 30:58:@10422.4]
  wire [2:0] _T_1980; // @[Cat.scala 30:58:@10424.4]
  wire [2:0] _T_1981; // @[Mux.scala 31:69:@10425.4]
  wire [2:0] _T_1982; // @[Mux.scala 31:69:@10426.4]
  wire [2:0] _T_1983; // @[Mux.scala 31:69:@10427.4]
  wire [2:0] _T_1984; // @[Mux.scala 31:69:@10428.4]
  wire [2:0] _T_1985; // @[Mux.scala 31:69:@10429.4]
  wire [2:0] _T_1986; // @[Mux.scala 31:69:@10430.4]
  wire [2:0] _T_1987; // @[Mux.scala 31:69:@10431.4]
  wire  _T_1992; // @[MemPrimitives.scala 110:210:@10438.4]
  wire  _T_1997; // @[MemPrimitives.scala 110:210:@10441.4]
  wire  _T_2002; // @[MemPrimitives.scala 110:210:@10444.4]
  wire  _T_2007; // @[MemPrimitives.scala 110:210:@10447.4]
  wire  _T_2011; // @[MemPrimitives.scala 123:41:@10457.4]
  wire  _T_2012; // @[MemPrimitives.scala 123:41:@10458.4]
  wire  _T_2013; // @[MemPrimitives.scala 123:41:@10459.4]
  wire  _T_2014; // @[MemPrimitives.scala 123:41:@10460.4]
  wire [2:0] _T_2016; // @[Cat.scala 30:58:@10462.4]
  wire [2:0] _T_2018; // @[Cat.scala 30:58:@10464.4]
  wire [2:0] _T_2020; // @[Cat.scala 30:58:@10466.4]
  wire [2:0] _T_2022; // @[Cat.scala 30:58:@10468.4]
  wire [2:0] _T_2023; // @[Mux.scala 31:69:@10469.4]
  wire [2:0] _T_2024; // @[Mux.scala 31:69:@10470.4]
  wire [2:0] _T_2025; // @[Mux.scala 31:69:@10471.4]
  wire  _T_2030; // @[MemPrimitives.scala 110:210:@10478.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:210:@10481.4]
  wire  _T_2040; // @[MemPrimitives.scala 110:210:@10484.4]
  wire  _T_2045; // @[MemPrimitives.scala 110:210:@10487.4]
  wire  _T_2049; // @[MemPrimitives.scala 123:41:@10497.4]
  wire  _T_2050; // @[MemPrimitives.scala 123:41:@10498.4]
  wire  _T_2051; // @[MemPrimitives.scala 123:41:@10499.4]
  wire  _T_2052; // @[MemPrimitives.scala 123:41:@10500.4]
  wire [2:0] _T_2054; // @[Cat.scala 30:58:@10502.4]
  wire [2:0] _T_2056; // @[Cat.scala 30:58:@10504.4]
  wire [2:0] _T_2058; // @[Cat.scala 30:58:@10506.4]
  wire [2:0] _T_2060; // @[Cat.scala 30:58:@10508.4]
  wire [2:0] _T_2061; // @[Mux.scala 31:69:@10509.4]
  wire [2:0] _T_2062; // @[Mux.scala 31:69:@10510.4]
  wire [2:0] _T_2063; // @[Mux.scala 31:69:@10511.4]
  wire  _T_2068; // @[MemPrimitives.scala 110:210:@10518.4]
  wire  _T_2073; // @[MemPrimitives.scala 110:210:@10521.4]
  wire  _T_2078; // @[MemPrimitives.scala 110:210:@10524.4]
  wire  _T_2083; // @[MemPrimitives.scala 110:210:@10527.4]
  wire  _T_2088; // @[MemPrimitives.scala 110:210:@10530.4]
  wire  _T_2093; // @[MemPrimitives.scala 110:210:@10533.4]
  wire  _T_2098; // @[MemPrimitives.scala 110:210:@10536.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:210:@10539.4]
  wire  _T_2107; // @[MemPrimitives.scala 123:41:@10553.4]
  wire  _T_2108; // @[MemPrimitives.scala 123:41:@10554.4]
  wire  _T_2109; // @[MemPrimitives.scala 123:41:@10555.4]
  wire  _T_2110; // @[MemPrimitives.scala 123:41:@10556.4]
  wire  _T_2111; // @[MemPrimitives.scala 123:41:@10557.4]
  wire  _T_2112; // @[MemPrimitives.scala 123:41:@10558.4]
  wire  _T_2113; // @[MemPrimitives.scala 123:41:@10559.4]
  wire  _T_2114; // @[MemPrimitives.scala 123:41:@10560.4]
  wire [2:0] _T_2116; // @[Cat.scala 30:58:@10562.4]
  wire [2:0] _T_2118; // @[Cat.scala 30:58:@10564.4]
  wire [2:0] _T_2120; // @[Cat.scala 30:58:@10566.4]
  wire [2:0] _T_2122; // @[Cat.scala 30:58:@10568.4]
  wire [2:0] _T_2124; // @[Cat.scala 30:58:@10570.4]
  wire [2:0] _T_2126; // @[Cat.scala 30:58:@10572.4]
  wire [2:0] _T_2128; // @[Cat.scala 30:58:@10574.4]
  wire [2:0] _T_2130; // @[Cat.scala 30:58:@10576.4]
  wire [2:0] _T_2131; // @[Mux.scala 31:69:@10577.4]
  wire [2:0] _T_2132; // @[Mux.scala 31:69:@10578.4]
  wire [2:0] _T_2133; // @[Mux.scala 31:69:@10579.4]
  wire [2:0] _T_2134; // @[Mux.scala 31:69:@10580.4]
  wire [2:0] _T_2135; // @[Mux.scala 31:69:@10581.4]
  wire [2:0] _T_2136; // @[Mux.scala 31:69:@10582.4]
  wire [2:0] _T_2137; // @[Mux.scala 31:69:@10583.4]
  wire  _T_2142; // @[MemPrimitives.scala 110:210:@10590.4]
  wire  _T_2147; // @[MemPrimitives.scala 110:210:@10593.4]
  wire  _T_2152; // @[MemPrimitives.scala 110:210:@10596.4]
  wire  _T_2157; // @[MemPrimitives.scala 110:210:@10599.4]
  wire  _T_2162; // @[MemPrimitives.scala 110:210:@10602.4]
  wire  _T_2167; // @[MemPrimitives.scala 110:210:@10605.4]
  wire  _T_2172; // @[MemPrimitives.scala 110:210:@10608.4]
  wire  _T_2177; // @[MemPrimitives.scala 110:210:@10611.4]
  wire  _T_2181; // @[MemPrimitives.scala 123:41:@10625.4]
  wire  _T_2182; // @[MemPrimitives.scala 123:41:@10626.4]
  wire  _T_2183; // @[MemPrimitives.scala 123:41:@10627.4]
  wire  _T_2184; // @[MemPrimitives.scala 123:41:@10628.4]
  wire  _T_2185; // @[MemPrimitives.scala 123:41:@10629.4]
  wire  _T_2186; // @[MemPrimitives.scala 123:41:@10630.4]
  wire  _T_2187; // @[MemPrimitives.scala 123:41:@10631.4]
  wire  _T_2188; // @[MemPrimitives.scala 123:41:@10632.4]
  wire [2:0] _T_2190; // @[Cat.scala 30:58:@10634.4]
  wire [2:0] _T_2192; // @[Cat.scala 30:58:@10636.4]
  wire [2:0] _T_2194; // @[Cat.scala 30:58:@10638.4]
  wire [2:0] _T_2196; // @[Cat.scala 30:58:@10640.4]
  wire [2:0] _T_2198; // @[Cat.scala 30:58:@10642.4]
  wire [2:0] _T_2200; // @[Cat.scala 30:58:@10644.4]
  wire [2:0] _T_2202; // @[Cat.scala 30:58:@10646.4]
  wire [2:0] _T_2204; // @[Cat.scala 30:58:@10648.4]
  wire [2:0] _T_2205; // @[Mux.scala 31:69:@10649.4]
  wire [2:0] _T_2206; // @[Mux.scala 31:69:@10650.4]
  wire [2:0] _T_2207; // @[Mux.scala 31:69:@10651.4]
  wire [2:0] _T_2208; // @[Mux.scala 31:69:@10652.4]
  wire [2:0] _T_2209; // @[Mux.scala 31:69:@10653.4]
  wire [2:0] _T_2210; // @[Mux.scala 31:69:@10654.4]
  wire [2:0] _T_2211; // @[Mux.scala 31:69:@10655.4]
  wire  _T_2243; // @[package.scala 96:25:@10696.4 package.scala 96:25:@10697.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@10706.4]
  wire  _T_2240; // @[package.scala 96:25:@10688.4 package.scala 96:25:@10689.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@10707.4]
  wire  _T_2237; // @[package.scala 96:25:@10680.4 package.scala 96:25:@10681.4]
  wire  _T_2278; // @[package.scala 96:25:@10744.4 package.scala 96:25:@10745.4]
  wire [7:0] _T_2282; // @[Mux.scala 31:69:@10754.4]
  wire  _T_2275; // @[package.scala 96:25:@10736.4 package.scala 96:25:@10737.4]
  wire [7:0] _T_2283; // @[Mux.scala 31:69:@10755.4]
  wire  _T_2272; // @[package.scala 96:25:@10728.4 package.scala 96:25:@10729.4]
  wire  _T_2313; // @[package.scala 96:25:@10792.4 package.scala 96:25:@10793.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@10802.4]
  wire  _T_2310; // @[package.scala 96:25:@10784.4 package.scala 96:25:@10785.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@10803.4]
  wire  _T_2307; // @[package.scala 96:25:@10776.4 package.scala 96:25:@10777.4]
  wire  _T_2348; // @[package.scala 96:25:@10840.4 package.scala 96:25:@10841.4]
  wire [7:0] _T_2352; // @[Mux.scala 31:69:@10850.4]
  wire  _T_2345; // @[package.scala 96:25:@10832.4 package.scala 96:25:@10833.4]
  wire [7:0] _T_2353; // @[Mux.scala 31:69:@10851.4]
  wire  _T_2342; // @[package.scala 96:25:@10824.4 package.scala 96:25:@10825.4]
  wire  _T_2383; // @[package.scala 96:25:@10888.4 package.scala 96:25:@10889.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@10898.4]
  wire  _T_2380; // @[package.scala 96:25:@10880.4 package.scala 96:25:@10881.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@10899.4]
  wire  _T_2377; // @[package.scala 96:25:@10872.4 package.scala 96:25:@10873.4]
  wire  _T_2418; // @[package.scala 96:25:@10936.4 package.scala 96:25:@10937.4]
  wire [7:0] _T_2422; // @[Mux.scala 31:69:@10946.4]
  wire  _T_2415; // @[package.scala 96:25:@10928.4 package.scala 96:25:@10929.4]
  wire [7:0] _T_2423; // @[Mux.scala 31:69:@10947.4]
  wire  _T_2412; // @[package.scala 96:25:@10920.4 package.scala 96:25:@10921.4]
  wire  _T_2453; // @[package.scala 96:25:@10984.4 package.scala 96:25:@10985.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@10994.4]
  wire  _T_2450; // @[package.scala 96:25:@10976.4 package.scala 96:25:@10977.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@10995.4]
  wire  _T_2447; // @[package.scala 96:25:@10968.4 package.scala 96:25:@10969.4]
  wire  _T_2488; // @[package.scala 96:25:@11032.4 package.scala 96:25:@11033.4]
  wire [7:0] _T_2492; // @[Mux.scala 31:69:@11042.4]
  wire  _T_2485; // @[package.scala 96:25:@11024.4 package.scala 96:25:@11025.4]
  wire [7:0] _T_2493; // @[Mux.scala 31:69:@11043.4]
  wire  _T_2482; // @[package.scala 96:25:@11016.4 package.scala 96:25:@11017.4]
  wire  _T_2523; // @[package.scala 96:25:@11080.4 package.scala 96:25:@11081.4]
  wire [7:0] _T_2527; // @[Mux.scala 31:69:@11090.4]
  wire  _T_2520; // @[package.scala 96:25:@11072.4 package.scala 96:25:@11073.4]
  wire [7:0] _T_2528; // @[Mux.scala 31:69:@11091.4]
  wire  _T_2517; // @[package.scala 96:25:@11064.4 package.scala 96:25:@11065.4]
  wire  _T_2558; // @[package.scala 96:25:@11128.4 package.scala 96:25:@11129.4]
  wire [7:0] _T_2562; // @[Mux.scala 31:69:@11138.4]
  wire  _T_2555; // @[package.scala 96:25:@11120.4 package.scala 96:25:@11121.4]
  wire [7:0] _T_2563; // @[Mux.scala 31:69:@11139.4]
  wire  _T_2552; // @[package.scala 96:25:@11112.4 package.scala 96:25:@11113.4]
  wire  _T_2593; // @[package.scala 96:25:@11176.4 package.scala 96:25:@11177.4]
  wire [7:0] _T_2597; // @[Mux.scala 31:69:@11186.4]
  wire  _T_2590; // @[package.scala 96:25:@11168.4 package.scala 96:25:@11169.4]
  wire [7:0] _T_2598; // @[Mux.scala 31:69:@11187.4]
  wire  _T_2587; // @[package.scala 96:25:@11160.4 package.scala 96:25:@11161.4]
  wire  _T_2628; // @[package.scala 96:25:@11224.4 package.scala 96:25:@11225.4]
  wire [7:0] _T_2632; // @[Mux.scala 31:69:@11234.4]
  wire  _T_2625; // @[package.scala 96:25:@11216.4 package.scala 96:25:@11217.4]
  wire [7:0] _T_2633; // @[Mux.scala 31:69:@11235.4]
  wire  _T_2622; // @[package.scala 96:25:@11208.4 package.scala 96:25:@11209.4]
  wire  _T_2663; // @[package.scala 96:25:@11272.4 package.scala 96:25:@11273.4]
  wire [7:0] _T_2667; // @[Mux.scala 31:69:@11282.4]
  wire  _T_2660; // @[package.scala 96:25:@11264.4 package.scala 96:25:@11265.4]
  wire [7:0] _T_2668; // @[Mux.scala 31:69:@11283.4]
  wire  _T_2657; // @[package.scala 96:25:@11256.4 package.scala 96:25:@11257.4]
  wire  _T_2698; // @[package.scala 96:25:@11320.4 package.scala 96:25:@11321.4]
  wire [7:0] _T_2702; // @[Mux.scala 31:69:@11330.4]
  wire  _T_2695; // @[package.scala 96:25:@11312.4 package.scala 96:25:@11313.4]
  wire [7:0] _T_2703; // @[Mux.scala 31:69:@11331.4]
  wire  _T_2692; // @[package.scala 96:25:@11304.4 package.scala 96:25:@11305.4]
  wire  _T_2733; // @[package.scala 96:25:@11368.4 package.scala 96:25:@11369.4]
  wire [7:0] _T_2737; // @[Mux.scala 31:69:@11378.4]
  wire  _T_2730; // @[package.scala 96:25:@11360.4 package.scala 96:25:@11361.4]
  wire [7:0] _T_2738; // @[Mux.scala 31:69:@11379.4]
  wire  _T_2727; // @[package.scala 96:25:@11352.4 package.scala 96:25:@11353.4]
  wire  _T_2768; // @[package.scala 96:25:@11416.4 package.scala 96:25:@11417.4]
  wire [7:0] _T_2772; // @[Mux.scala 31:69:@11426.4]
  wire  _T_2765; // @[package.scala 96:25:@11408.4 package.scala 96:25:@11409.4]
  wire [7:0] _T_2773; // @[Mux.scala 31:69:@11427.4]
  wire  _T_2762; // @[package.scala 96:25:@11400.4 package.scala 96:25:@11401.4]
  wire  _T_2803; // @[package.scala 96:25:@11464.4 package.scala 96:25:@11465.4]
  wire [7:0] _T_2807; // @[Mux.scala 31:69:@11474.4]
  wire  _T_2800; // @[package.scala 96:25:@11456.4 package.scala 96:25:@11457.4]
  wire [7:0] _T_2808; // @[Mux.scala 31:69:@11475.4]
  wire  _T_2797; // @[package.scala 96:25:@11448.4 package.scala 96:25:@11449.4]
  wire  _T_2838; // @[package.scala 96:25:@11512.4 package.scala 96:25:@11513.4]
  wire [7:0] _T_2842; // @[Mux.scala 31:69:@11522.4]
  wire  _T_2835; // @[package.scala 96:25:@11504.4 package.scala 96:25:@11505.4]
  wire [7:0] _T_2843; // @[Mux.scala 31:69:@11523.4]
  wire  _T_2832; // @[package.scala 96:25:@11496.4 package.scala 96:25:@11497.4]
  wire  _T_2873; // @[package.scala 96:25:@11560.4 package.scala 96:25:@11561.4]
  wire [7:0] _T_2877; // @[Mux.scala 31:69:@11570.4]
  wire  _T_2870; // @[package.scala 96:25:@11552.4 package.scala 96:25:@11553.4]
  wire [7:0] _T_2878; // @[Mux.scala 31:69:@11571.4]
  wire  _T_2867; // @[package.scala 96:25:@11544.4 package.scala 96:25:@11545.4]
  wire  _T_2908; // @[package.scala 96:25:@11608.4 package.scala 96:25:@11609.4]
  wire [7:0] _T_2912; // @[Mux.scala 31:69:@11618.4]
  wire  _T_2905; // @[package.scala 96:25:@11600.4 package.scala 96:25:@11601.4]
  wire [7:0] _T_2913; // @[Mux.scala 31:69:@11619.4]
  wire  _T_2902; // @[package.scala 96:25:@11592.4 package.scala 96:25:@11593.4]
  wire  _T_2943; // @[package.scala 96:25:@11656.4 package.scala 96:25:@11657.4]
  wire [7:0] _T_2947; // @[Mux.scala 31:69:@11666.4]
  wire  _T_2940; // @[package.scala 96:25:@11648.4 package.scala 96:25:@11649.4]
  wire [7:0] _T_2948; // @[Mux.scala 31:69:@11667.4]
  wire  _T_2937; // @[package.scala 96:25:@11640.4 package.scala 96:25:@11641.4]
  wire  _T_2978; // @[package.scala 96:25:@11704.4 package.scala 96:25:@11705.4]
  wire [7:0] _T_2982; // @[Mux.scala 31:69:@11714.4]
  wire  _T_2975; // @[package.scala 96:25:@11696.4 package.scala 96:25:@11697.4]
  wire [7:0] _T_2983; // @[Mux.scala 31:69:@11715.4]
  wire  _T_2972; // @[package.scala 96:25:@11688.4 package.scala 96:25:@11689.4]
  wire  _T_3013; // @[package.scala 96:25:@11752.4 package.scala 96:25:@11753.4]
  wire [7:0] _T_3017; // @[Mux.scala 31:69:@11762.4]
  wire  _T_3010; // @[package.scala 96:25:@11744.4 package.scala 96:25:@11745.4]
  wire [7:0] _T_3018; // @[Mux.scala 31:69:@11763.4]
  wire  _T_3007; // @[package.scala 96:25:@11736.4 package.scala 96:25:@11737.4]
  wire  _T_3048; // @[package.scala 96:25:@11800.4 package.scala 96:25:@11801.4]
  wire [7:0] _T_3052; // @[Mux.scala 31:69:@11810.4]
  wire  _T_3045; // @[package.scala 96:25:@11792.4 package.scala 96:25:@11793.4]
  wire [7:0] _T_3053; // @[Mux.scala 31:69:@11811.4]
  wire  _T_3042; // @[package.scala 96:25:@11784.4 package.scala 96:25:@11785.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@9238.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@9254.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@9270.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@9286.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@9302.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@9318.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@9334.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@9350.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@9366.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@9382.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@9398.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@9414.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@9430.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@9446.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@9462.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@9478.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@9778.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@9818.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_2 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@9870.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7)
  );
  StickySelects_2 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@9942.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@10002.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@10042.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_2 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@10094.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7)
  );
  StickySelects_2 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@10166.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@10226.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@10266.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_2 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@10318.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7)
  );
  StickySelects_2 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@10390.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@10450.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@10490.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3)
  );
  StickySelects_2 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@10542.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7)
  );
  StickySelects_2 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@10614.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@10675.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@10683.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@10691.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@10699.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@10723.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@10731.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@10739.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@10747.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@10771.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@10779.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@10787.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@10795.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@10819.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@10827.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@10835.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@10843.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@10867.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@10875.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@10883.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@10891.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@10915.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@10923.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@10931.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@10939.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@10963.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@10971.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@10979.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@10987.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@11011.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@11019.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@11027.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@11035.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@11059.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@11067.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@11075.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@11083.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@11107.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@11115.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@11123.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@11131.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@11155.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@11163.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@11171.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@11179.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@11203.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@11211.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@11219.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@11227.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@11251.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@11259.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@11267.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@11275.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@11299.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@11307.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@11315.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@11323.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@11347.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@11355.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@11363.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@11371.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@11395.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@11403.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@11411.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@11419.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@11443.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@11451.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@11459.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@11467.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@11491.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@11499.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@11507.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@11515.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_72 ( // @[package.scala 93:22:@11539.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_73 ( // @[package.scala 93:22:@11547.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_74 ( // @[package.scala 93:22:@11555.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_75 ( // @[package.scala 93:22:@11563.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_76 ( // @[package.scala 93:22:@11587.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_77 ( // @[package.scala 93:22:@11595.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_78 ( // @[package.scala 93:22:@11603.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_79 ( // @[package.scala 93:22:@11611.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_80 ( // @[package.scala 93:22:@11635.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_81 ( // @[package.scala 93:22:@11643.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_82 ( // @[package.scala 93:22:@11651.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_83 ( // @[package.scala 93:22:@11659.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_84 ( // @[package.scala 93:22:@11683.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_85 ( // @[package.scala 93:22:@11691.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_86 ( // @[package.scala 93:22:@11699.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_87 ( // @[package.scala 93:22:@11707.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_88 ( // @[package.scala 93:22:@11731.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_89 ( // @[package.scala 93:22:@11739.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_90 ( // @[package.scala 93:22:@11747.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_91 ( // @[package.scala 93:22:@11755.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_92 ( // @[package.scala 93:22:@11779.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_93 ( // @[package.scala 93:22:@11787.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_94 ( // @[package.scala 93:22:@11795.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_95 ( // @[package.scala 93:22:@11803.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_1032 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9494.4]
  assign _T_1035 = io_wPort_1_en_0 & _T_1032; // @[MemPrimitives.scala 83:102:@9496.4]
  assign _T_1037 = io_wPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9497.4]
  assign _T_1040 = io_wPort_4_en_0 & _T_1037; // @[MemPrimitives.scala 83:102:@9499.4]
  assign _T_1042 = {_T_1035,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9501.4]
  assign _T_1044 = {_T_1040,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9503.4]
  assign _T_1045 = _T_1035 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@9504.4]
  assign _T_1050 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9511.4]
  assign _T_1053 = io_wPort_2_en_0 & _T_1050; // @[MemPrimitives.scala 83:102:@9513.4]
  assign _T_1055 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9514.4]
  assign _T_1058 = io_wPort_3_en_0 & _T_1055; // @[MemPrimitives.scala 83:102:@9516.4]
  assign _T_1060 = {_T_1053,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9518.4]
  assign _T_1062 = {_T_1058,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9520.4]
  assign _T_1063 = _T_1053 ? _T_1060 : _T_1062; // @[Mux.scala 31:69:@9521.4]
  assign _T_1068 = io_wPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9528.4]
  assign _T_1071 = io_wPort_5_en_0 & _T_1068; // @[MemPrimitives.scala 83:102:@9530.4]
  assign _T_1073 = io_wPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9531.4]
  assign _T_1076 = io_wPort_7_en_0 & _T_1073; // @[MemPrimitives.scala 83:102:@9533.4]
  assign _T_1078 = {_T_1071,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9535.4]
  assign _T_1080 = {_T_1076,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9537.4]
  assign _T_1081 = _T_1071 ? _T_1078 : _T_1080; // @[Mux.scala 31:69:@9538.4]
  assign _T_1086 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9545.4]
  assign _T_1089 = io_wPort_0_en_0 & _T_1086; // @[MemPrimitives.scala 83:102:@9547.4]
  assign _T_1091 = io_wPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@9548.4]
  assign _T_1094 = io_wPort_6_en_0 & _T_1091; // @[MemPrimitives.scala 83:102:@9550.4]
  assign _T_1096 = {_T_1089,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9552.4]
  assign _T_1098 = {_T_1094,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9554.4]
  assign _T_1099 = _T_1089 ? _T_1096 : _T_1098; // @[Mux.scala 31:69:@9555.4]
  assign _T_1104 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9562.4]
  assign _T_1107 = io_wPort_1_en_0 & _T_1104; // @[MemPrimitives.scala 83:102:@9564.4]
  assign _T_1109 = io_wPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9565.4]
  assign _T_1112 = io_wPort_4_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@9567.4]
  assign _T_1114 = {_T_1107,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9569.4]
  assign _T_1116 = {_T_1112,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9571.4]
  assign _T_1117 = _T_1107 ? _T_1114 : _T_1116; // @[Mux.scala 31:69:@9572.4]
  assign _T_1122 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9579.4]
  assign _T_1125 = io_wPort_2_en_0 & _T_1122; // @[MemPrimitives.scala 83:102:@9581.4]
  assign _T_1127 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9582.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1127; // @[MemPrimitives.scala 83:102:@9584.4]
  assign _T_1132 = {_T_1125,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9586.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9588.4]
  assign _T_1135 = _T_1125 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@9589.4]
  assign _T_1140 = io_wPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9596.4]
  assign _T_1143 = io_wPort_5_en_0 & _T_1140; // @[MemPrimitives.scala 83:102:@9598.4]
  assign _T_1145 = io_wPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9599.4]
  assign _T_1148 = io_wPort_7_en_0 & _T_1145; // @[MemPrimitives.scala 83:102:@9601.4]
  assign _T_1150 = {_T_1143,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9603.4]
  assign _T_1152 = {_T_1148,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9605.4]
  assign _T_1153 = _T_1143 ? _T_1150 : _T_1152; // @[Mux.scala 31:69:@9606.4]
  assign _T_1158 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9613.4]
  assign _T_1161 = io_wPort_0_en_0 & _T_1158; // @[MemPrimitives.scala 83:102:@9615.4]
  assign _T_1163 = io_wPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@9616.4]
  assign _T_1166 = io_wPort_6_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@9618.4]
  assign _T_1168 = {_T_1161,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9620.4]
  assign _T_1170 = {_T_1166,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9622.4]
  assign _T_1171 = _T_1161 ? _T_1168 : _T_1170; // @[Mux.scala 31:69:@9623.4]
  assign _T_1176 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9630.4]
  assign _T_1179 = io_wPort_1_en_0 & _T_1176; // @[MemPrimitives.scala 83:102:@9632.4]
  assign _T_1181 = io_wPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9633.4]
  assign _T_1184 = io_wPort_4_en_0 & _T_1181; // @[MemPrimitives.scala 83:102:@9635.4]
  assign _T_1186 = {_T_1179,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9637.4]
  assign _T_1188 = {_T_1184,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9639.4]
  assign _T_1189 = _T_1179 ? _T_1186 : _T_1188; // @[Mux.scala 31:69:@9640.4]
  assign _T_1194 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9647.4]
  assign _T_1197 = io_wPort_2_en_0 & _T_1194; // @[MemPrimitives.scala 83:102:@9649.4]
  assign _T_1199 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9650.4]
  assign _T_1202 = io_wPort_3_en_0 & _T_1199; // @[MemPrimitives.scala 83:102:@9652.4]
  assign _T_1204 = {_T_1197,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9654.4]
  assign _T_1206 = {_T_1202,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9656.4]
  assign _T_1207 = _T_1197 ? _T_1204 : _T_1206; // @[Mux.scala 31:69:@9657.4]
  assign _T_1212 = io_wPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9664.4]
  assign _T_1215 = io_wPort_5_en_0 & _T_1212; // @[MemPrimitives.scala 83:102:@9666.4]
  assign _T_1217 = io_wPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9667.4]
  assign _T_1220 = io_wPort_7_en_0 & _T_1217; // @[MemPrimitives.scala 83:102:@9669.4]
  assign _T_1222 = {_T_1215,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9671.4]
  assign _T_1224 = {_T_1220,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9673.4]
  assign _T_1225 = _T_1215 ? _T_1222 : _T_1224; // @[Mux.scala 31:69:@9674.4]
  assign _T_1230 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9681.4]
  assign _T_1233 = io_wPort_0_en_0 & _T_1230; // @[MemPrimitives.scala 83:102:@9683.4]
  assign _T_1235 = io_wPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@9684.4]
  assign _T_1238 = io_wPort_6_en_0 & _T_1235; // @[MemPrimitives.scala 83:102:@9686.4]
  assign _T_1240 = {_T_1233,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9688.4]
  assign _T_1242 = {_T_1238,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9690.4]
  assign _T_1243 = _T_1233 ? _T_1240 : _T_1242; // @[Mux.scala 31:69:@9691.4]
  assign _T_1248 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9698.4]
  assign _T_1251 = io_wPort_1_en_0 & _T_1248; // @[MemPrimitives.scala 83:102:@9700.4]
  assign _T_1253 = io_wPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9701.4]
  assign _T_1256 = io_wPort_4_en_0 & _T_1253; // @[MemPrimitives.scala 83:102:@9703.4]
  assign _T_1258 = {_T_1251,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@9705.4]
  assign _T_1260 = {_T_1256,io_wPort_4_data_0,io_wPort_4_ofs_0}; // @[Cat.scala 30:58:@9707.4]
  assign _T_1261 = _T_1251 ? _T_1258 : _T_1260; // @[Mux.scala 31:69:@9708.4]
  assign _T_1266 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9715.4]
  assign _T_1269 = io_wPort_2_en_0 & _T_1266; // @[MemPrimitives.scala 83:102:@9717.4]
  assign _T_1271 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9718.4]
  assign _T_1274 = io_wPort_3_en_0 & _T_1271; // @[MemPrimitives.scala 83:102:@9720.4]
  assign _T_1276 = {_T_1269,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@9722.4]
  assign _T_1278 = {_T_1274,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@9724.4]
  assign _T_1279 = _T_1269 ? _T_1276 : _T_1278; // @[Mux.scala 31:69:@9725.4]
  assign _T_1284 = io_wPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9732.4]
  assign _T_1287 = io_wPort_5_en_0 & _T_1284; // @[MemPrimitives.scala 83:102:@9734.4]
  assign _T_1289 = io_wPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9735.4]
  assign _T_1292 = io_wPort_7_en_0 & _T_1289; // @[MemPrimitives.scala 83:102:@9737.4]
  assign _T_1294 = {_T_1287,io_wPort_5_data_0,io_wPort_5_ofs_0}; // @[Cat.scala 30:58:@9739.4]
  assign _T_1296 = {_T_1292,io_wPort_7_data_0,io_wPort_7_ofs_0}; // @[Cat.scala 30:58:@9741.4]
  assign _T_1297 = _T_1287 ? _T_1294 : _T_1296; // @[Mux.scala 31:69:@9742.4]
  assign _T_1302 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9749.4]
  assign _T_1305 = io_wPort_0_en_0 & _T_1302; // @[MemPrimitives.scala 83:102:@9751.4]
  assign _T_1307 = io_wPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@9752.4]
  assign _T_1310 = io_wPort_6_en_0 & _T_1307; // @[MemPrimitives.scala 83:102:@9754.4]
  assign _T_1312 = {_T_1305,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@9756.4]
  assign _T_1314 = {_T_1310,io_wPort_6_data_0,io_wPort_6_ofs_0}; // @[Cat.scala 30:58:@9758.4]
  assign _T_1315 = _T_1305 ? _T_1312 : _T_1314; // @[Mux.scala 31:69:@9759.4]
  assign _T_1320 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9766.4]
  assign _T_1325 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9769.4]
  assign _T_1330 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9772.4]
  assign _T_1335 = io_rPort_23_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9775.4]
  assign _T_1339 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@9785.4]
  assign _T_1340 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@9786.4]
  assign _T_1341 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@9787.4]
  assign _T_1342 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@9788.4]
  assign _T_1344 = {_T_1339,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9790.4]
  assign _T_1346 = {_T_1340,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9792.4]
  assign _T_1348 = {_T_1341,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9794.4]
  assign _T_1350 = {_T_1342,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@9796.4]
  assign _T_1351 = _T_1341 ? _T_1348 : _T_1350; // @[Mux.scala 31:69:@9797.4]
  assign _T_1352 = _T_1340 ? _T_1346 : _T_1351; // @[Mux.scala 31:69:@9798.4]
  assign _T_1353 = _T_1339 ? _T_1344 : _T_1352; // @[Mux.scala 31:69:@9799.4]
  assign _T_1358 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9806.4]
  assign _T_1363 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9809.4]
  assign _T_1368 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9812.4]
  assign _T_1373 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9815.4]
  assign _T_1377 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@9825.4]
  assign _T_1378 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@9826.4]
  assign _T_1379 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@9827.4]
  assign _T_1380 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@9828.4]
  assign _T_1382 = {_T_1377,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9830.4]
  assign _T_1384 = {_T_1378,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9832.4]
  assign _T_1386 = {_T_1379,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@9834.4]
  assign _T_1388 = {_T_1380,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@9836.4]
  assign _T_1389 = _T_1379 ? _T_1386 : _T_1388; // @[Mux.scala 31:69:@9837.4]
  assign _T_1390 = _T_1378 ? _T_1384 : _T_1389; // @[Mux.scala 31:69:@9838.4]
  assign _T_1391 = _T_1377 ? _T_1382 : _T_1390; // @[Mux.scala 31:69:@9839.4]
  assign _T_1396 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9846.4]
  assign _T_1401 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9849.4]
  assign _T_1406 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9852.4]
  assign _T_1411 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9855.4]
  assign _T_1416 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9858.4]
  assign _T_1421 = io_rPort_19_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9861.4]
  assign _T_1426 = io_rPort_20_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9864.4]
  assign _T_1431 = io_rPort_22_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9867.4]
  assign _T_1435 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@9881.4]
  assign _T_1436 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@9882.4]
  assign _T_1437 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@9883.4]
  assign _T_1438 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@9884.4]
  assign _T_1439 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@9885.4]
  assign _T_1440 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@9886.4]
  assign _T_1441 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@9887.4]
  assign _T_1442 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@9888.4]
  assign _T_1444 = {_T_1435,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9890.4]
  assign _T_1446 = {_T_1436,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9892.4]
  assign _T_1448 = {_T_1437,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9894.4]
  assign _T_1450 = {_T_1438,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@9896.4]
  assign _T_1452 = {_T_1439,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@9898.4]
  assign _T_1454 = {_T_1440,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@9900.4]
  assign _T_1456 = {_T_1441,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@9902.4]
  assign _T_1458 = {_T_1442,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@9904.4]
  assign _T_1459 = _T_1441 ? _T_1456 : _T_1458; // @[Mux.scala 31:69:@9905.4]
  assign _T_1460 = _T_1440 ? _T_1454 : _T_1459; // @[Mux.scala 31:69:@9906.4]
  assign _T_1461 = _T_1439 ? _T_1452 : _T_1460; // @[Mux.scala 31:69:@9907.4]
  assign _T_1462 = _T_1438 ? _T_1450 : _T_1461; // @[Mux.scala 31:69:@9908.4]
  assign _T_1463 = _T_1437 ? _T_1448 : _T_1462; // @[Mux.scala 31:69:@9909.4]
  assign _T_1464 = _T_1436 ? _T_1446 : _T_1463; // @[Mux.scala 31:69:@9910.4]
  assign _T_1465 = _T_1435 ? _T_1444 : _T_1464; // @[Mux.scala 31:69:@9911.4]
  assign _T_1470 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9918.4]
  assign _T_1475 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9921.4]
  assign _T_1480 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9924.4]
  assign _T_1485 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9927.4]
  assign _T_1490 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9930.4]
  assign _T_1495 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9933.4]
  assign _T_1500 = io_rPort_18_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9936.4]
  assign _T_1505 = io_rPort_21_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@9939.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@9953.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@9954.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@9955.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@9956.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@9957.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@9958.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@9959.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@9960.4]
  assign _T_1518 = {_T_1509,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9962.4]
  assign _T_1520 = {_T_1510,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9964.4]
  assign _T_1522 = {_T_1511,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9966.4]
  assign _T_1524 = {_T_1512,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9968.4]
  assign _T_1526 = {_T_1513,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@9970.4]
  assign _T_1528 = {_T_1514,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@9972.4]
  assign _T_1530 = {_T_1515,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@9974.4]
  assign _T_1532 = {_T_1516,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@9976.4]
  assign _T_1533 = _T_1515 ? _T_1530 : _T_1532; // @[Mux.scala 31:69:@9977.4]
  assign _T_1534 = _T_1514 ? _T_1528 : _T_1533; // @[Mux.scala 31:69:@9978.4]
  assign _T_1535 = _T_1513 ? _T_1526 : _T_1534; // @[Mux.scala 31:69:@9979.4]
  assign _T_1536 = _T_1512 ? _T_1524 : _T_1535; // @[Mux.scala 31:69:@9980.4]
  assign _T_1537 = _T_1511 ? _T_1522 : _T_1536; // @[Mux.scala 31:69:@9981.4]
  assign _T_1538 = _T_1510 ? _T_1520 : _T_1537; // @[Mux.scala 31:69:@9982.4]
  assign _T_1539 = _T_1509 ? _T_1518 : _T_1538; // @[Mux.scala 31:69:@9983.4]
  assign _T_1544 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9990.4]
  assign _T_1549 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9993.4]
  assign _T_1554 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9996.4]
  assign _T_1559 = io_rPort_23_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@9999.4]
  assign _T_1563 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@10009.4]
  assign _T_1564 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@10010.4]
  assign _T_1565 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@10011.4]
  assign _T_1566 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@10012.4]
  assign _T_1568 = {_T_1563,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10014.4]
  assign _T_1570 = {_T_1564,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10016.4]
  assign _T_1572 = {_T_1565,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10018.4]
  assign _T_1574 = {_T_1566,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10020.4]
  assign _T_1575 = _T_1565 ? _T_1572 : _T_1574; // @[Mux.scala 31:69:@10021.4]
  assign _T_1576 = _T_1564 ? _T_1570 : _T_1575; // @[Mux.scala 31:69:@10022.4]
  assign _T_1577 = _T_1563 ? _T_1568 : _T_1576; // @[Mux.scala 31:69:@10023.4]
  assign _T_1582 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10030.4]
  assign _T_1587 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10033.4]
  assign _T_1592 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10036.4]
  assign _T_1597 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10039.4]
  assign _T_1601 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@10049.4]
  assign _T_1602 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@10050.4]
  assign _T_1603 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@10051.4]
  assign _T_1604 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@10052.4]
  assign _T_1606 = {_T_1601,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10054.4]
  assign _T_1608 = {_T_1602,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10056.4]
  assign _T_1610 = {_T_1603,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10058.4]
  assign _T_1612 = {_T_1604,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10060.4]
  assign _T_1613 = _T_1603 ? _T_1610 : _T_1612; // @[Mux.scala 31:69:@10061.4]
  assign _T_1614 = _T_1602 ? _T_1608 : _T_1613; // @[Mux.scala 31:69:@10062.4]
  assign _T_1615 = _T_1601 ? _T_1606 : _T_1614; // @[Mux.scala 31:69:@10063.4]
  assign _T_1620 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10070.4]
  assign _T_1625 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10073.4]
  assign _T_1630 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10076.4]
  assign _T_1635 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10079.4]
  assign _T_1640 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10082.4]
  assign _T_1645 = io_rPort_19_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10085.4]
  assign _T_1650 = io_rPort_20_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10088.4]
  assign _T_1655 = io_rPort_22_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10091.4]
  assign _T_1659 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@10105.4]
  assign _T_1660 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@10106.4]
  assign _T_1661 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@10107.4]
  assign _T_1662 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@10108.4]
  assign _T_1663 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@10109.4]
  assign _T_1664 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@10110.4]
  assign _T_1665 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@10111.4]
  assign _T_1666 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@10112.4]
  assign _T_1668 = {_T_1659,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10114.4]
  assign _T_1670 = {_T_1660,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10116.4]
  assign _T_1672 = {_T_1661,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10118.4]
  assign _T_1674 = {_T_1662,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10120.4]
  assign _T_1676 = {_T_1663,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10122.4]
  assign _T_1678 = {_T_1664,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10124.4]
  assign _T_1680 = {_T_1665,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10126.4]
  assign _T_1682 = {_T_1666,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10128.4]
  assign _T_1683 = _T_1665 ? _T_1680 : _T_1682; // @[Mux.scala 31:69:@10129.4]
  assign _T_1684 = _T_1664 ? _T_1678 : _T_1683; // @[Mux.scala 31:69:@10130.4]
  assign _T_1685 = _T_1663 ? _T_1676 : _T_1684; // @[Mux.scala 31:69:@10131.4]
  assign _T_1686 = _T_1662 ? _T_1674 : _T_1685; // @[Mux.scala 31:69:@10132.4]
  assign _T_1687 = _T_1661 ? _T_1672 : _T_1686; // @[Mux.scala 31:69:@10133.4]
  assign _T_1688 = _T_1660 ? _T_1670 : _T_1687; // @[Mux.scala 31:69:@10134.4]
  assign _T_1689 = _T_1659 ? _T_1668 : _T_1688; // @[Mux.scala 31:69:@10135.4]
  assign _T_1694 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10142.4]
  assign _T_1699 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10145.4]
  assign _T_1704 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10148.4]
  assign _T_1709 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10151.4]
  assign _T_1714 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10154.4]
  assign _T_1719 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10157.4]
  assign _T_1724 = io_rPort_18_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10160.4]
  assign _T_1729 = io_rPort_21_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@10163.4]
  assign _T_1733 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@10177.4]
  assign _T_1734 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@10178.4]
  assign _T_1735 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@10179.4]
  assign _T_1736 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@10180.4]
  assign _T_1737 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@10181.4]
  assign _T_1738 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@10182.4]
  assign _T_1739 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@10183.4]
  assign _T_1740 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@10184.4]
  assign _T_1742 = {_T_1733,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10186.4]
  assign _T_1744 = {_T_1734,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10188.4]
  assign _T_1746 = {_T_1735,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10190.4]
  assign _T_1748 = {_T_1736,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10192.4]
  assign _T_1750 = {_T_1737,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10194.4]
  assign _T_1752 = {_T_1738,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10196.4]
  assign _T_1754 = {_T_1739,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10198.4]
  assign _T_1756 = {_T_1740,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10200.4]
  assign _T_1757 = _T_1739 ? _T_1754 : _T_1756; // @[Mux.scala 31:69:@10201.4]
  assign _T_1758 = _T_1738 ? _T_1752 : _T_1757; // @[Mux.scala 31:69:@10202.4]
  assign _T_1759 = _T_1737 ? _T_1750 : _T_1758; // @[Mux.scala 31:69:@10203.4]
  assign _T_1760 = _T_1736 ? _T_1748 : _T_1759; // @[Mux.scala 31:69:@10204.4]
  assign _T_1761 = _T_1735 ? _T_1746 : _T_1760; // @[Mux.scala 31:69:@10205.4]
  assign _T_1762 = _T_1734 ? _T_1744 : _T_1761; // @[Mux.scala 31:69:@10206.4]
  assign _T_1763 = _T_1733 ? _T_1742 : _T_1762; // @[Mux.scala 31:69:@10207.4]
  assign _T_1768 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10214.4]
  assign _T_1773 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10217.4]
  assign _T_1778 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10220.4]
  assign _T_1783 = io_rPort_23_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10223.4]
  assign _T_1787 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@10233.4]
  assign _T_1788 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@10234.4]
  assign _T_1789 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@10235.4]
  assign _T_1790 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@10236.4]
  assign _T_1792 = {_T_1787,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10238.4]
  assign _T_1794 = {_T_1788,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10240.4]
  assign _T_1796 = {_T_1789,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10242.4]
  assign _T_1798 = {_T_1790,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10244.4]
  assign _T_1799 = _T_1789 ? _T_1796 : _T_1798; // @[Mux.scala 31:69:@10245.4]
  assign _T_1800 = _T_1788 ? _T_1794 : _T_1799; // @[Mux.scala 31:69:@10246.4]
  assign _T_1801 = _T_1787 ? _T_1792 : _T_1800; // @[Mux.scala 31:69:@10247.4]
  assign _T_1806 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10254.4]
  assign _T_1811 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10257.4]
  assign _T_1816 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10260.4]
  assign _T_1821 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10263.4]
  assign _T_1825 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@10273.4]
  assign _T_1826 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@10274.4]
  assign _T_1827 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@10275.4]
  assign _T_1828 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@10276.4]
  assign _T_1830 = {_T_1825,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10278.4]
  assign _T_1832 = {_T_1826,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10280.4]
  assign _T_1834 = {_T_1827,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10282.4]
  assign _T_1836 = {_T_1828,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10284.4]
  assign _T_1837 = _T_1827 ? _T_1834 : _T_1836; // @[Mux.scala 31:69:@10285.4]
  assign _T_1838 = _T_1826 ? _T_1832 : _T_1837; // @[Mux.scala 31:69:@10286.4]
  assign _T_1839 = _T_1825 ? _T_1830 : _T_1838; // @[Mux.scala 31:69:@10287.4]
  assign _T_1844 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10294.4]
  assign _T_1849 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10297.4]
  assign _T_1854 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10300.4]
  assign _T_1859 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10303.4]
  assign _T_1864 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10306.4]
  assign _T_1869 = io_rPort_19_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10309.4]
  assign _T_1874 = io_rPort_20_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10312.4]
  assign _T_1879 = io_rPort_22_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10315.4]
  assign _T_1883 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@10329.4]
  assign _T_1884 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@10330.4]
  assign _T_1885 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@10331.4]
  assign _T_1886 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@10332.4]
  assign _T_1887 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@10333.4]
  assign _T_1888 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@10334.4]
  assign _T_1889 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@10335.4]
  assign _T_1890 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@10336.4]
  assign _T_1892 = {_T_1883,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10338.4]
  assign _T_1894 = {_T_1884,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10340.4]
  assign _T_1896 = {_T_1885,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10342.4]
  assign _T_1898 = {_T_1886,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10344.4]
  assign _T_1900 = {_T_1887,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10346.4]
  assign _T_1902 = {_T_1888,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10348.4]
  assign _T_1904 = {_T_1889,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10350.4]
  assign _T_1906 = {_T_1890,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10352.4]
  assign _T_1907 = _T_1889 ? _T_1904 : _T_1906; // @[Mux.scala 31:69:@10353.4]
  assign _T_1908 = _T_1888 ? _T_1902 : _T_1907; // @[Mux.scala 31:69:@10354.4]
  assign _T_1909 = _T_1887 ? _T_1900 : _T_1908; // @[Mux.scala 31:69:@10355.4]
  assign _T_1910 = _T_1886 ? _T_1898 : _T_1909; // @[Mux.scala 31:69:@10356.4]
  assign _T_1911 = _T_1885 ? _T_1896 : _T_1910; // @[Mux.scala 31:69:@10357.4]
  assign _T_1912 = _T_1884 ? _T_1894 : _T_1911; // @[Mux.scala 31:69:@10358.4]
  assign _T_1913 = _T_1883 ? _T_1892 : _T_1912; // @[Mux.scala 31:69:@10359.4]
  assign _T_1918 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10366.4]
  assign _T_1923 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10369.4]
  assign _T_1928 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10372.4]
  assign _T_1933 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10375.4]
  assign _T_1938 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10378.4]
  assign _T_1943 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10381.4]
  assign _T_1948 = io_rPort_18_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10384.4]
  assign _T_1953 = io_rPort_21_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@10387.4]
  assign _T_1957 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@10401.4]
  assign _T_1958 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@10402.4]
  assign _T_1959 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@10403.4]
  assign _T_1960 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@10404.4]
  assign _T_1961 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@10405.4]
  assign _T_1962 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@10406.4]
  assign _T_1963 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@10407.4]
  assign _T_1964 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@10408.4]
  assign _T_1966 = {_T_1957,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10410.4]
  assign _T_1968 = {_T_1958,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10412.4]
  assign _T_1970 = {_T_1959,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10414.4]
  assign _T_1972 = {_T_1960,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10416.4]
  assign _T_1974 = {_T_1961,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10418.4]
  assign _T_1976 = {_T_1962,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10420.4]
  assign _T_1978 = {_T_1963,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10422.4]
  assign _T_1980 = {_T_1964,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10424.4]
  assign _T_1981 = _T_1963 ? _T_1978 : _T_1980; // @[Mux.scala 31:69:@10425.4]
  assign _T_1982 = _T_1962 ? _T_1976 : _T_1981; // @[Mux.scala 31:69:@10426.4]
  assign _T_1983 = _T_1961 ? _T_1974 : _T_1982; // @[Mux.scala 31:69:@10427.4]
  assign _T_1984 = _T_1960 ? _T_1972 : _T_1983; // @[Mux.scala 31:69:@10428.4]
  assign _T_1985 = _T_1959 ? _T_1970 : _T_1984; // @[Mux.scala 31:69:@10429.4]
  assign _T_1986 = _T_1958 ? _T_1968 : _T_1985; // @[Mux.scala 31:69:@10430.4]
  assign _T_1987 = _T_1957 ? _T_1966 : _T_1986; // @[Mux.scala 31:69:@10431.4]
  assign _T_1992 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10438.4]
  assign _T_1997 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10441.4]
  assign _T_2002 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10444.4]
  assign _T_2007 = io_rPort_23_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10447.4]
  assign _T_2011 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@10457.4]
  assign _T_2012 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@10458.4]
  assign _T_2013 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@10459.4]
  assign _T_2014 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@10460.4]
  assign _T_2016 = {_T_2011,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@10462.4]
  assign _T_2018 = {_T_2012,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@10464.4]
  assign _T_2020 = {_T_2013,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@10466.4]
  assign _T_2022 = {_T_2014,io_rPort_23_backpressure,io_rPort_23_ofs_0}; // @[Cat.scala 30:58:@10468.4]
  assign _T_2023 = _T_2013 ? _T_2020 : _T_2022; // @[Mux.scala 31:69:@10469.4]
  assign _T_2024 = _T_2012 ? _T_2018 : _T_2023; // @[Mux.scala 31:69:@10470.4]
  assign _T_2025 = _T_2011 ? _T_2016 : _T_2024; // @[Mux.scala 31:69:@10471.4]
  assign _T_2030 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10478.4]
  assign _T_2035 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10481.4]
  assign _T_2040 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10484.4]
  assign _T_2045 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10487.4]
  assign _T_2049 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@10497.4]
  assign _T_2050 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@10498.4]
  assign _T_2051 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@10499.4]
  assign _T_2052 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@10500.4]
  assign _T_2054 = {_T_2049,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@10502.4]
  assign _T_2056 = {_T_2050,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@10504.4]
  assign _T_2058 = {_T_2051,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@10506.4]
  assign _T_2060 = {_T_2052,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@10508.4]
  assign _T_2061 = _T_2051 ? _T_2058 : _T_2060; // @[Mux.scala 31:69:@10509.4]
  assign _T_2062 = _T_2050 ? _T_2056 : _T_2061; // @[Mux.scala 31:69:@10510.4]
  assign _T_2063 = _T_2049 ? _T_2054 : _T_2062; // @[Mux.scala 31:69:@10511.4]
  assign _T_2068 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10518.4]
  assign _T_2073 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10521.4]
  assign _T_2078 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10524.4]
  assign _T_2083 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10527.4]
  assign _T_2088 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10530.4]
  assign _T_2093 = io_rPort_19_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10533.4]
  assign _T_2098 = io_rPort_20_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10536.4]
  assign _T_2103 = io_rPort_22_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10539.4]
  assign _T_2107 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@10553.4]
  assign _T_2108 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@10554.4]
  assign _T_2109 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@10555.4]
  assign _T_2110 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@10556.4]
  assign _T_2111 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@10557.4]
  assign _T_2112 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@10558.4]
  assign _T_2113 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 123:41:@10559.4]
  assign _T_2114 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 123:41:@10560.4]
  assign _T_2116 = {_T_2107,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@10562.4]
  assign _T_2118 = {_T_2108,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@10564.4]
  assign _T_2120 = {_T_2109,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@10566.4]
  assign _T_2122 = {_T_2110,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@10568.4]
  assign _T_2124 = {_T_2111,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@10570.4]
  assign _T_2126 = {_T_2112,io_rPort_19_backpressure,io_rPort_19_ofs_0}; // @[Cat.scala 30:58:@10572.4]
  assign _T_2128 = {_T_2113,io_rPort_20_backpressure,io_rPort_20_ofs_0}; // @[Cat.scala 30:58:@10574.4]
  assign _T_2130 = {_T_2114,io_rPort_22_backpressure,io_rPort_22_ofs_0}; // @[Cat.scala 30:58:@10576.4]
  assign _T_2131 = _T_2113 ? _T_2128 : _T_2130; // @[Mux.scala 31:69:@10577.4]
  assign _T_2132 = _T_2112 ? _T_2126 : _T_2131; // @[Mux.scala 31:69:@10578.4]
  assign _T_2133 = _T_2111 ? _T_2124 : _T_2132; // @[Mux.scala 31:69:@10579.4]
  assign _T_2134 = _T_2110 ? _T_2122 : _T_2133; // @[Mux.scala 31:69:@10580.4]
  assign _T_2135 = _T_2109 ? _T_2120 : _T_2134; // @[Mux.scala 31:69:@10581.4]
  assign _T_2136 = _T_2108 ? _T_2118 : _T_2135; // @[Mux.scala 31:69:@10582.4]
  assign _T_2137 = _T_2107 ? _T_2116 : _T_2136; // @[Mux.scala 31:69:@10583.4]
  assign _T_2142 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10590.4]
  assign _T_2147 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10593.4]
  assign _T_2152 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10596.4]
  assign _T_2157 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10599.4]
  assign _T_2162 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10602.4]
  assign _T_2167 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10605.4]
  assign _T_2172 = io_rPort_18_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10608.4]
  assign _T_2177 = io_rPort_21_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@10611.4]
  assign _T_2181 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@10625.4]
  assign _T_2182 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@10626.4]
  assign _T_2183 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@10627.4]
  assign _T_2184 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@10628.4]
  assign _T_2185 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@10629.4]
  assign _T_2186 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@10630.4]
  assign _T_2187 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 123:41:@10631.4]
  assign _T_2188 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 123:41:@10632.4]
  assign _T_2190 = {_T_2181,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@10634.4]
  assign _T_2192 = {_T_2182,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@10636.4]
  assign _T_2194 = {_T_2183,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@10638.4]
  assign _T_2196 = {_T_2184,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@10640.4]
  assign _T_2198 = {_T_2185,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@10642.4]
  assign _T_2200 = {_T_2186,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@10644.4]
  assign _T_2202 = {_T_2187,io_rPort_18_backpressure,io_rPort_18_ofs_0}; // @[Cat.scala 30:58:@10646.4]
  assign _T_2204 = {_T_2188,io_rPort_21_backpressure,io_rPort_21_ofs_0}; // @[Cat.scala 30:58:@10648.4]
  assign _T_2205 = _T_2187 ? _T_2202 : _T_2204; // @[Mux.scala 31:69:@10649.4]
  assign _T_2206 = _T_2186 ? _T_2200 : _T_2205; // @[Mux.scala 31:69:@10650.4]
  assign _T_2207 = _T_2185 ? _T_2198 : _T_2206; // @[Mux.scala 31:69:@10651.4]
  assign _T_2208 = _T_2184 ? _T_2196 : _T_2207; // @[Mux.scala 31:69:@10652.4]
  assign _T_2209 = _T_2183 ? _T_2194 : _T_2208; // @[Mux.scala 31:69:@10653.4]
  assign _T_2210 = _T_2182 ? _T_2192 : _T_2209; // @[Mux.scala 31:69:@10654.4]
  assign _T_2211 = _T_2181 ? _T_2190 : _T_2210; // @[Mux.scala 31:69:@10655.4]
  assign _T_2243 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@10696.4 package.scala 96:25:@10697.4]
  assign _T_2247 = _T_2243 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@10706.4]
  assign _T_2240 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@10688.4 package.scala 96:25:@10689.4]
  assign _T_2248 = _T_2240 ? Mem1D_5_io_output : _T_2247; // @[Mux.scala 31:69:@10707.4]
  assign _T_2237 = RetimeWrapper_io_out; // @[package.scala 96:25:@10680.4 package.scala 96:25:@10681.4]
  assign _T_2278 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@10744.4 package.scala 96:25:@10745.4]
  assign _T_2282 = _T_2278 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10754.4]
  assign _T_2275 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@10736.4 package.scala 96:25:@10737.4]
  assign _T_2283 = _T_2275 ? Mem1D_7_io_output : _T_2282; // @[Mux.scala 31:69:@10755.4]
  assign _T_2272 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@10728.4 package.scala 96:25:@10729.4]
  assign _T_2313 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@10792.4 package.scala 96:25:@10793.4]
  assign _T_2317 = _T_2313 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@10802.4]
  assign _T_2310 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@10784.4 package.scala 96:25:@10785.4]
  assign _T_2318 = _T_2310 ? Mem1D_4_io_output : _T_2317; // @[Mux.scala 31:69:@10803.4]
  assign _T_2307 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@10776.4 package.scala 96:25:@10777.4]
  assign _T_2348 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@10840.4 package.scala 96:25:@10841.4]
  assign _T_2352 = _T_2348 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10850.4]
  assign _T_2345 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@10832.4 package.scala 96:25:@10833.4]
  assign _T_2353 = _T_2345 ? Mem1D_6_io_output : _T_2352; // @[Mux.scala 31:69:@10851.4]
  assign _T_2342 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@10824.4 package.scala 96:25:@10825.4]
  assign _T_2383 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@10888.4 package.scala 96:25:@10889.4]
  assign _T_2387 = _T_2383 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@10898.4]
  assign _T_2380 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@10880.4 package.scala 96:25:@10881.4]
  assign _T_2388 = _T_2380 ? Mem1D_4_io_output : _T_2387; // @[Mux.scala 31:69:@10899.4]
  assign _T_2377 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@10872.4 package.scala 96:25:@10873.4]
  assign _T_2418 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@10936.4 package.scala 96:25:@10937.4]
  assign _T_2422 = _T_2418 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@10946.4]
  assign _T_2415 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@10928.4 package.scala 96:25:@10929.4]
  assign _T_2423 = _T_2415 ? Mem1D_7_io_output : _T_2422; // @[Mux.scala 31:69:@10947.4]
  assign _T_2412 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@10920.4 package.scala 96:25:@10921.4]
  assign _T_2453 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@10984.4 package.scala 96:25:@10985.4]
  assign _T_2457 = _T_2453 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10994.4]
  assign _T_2450 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@10976.4 package.scala 96:25:@10977.4]
  assign _T_2458 = _T_2450 ? Mem1D_6_io_output : _T_2457; // @[Mux.scala 31:69:@10995.4]
  assign _T_2447 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@10968.4 package.scala 96:25:@10969.4]
  assign _T_2488 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@11032.4 package.scala 96:25:@11033.4]
  assign _T_2492 = _T_2488 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11042.4]
  assign _T_2485 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@11024.4 package.scala 96:25:@11025.4]
  assign _T_2493 = _T_2485 ? Mem1D_7_io_output : _T_2492; // @[Mux.scala 31:69:@11043.4]
  assign _T_2482 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@11016.4 package.scala 96:25:@11017.4]
  assign _T_2523 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@11080.4 package.scala 96:25:@11081.4]
  assign _T_2527 = _T_2523 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11090.4]
  assign _T_2520 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@11072.4 package.scala 96:25:@11073.4]
  assign _T_2528 = _T_2520 ? Mem1D_5_io_output : _T_2527; // @[Mux.scala 31:69:@11091.4]
  assign _T_2517 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@11064.4 package.scala 96:25:@11065.4]
  assign _T_2558 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@11128.4 package.scala 96:25:@11129.4]
  assign _T_2562 = _T_2558 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11138.4]
  assign _T_2555 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@11120.4 package.scala 96:25:@11121.4]
  assign _T_2563 = _T_2555 ? Mem1D_6_io_output : _T_2562; // @[Mux.scala 31:69:@11139.4]
  assign _T_2552 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@11112.4 package.scala 96:25:@11113.4]
  assign _T_2593 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@11176.4 package.scala 96:25:@11177.4]
  assign _T_2597 = _T_2593 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11186.4]
  assign _T_2590 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@11168.4 package.scala 96:25:@11169.4]
  assign _T_2598 = _T_2590 ? Mem1D_4_io_output : _T_2597; // @[Mux.scala 31:69:@11187.4]
  assign _T_2587 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@11160.4 package.scala 96:25:@11161.4]
  assign _T_2628 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@11224.4 package.scala 96:25:@11225.4]
  assign _T_2632 = _T_2628 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11234.4]
  assign _T_2625 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@11216.4 package.scala 96:25:@11217.4]
  assign _T_2633 = _T_2625 ? Mem1D_7_io_output : _T_2632; // @[Mux.scala 31:69:@11235.4]
  assign _T_2622 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@11208.4 package.scala 96:25:@11209.4]
  assign _T_2663 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@11272.4 package.scala 96:25:@11273.4]
  assign _T_2667 = _T_2663 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11282.4]
  assign _T_2660 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@11264.4 package.scala 96:25:@11265.4]
  assign _T_2668 = _T_2660 ? Mem1D_6_io_output : _T_2667; // @[Mux.scala 31:69:@11283.4]
  assign _T_2657 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@11256.4 package.scala 96:25:@11257.4]
  assign _T_2698 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@11320.4 package.scala 96:25:@11321.4]
  assign _T_2702 = _T_2698 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11330.4]
  assign _T_2695 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@11312.4 package.scala 96:25:@11313.4]
  assign _T_2703 = _T_2695 ? Mem1D_6_io_output : _T_2702; // @[Mux.scala 31:69:@11331.4]
  assign _T_2692 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@11304.4 package.scala 96:25:@11305.4]
  assign _T_2733 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@11368.4 package.scala 96:25:@11369.4]
  assign _T_2737 = _T_2733 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11378.4]
  assign _T_2730 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@11360.4 package.scala 96:25:@11361.4]
  assign _T_2738 = _T_2730 ? Mem1D_7_io_output : _T_2737; // @[Mux.scala 31:69:@11379.4]
  assign _T_2727 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@11352.4 package.scala 96:25:@11353.4]
  assign _T_2768 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@11416.4 package.scala 96:25:@11417.4]
  assign _T_2772 = _T_2768 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11426.4]
  assign _T_2765 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@11408.4 package.scala 96:25:@11409.4]
  assign _T_2773 = _T_2765 ? Mem1D_5_io_output : _T_2772; // @[Mux.scala 31:69:@11427.4]
  assign _T_2762 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@11400.4 package.scala 96:25:@11401.4]
  assign _T_2803 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@11464.4 package.scala 96:25:@11465.4]
  assign _T_2807 = _T_2803 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@11474.4]
  assign _T_2800 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@11456.4 package.scala 96:25:@11457.4]
  assign _T_2808 = _T_2800 ? Mem1D_5_io_output : _T_2807; // @[Mux.scala 31:69:@11475.4]
  assign _T_2797 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@11448.4 package.scala 96:25:@11449.4]
  assign _T_2838 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@11512.4 package.scala 96:25:@11513.4]
  assign _T_2842 = _T_2838 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11522.4]
  assign _T_2835 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@11504.4 package.scala 96:25:@11505.4]
  assign _T_2843 = _T_2835 ? Mem1D_7_io_output : _T_2842; // @[Mux.scala 31:69:@11523.4]
  assign _T_2832 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@11496.4 package.scala 96:25:@11497.4]
  assign _T_2873 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@11560.4 package.scala 96:25:@11561.4]
  assign _T_2877 = _T_2873 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11570.4]
  assign _T_2870 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@11552.4 package.scala 96:25:@11553.4]
  assign _T_2878 = _T_2870 ? Mem1D_7_io_output : _T_2877; // @[Mux.scala 31:69:@11571.4]
  assign _T_2867 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@11544.4 package.scala 96:25:@11545.4]
  assign _T_2908 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@11608.4 package.scala 96:25:@11609.4]
  assign _T_2912 = _T_2908 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11618.4]
  assign _T_2905 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@11600.4 package.scala 96:25:@11601.4]
  assign _T_2913 = _T_2905 ? Mem1D_6_io_output : _T_2912; // @[Mux.scala 31:69:@11619.4]
  assign _T_2902 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@11592.4 package.scala 96:25:@11593.4]
  assign _T_2943 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@11656.4 package.scala 96:25:@11657.4]
  assign _T_2947 = _T_2943 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11666.4]
  assign _T_2940 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@11648.4 package.scala 96:25:@11649.4]
  assign _T_2948 = _T_2940 ? Mem1D_6_io_output : _T_2947; // @[Mux.scala 31:69:@11667.4]
  assign _T_2937 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@11640.4 package.scala 96:25:@11641.4]
  assign _T_2978 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@11704.4 package.scala 96:25:@11705.4]
  assign _T_2982 = _T_2978 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@11714.4]
  assign _T_2975 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@11696.4 package.scala 96:25:@11697.4]
  assign _T_2983 = _T_2975 ? Mem1D_7_io_output : _T_2982; // @[Mux.scala 31:69:@11715.4]
  assign _T_2972 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@11688.4 package.scala 96:25:@11689.4]
  assign _T_3013 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@11752.4 package.scala 96:25:@11753.4]
  assign _T_3017 = _T_3013 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@11762.4]
  assign _T_3010 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@11744.4 package.scala 96:25:@11745.4]
  assign _T_3018 = _T_3010 ? Mem1D_6_io_output : _T_3017; // @[Mux.scala 31:69:@11763.4]
  assign _T_3007 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@11736.4 package.scala 96:25:@11737.4]
  assign _T_3048 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@11800.4 package.scala 96:25:@11801.4]
  assign _T_3052 = _T_3048 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@11810.4]
  assign _T_3045 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@11792.4 package.scala 96:25:@11793.4]
  assign _T_3053 = _T_3045 ? Mem1D_4_io_output : _T_3052; // @[Mux.scala 31:69:@11811.4]
  assign _T_3042 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@11784.4 package.scala 96:25:@11785.4]
  assign io_rPort_23_output_0 = _T_3042 ? Mem1D_io_output : _T_3053; // @[MemPrimitives.scala 148:13:@11813.4]
  assign io_rPort_22_output_0 = _T_3007 ? Mem1D_2_io_output : _T_3018; // @[MemPrimitives.scala 148:13:@11765.4]
  assign io_rPort_21_output_0 = _T_2972 ? Mem1D_3_io_output : _T_2983; // @[MemPrimitives.scala 148:13:@11717.4]
  assign io_rPort_20_output_0 = _T_2937 ? Mem1D_2_io_output : _T_2948; // @[MemPrimitives.scala 148:13:@11669.4]
  assign io_rPort_19_output_0 = _T_2902 ? Mem1D_2_io_output : _T_2913; // @[MemPrimitives.scala 148:13:@11621.4]
  assign io_rPort_18_output_0 = _T_2867 ? Mem1D_3_io_output : _T_2878; // @[MemPrimitives.scala 148:13:@11573.4]
  assign io_rPort_17_output_0 = _T_2832 ? Mem1D_3_io_output : _T_2843; // @[MemPrimitives.scala 148:13:@11525.4]
  assign io_rPort_16_output_0 = _T_2797 ? Mem1D_1_io_output : _T_2808; // @[MemPrimitives.scala 148:13:@11477.4]
  assign io_rPort_15_output_0 = _T_2762 ? Mem1D_1_io_output : _T_2773; // @[MemPrimitives.scala 148:13:@11429.4]
  assign io_rPort_14_output_0 = _T_2727 ? Mem1D_3_io_output : _T_2738; // @[MemPrimitives.scala 148:13:@11381.4]
  assign io_rPort_13_output_0 = _T_2692 ? Mem1D_2_io_output : _T_2703; // @[MemPrimitives.scala 148:13:@11333.4]
  assign io_rPort_12_output_0 = _T_2657 ? Mem1D_2_io_output : _T_2668; // @[MemPrimitives.scala 148:13:@11285.4]
  assign io_rPort_11_output_0 = _T_2622 ? Mem1D_3_io_output : _T_2633; // @[MemPrimitives.scala 148:13:@11237.4]
  assign io_rPort_10_output_0 = _T_2587 ? Mem1D_io_output : _T_2598; // @[MemPrimitives.scala 148:13:@11189.4]
  assign io_rPort_9_output_0 = _T_2552 ? Mem1D_2_io_output : _T_2563; // @[MemPrimitives.scala 148:13:@11141.4]
  assign io_rPort_8_output_0 = _T_2517 ? Mem1D_1_io_output : _T_2528; // @[MemPrimitives.scala 148:13:@11093.4]
  assign io_rPort_7_output_0 = _T_2482 ? Mem1D_3_io_output : _T_2493; // @[MemPrimitives.scala 148:13:@11045.4]
  assign io_rPort_6_output_0 = _T_2447 ? Mem1D_2_io_output : _T_2458; // @[MemPrimitives.scala 148:13:@10997.4]
  assign io_rPort_5_output_0 = _T_2412 ? Mem1D_3_io_output : _T_2423; // @[MemPrimitives.scala 148:13:@10949.4]
  assign io_rPort_4_output_0 = _T_2377 ? Mem1D_io_output : _T_2388; // @[MemPrimitives.scala 148:13:@10901.4]
  assign io_rPort_3_output_0 = _T_2342 ? Mem1D_2_io_output : _T_2353; // @[MemPrimitives.scala 148:13:@10853.4]
  assign io_rPort_2_output_0 = _T_2307 ? Mem1D_io_output : _T_2318; // @[MemPrimitives.scala 148:13:@10805.4]
  assign io_rPort_1_output_0 = _T_2272 ? Mem1D_3_io_output : _T_2283; // @[MemPrimitives.scala 148:13:@10757.4]
  assign io_rPort_0_output_0 = _T_2237 ? Mem1D_1_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@10709.4]
  assign Mem1D_clock = clock; // @[:@9239.4]
  assign Mem1D_reset = reset; // @[:@9240.4]
  assign Mem1D_io_r_ofs_0 = _T_1353[0]; // @[MemPrimitives.scala 127:28:@9803.4]
  assign Mem1D_io_r_backpressure = _T_1353[1]; // @[MemPrimitives.scala 128:32:@9804.4]
  assign Mem1D_io_w_ofs_0 = _T_1045[0]; // @[MemPrimitives.scala 94:28:@9508.4]
  assign Mem1D_io_w_data_0 = _T_1045[8:1]; // @[MemPrimitives.scala 95:29:@9509.4]
  assign Mem1D_io_w_en_0 = _T_1045[9]; // @[MemPrimitives.scala 96:27:@9510.4]
  assign Mem1D_1_clock = clock; // @[:@9255.4]
  assign Mem1D_1_reset = reset; // @[:@9256.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1391[0]; // @[MemPrimitives.scala 127:28:@9843.4]
  assign Mem1D_1_io_r_backpressure = _T_1391[1]; // @[MemPrimitives.scala 128:32:@9844.4]
  assign Mem1D_1_io_w_ofs_0 = _T_1063[0]; // @[MemPrimitives.scala 94:28:@9525.4]
  assign Mem1D_1_io_w_data_0 = _T_1063[8:1]; // @[MemPrimitives.scala 95:29:@9526.4]
  assign Mem1D_1_io_w_en_0 = _T_1063[9]; // @[MemPrimitives.scala 96:27:@9527.4]
  assign Mem1D_2_clock = clock; // @[:@9271.4]
  assign Mem1D_2_reset = reset; // @[:@9272.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1465[0]; // @[MemPrimitives.scala 127:28:@9915.4]
  assign Mem1D_2_io_r_backpressure = _T_1465[1]; // @[MemPrimitives.scala 128:32:@9916.4]
  assign Mem1D_2_io_w_ofs_0 = _T_1081[0]; // @[MemPrimitives.scala 94:28:@9542.4]
  assign Mem1D_2_io_w_data_0 = _T_1081[8:1]; // @[MemPrimitives.scala 95:29:@9543.4]
  assign Mem1D_2_io_w_en_0 = _T_1081[9]; // @[MemPrimitives.scala 96:27:@9544.4]
  assign Mem1D_3_clock = clock; // @[:@9287.4]
  assign Mem1D_3_reset = reset; // @[:@9288.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1539[0]; // @[MemPrimitives.scala 127:28:@9987.4]
  assign Mem1D_3_io_r_backpressure = _T_1539[1]; // @[MemPrimitives.scala 128:32:@9988.4]
  assign Mem1D_3_io_w_ofs_0 = _T_1099[0]; // @[MemPrimitives.scala 94:28:@9559.4]
  assign Mem1D_3_io_w_data_0 = _T_1099[8:1]; // @[MemPrimitives.scala 95:29:@9560.4]
  assign Mem1D_3_io_w_en_0 = _T_1099[9]; // @[MemPrimitives.scala 96:27:@9561.4]
  assign Mem1D_4_clock = clock; // @[:@9303.4]
  assign Mem1D_4_reset = reset; // @[:@9304.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1577[0]; // @[MemPrimitives.scala 127:28:@10027.4]
  assign Mem1D_4_io_r_backpressure = _T_1577[1]; // @[MemPrimitives.scala 128:32:@10028.4]
  assign Mem1D_4_io_w_ofs_0 = _T_1117[0]; // @[MemPrimitives.scala 94:28:@9576.4]
  assign Mem1D_4_io_w_data_0 = _T_1117[8:1]; // @[MemPrimitives.scala 95:29:@9577.4]
  assign Mem1D_4_io_w_en_0 = _T_1117[9]; // @[MemPrimitives.scala 96:27:@9578.4]
  assign Mem1D_5_clock = clock; // @[:@9319.4]
  assign Mem1D_5_reset = reset; // @[:@9320.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1615[0]; // @[MemPrimitives.scala 127:28:@10067.4]
  assign Mem1D_5_io_r_backpressure = _T_1615[1]; // @[MemPrimitives.scala 128:32:@10068.4]
  assign Mem1D_5_io_w_ofs_0 = _T_1135[0]; // @[MemPrimitives.scala 94:28:@9593.4]
  assign Mem1D_5_io_w_data_0 = _T_1135[8:1]; // @[MemPrimitives.scala 95:29:@9594.4]
  assign Mem1D_5_io_w_en_0 = _T_1135[9]; // @[MemPrimitives.scala 96:27:@9595.4]
  assign Mem1D_6_clock = clock; // @[:@9335.4]
  assign Mem1D_6_reset = reset; // @[:@9336.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1689[0]; // @[MemPrimitives.scala 127:28:@10139.4]
  assign Mem1D_6_io_r_backpressure = _T_1689[1]; // @[MemPrimitives.scala 128:32:@10140.4]
  assign Mem1D_6_io_w_ofs_0 = _T_1153[0]; // @[MemPrimitives.scala 94:28:@9610.4]
  assign Mem1D_6_io_w_data_0 = _T_1153[8:1]; // @[MemPrimitives.scala 95:29:@9611.4]
  assign Mem1D_6_io_w_en_0 = _T_1153[9]; // @[MemPrimitives.scala 96:27:@9612.4]
  assign Mem1D_7_clock = clock; // @[:@9351.4]
  assign Mem1D_7_reset = reset; // @[:@9352.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1763[0]; // @[MemPrimitives.scala 127:28:@10211.4]
  assign Mem1D_7_io_r_backpressure = _T_1763[1]; // @[MemPrimitives.scala 128:32:@10212.4]
  assign Mem1D_7_io_w_ofs_0 = _T_1171[0]; // @[MemPrimitives.scala 94:28:@9627.4]
  assign Mem1D_7_io_w_data_0 = _T_1171[8:1]; // @[MemPrimitives.scala 95:29:@9628.4]
  assign Mem1D_7_io_w_en_0 = _T_1171[9]; // @[MemPrimitives.scala 96:27:@9629.4]
  assign Mem1D_8_clock = clock; // @[:@9367.4]
  assign Mem1D_8_reset = reset; // @[:@9368.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1801[0]; // @[MemPrimitives.scala 127:28:@10251.4]
  assign Mem1D_8_io_r_backpressure = _T_1801[1]; // @[MemPrimitives.scala 128:32:@10252.4]
  assign Mem1D_8_io_w_ofs_0 = _T_1189[0]; // @[MemPrimitives.scala 94:28:@9644.4]
  assign Mem1D_8_io_w_data_0 = _T_1189[8:1]; // @[MemPrimitives.scala 95:29:@9645.4]
  assign Mem1D_8_io_w_en_0 = _T_1189[9]; // @[MemPrimitives.scala 96:27:@9646.4]
  assign Mem1D_9_clock = clock; // @[:@9383.4]
  assign Mem1D_9_reset = reset; // @[:@9384.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1839[0]; // @[MemPrimitives.scala 127:28:@10291.4]
  assign Mem1D_9_io_r_backpressure = _T_1839[1]; // @[MemPrimitives.scala 128:32:@10292.4]
  assign Mem1D_9_io_w_ofs_0 = _T_1207[0]; // @[MemPrimitives.scala 94:28:@9661.4]
  assign Mem1D_9_io_w_data_0 = _T_1207[8:1]; // @[MemPrimitives.scala 95:29:@9662.4]
  assign Mem1D_9_io_w_en_0 = _T_1207[9]; // @[MemPrimitives.scala 96:27:@9663.4]
  assign Mem1D_10_clock = clock; // @[:@9399.4]
  assign Mem1D_10_reset = reset; // @[:@9400.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1913[0]; // @[MemPrimitives.scala 127:28:@10363.4]
  assign Mem1D_10_io_r_backpressure = _T_1913[1]; // @[MemPrimitives.scala 128:32:@10364.4]
  assign Mem1D_10_io_w_ofs_0 = _T_1225[0]; // @[MemPrimitives.scala 94:28:@9678.4]
  assign Mem1D_10_io_w_data_0 = _T_1225[8:1]; // @[MemPrimitives.scala 95:29:@9679.4]
  assign Mem1D_10_io_w_en_0 = _T_1225[9]; // @[MemPrimitives.scala 96:27:@9680.4]
  assign Mem1D_11_clock = clock; // @[:@9415.4]
  assign Mem1D_11_reset = reset; // @[:@9416.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1987[0]; // @[MemPrimitives.scala 127:28:@10435.4]
  assign Mem1D_11_io_r_backpressure = _T_1987[1]; // @[MemPrimitives.scala 128:32:@10436.4]
  assign Mem1D_11_io_w_ofs_0 = _T_1243[0]; // @[MemPrimitives.scala 94:28:@9695.4]
  assign Mem1D_11_io_w_data_0 = _T_1243[8:1]; // @[MemPrimitives.scala 95:29:@9696.4]
  assign Mem1D_11_io_w_en_0 = _T_1243[9]; // @[MemPrimitives.scala 96:27:@9697.4]
  assign Mem1D_12_clock = clock; // @[:@9431.4]
  assign Mem1D_12_reset = reset; // @[:@9432.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2025[0]; // @[MemPrimitives.scala 127:28:@10475.4]
  assign Mem1D_12_io_r_backpressure = _T_2025[1]; // @[MemPrimitives.scala 128:32:@10476.4]
  assign Mem1D_12_io_w_ofs_0 = _T_1261[0]; // @[MemPrimitives.scala 94:28:@9712.4]
  assign Mem1D_12_io_w_data_0 = _T_1261[8:1]; // @[MemPrimitives.scala 95:29:@9713.4]
  assign Mem1D_12_io_w_en_0 = _T_1261[9]; // @[MemPrimitives.scala 96:27:@9714.4]
  assign Mem1D_13_clock = clock; // @[:@9447.4]
  assign Mem1D_13_reset = reset; // @[:@9448.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2063[0]; // @[MemPrimitives.scala 127:28:@10515.4]
  assign Mem1D_13_io_r_backpressure = _T_2063[1]; // @[MemPrimitives.scala 128:32:@10516.4]
  assign Mem1D_13_io_w_ofs_0 = _T_1279[0]; // @[MemPrimitives.scala 94:28:@9729.4]
  assign Mem1D_13_io_w_data_0 = _T_1279[8:1]; // @[MemPrimitives.scala 95:29:@9730.4]
  assign Mem1D_13_io_w_en_0 = _T_1279[9]; // @[MemPrimitives.scala 96:27:@9731.4]
  assign Mem1D_14_clock = clock; // @[:@9463.4]
  assign Mem1D_14_reset = reset; // @[:@9464.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2137[0]; // @[MemPrimitives.scala 127:28:@10587.4]
  assign Mem1D_14_io_r_backpressure = _T_2137[1]; // @[MemPrimitives.scala 128:32:@10588.4]
  assign Mem1D_14_io_w_ofs_0 = _T_1297[0]; // @[MemPrimitives.scala 94:28:@9746.4]
  assign Mem1D_14_io_w_data_0 = _T_1297[8:1]; // @[MemPrimitives.scala 95:29:@9747.4]
  assign Mem1D_14_io_w_en_0 = _T_1297[9]; // @[MemPrimitives.scala 96:27:@9748.4]
  assign Mem1D_15_clock = clock; // @[:@9479.4]
  assign Mem1D_15_reset = reset; // @[:@9480.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2211[0]; // @[MemPrimitives.scala 127:28:@10659.4]
  assign Mem1D_15_io_r_backpressure = _T_2211[1]; // @[MemPrimitives.scala 128:32:@10660.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1315[0]; // @[MemPrimitives.scala 94:28:@9763.4]
  assign Mem1D_15_io_w_data_0 = _T_1315[8:1]; // @[MemPrimitives.scala 95:29:@9764.4]
  assign Mem1D_15_io_w_en_0 = _T_1315[9]; // @[MemPrimitives.scala 96:27:@9765.4]
  assign StickySelects_clock = clock; // @[:@9779.4]
  assign StickySelects_reset = reset; // @[:@9780.4]
  assign StickySelects_io_ins_0 = io_rPort_2_en_0 & _T_1320; // @[MemPrimitives.scala 122:60:@9781.4]
  assign StickySelects_io_ins_1 = io_rPort_4_en_0 & _T_1325; // @[MemPrimitives.scala 122:60:@9782.4]
  assign StickySelects_io_ins_2 = io_rPort_10_en_0 & _T_1330; // @[MemPrimitives.scala 122:60:@9783.4]
  assign StickySelects_io_ins_3 = io_rPort_23_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@9784.4]
  assign StickySelects_1_clock = clock; // @[:@9819.4]
  assign StickySelects_1_reset = reset; // @[:@9820.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_1358; // @[MemPrimitives.scala 122:60:@9821.4]
  assign StickySelects_1_io_ins_1 = io_rPort_8_en_0 & _T_1363; // @[MemPrimitives.scala 122:60:@9822.4]
  assign StickySelects_1_io_ins_2 = io_rPort_15_en_0 & _T_1368; // @[MemPrimitives.scala 122:60:@9823.4]
  assign StickySelects_1_io_ins_3 = io_rPort_16_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@9824.4]
  assign StickySelects_2_clock = clock; // @[:@9871.4]
  assign StickySelects_2_reset = reset; // @[:@9872.4]
  assign StickySelects_2_io_ins_0 = io_rPort_3_en_0 & _T_1396; // @[MemPrimitives.scala 122:60:@9873.4]
  assign StickySelects_2_io_ins_1 = io_rPort_6_en_0 & _T_1401; // @[MemPrimitives.scala 122:60:@9874.4]
  assign StickySelects_2_io_ins_2 = io_rPort_9_en_0 & _T_1406; // @[MemPrimitives.scala 122:60:@9875.4]
  assign StickySelects_2_io_ins_3 = io_rPort_12_en_0 & _T_1411; // @[MemPrimitives.scala 122:60:@9876.4]
  assign StickySelects_2_io_ins_4 = io_rPort_13_en_0 & _T_1416; // @[MemPrimitives.scala 122:60:@9877.4]
  assign StickySelects_2_io_ins_5 = io_rPort_19_en_0 & _T_1421; // @[MemPrimitives.scala 122:60:@9878.4]
  assign StickySelects_2_io_ins_6 = io_rPort_20_en_0 & _T_1426; // @[MemPrimitives.scala 122:60:@9879.4]
  assign StickySelects_2_io_ins_7 = io_rPort_22_en_0 & _T_1431; // @[MemPrimitives.scala 122:60:@9880.4]
  assign StickySelects_3_clock = clock; // @[:@9943.4]
  assign StickySelects_3_reset = reset; // @[:@9944.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_1470; // @[MemPrimitives.scala 122:60:@9945.4]
  assign StickySelects_3_io_ins_1 = io_rPort_5_en_0 & _T_1475; // @[MemPrimitives.scala 122:60:@9946.4]
  assign StickySelects_3_io_ins_2 = io_rPort_7_en_0 & _T_1480; // @[MemPrimitives.scala 122:60:@9947.4]
  assign StickySelects_3_io_ins_3 = io_rPort_11_en_0 & _T_1485; // @[MemPrimitives.scala 122:60:@9948.4]
  assign StickySelects_3_io_ins_4 = io_rPort_14_en_0 & _T_1490; // @[MemPrimitives.scala 122:60:@9949.4]
  assign StickySelects_3_io_ins_5 = io_rPort_17_en_0 & _T_1495; // @[MemPrimitives.scala 122:60:@9950.4]
  assign StickySelects_3_io_ins_6 = io_rPort_18_en_0 & _T_1500; // @[MemPrimitives.scala 122:60:@9951.4]
  assign StickySelects_3_io_ins_7 = io_rPort_21_en_0 & _T_1505; // @[MemPrimitives.scala 122:60:@9952.4]
  assign StickySelects_4_clock = clock; // @[:@10003.4]
  assign StickySelects_4_reset = reset; // @[:@10004.4]
  assign StickySelects_4_io_ins_0 = io_rPort_2_en_0 & _T_1544; // @[MemPrimitives.scala 122:60:@10005.4]
  assign StickySelects_4_io_ins_1 = io_rPort_4_en_0 & _T_1549; // @[MemPrimitives.scala 122:60:@10006.4]
  assign StickySelects_4_io_ins_2 = io_rPort_10_en_0 & _T_1554; // @[MemPrimitives.scala 122:60:@10007.4]
  assign StickySelects_4_io_ins_3 = io_rPort_23_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@10008.4]
  assign StickySelects_5_clock = clock; // @[:@10043.4]
  assign StickySelects_5_reset = reset; // @[:@10044.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_1582; // @[MemPrimitives.scala 122:60:@10045.4]
  assign StickySelects_5_io_ins_1 = io_rPort_8_en_0 & _T_1587; // @[MemPrimitives.scala 122:60:@10046.4]
  assign StickySelects_5_io_ins_2 = io_rPort_15_en_0 & _T_1592; // @[MemPrimitives.scala 122:60:@10047.4]
  assign StickySelects_5_io_ins_3 = io_rPort_16_en_0 & _T_1597; // @[MemPrimitives.scala 122:60:@10048.4]
  assign StickySelects_6_clock = clock; // @[:@10095.4]
  assign StickySelects_6_reset = reset; // @[:@10096.4]
  assign StickySelects_6_io_ins_0 = io_rPort_3_en_0 & _T_1620; // @[MemPrimitives.scala 122:60:@10097.4]
  assign StickySelects_6_io_ins_1 = io_rPort_6_en_0 & _T_1625; // @[MemPrimitives.scala 122:60:@10098.4]
  assign StickySelects_6_io_ins_2 = io_rPort_9_en_0 & _T_1630; // @[MemPrimitives.scala 122:60:@10099.4]
  assign StickySelects_6_io_ins_3 = io_rPort_12_en_0 & _T_1635; // @[MemPrimitives.scala 122:60:@10100.4]
  assign StickySelects_6_io_ins_4 = io_rPort_13_en_0 & _T_1640; // @[MemPrimitives.scala 122:60:@10101.4]
  assign StickySelects_6_io_ins_5 = io_rPort_19_en_0 & _T_1645; // @[MemPrimitives.scala 122:60:@10102.4]
  assign StickySelects_6_io_ins_6 = io_rPort_20_en_0 & _T_1650; // @[MemPrimitives.scala 122:60:@10103.4]
  assign StickySelects_6_io_ins_7 = io_rPort_22_en_0 & _T_1655; // @[MemPrimitives.scala 122:60:@10104.4]
  assign StickySelects_7_clock = clock; // @[:@10167.4]
  assign StickySelects_7_reset = reset; // @[:@10168.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1694; // @[MemPrimitives.scala 122:60:@10169.4]
  assign StickySelects_7_io_ins_1 = io_rPort_5_en_0 & _T_1699; // @[MemPrimitives.scala 122:60:@10170.4]
  assign StickySelects_7_io_ins_2 = io_rPort_7_en_0 & _T_1704; // @[MemPrimitives.scala 122:60:@10171.4]
  assign StickySelects_7_io_ins_3 = io_rPort_11_en_0 & _T_1709; // @[MemPrimitives.scala 122:60:@10172.4]
  assign StickySelects_7_io_ins_4 = io_rPort_14_en_0 & _T_1714; // @[MemPrimitives.scala 122:60:@10173.4]
  assign StickySelects_7_io_ins_5 = io_rPort_17_en_0 & _T_1719; // @[MemPrimitives.scala 122:60:@10174.4]
  assign StickySelects_7_io_ins_6 = io_rPort_18_en_0 & _T_1724; // @[MemPrimitives.scala 122:60:@10175.4]
  assign StickySelects_7_io_ins_7 = io_rPort_21_en_0 & _T_1729; // @[MemPrimitives.scala 122:60:@10176.4]
  assign StickySelects_8_clock = clock; // @[:@10227.4]
  assign StickySelects_8_reset = reset; // @[:@10228.4]
  assign StickySelects_8_io_ins_0 = io_rPort_2_en_0 & _T_1768; // @[MemPrimitives.scala 122:60:@10229.4]
  assign StickySelects_8_io_ins_1 = io_rPort_4_en_0 & _T_1773; // @[MemPrimitives.scala 122:60:@10230.4]
  assign StickySelects_8_io_ins_2 = io_rPort_10_en_0 & _T_1778; // @[MemPrimitives.scala 122:60:@10231.4]
  assign StickySelects_8_io_ins_3 = io_rPort_23_en_0 & _T_1783; // @[MemPrimitives.scala 122:60:@10232.4]
  assign StickySelects_9_clock = clock; // @[:@10267.4]
  assign StickySelects_9_reset = reset; // @[:@10268.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1806; // @[MemPrimitives.scala 122:60:@10269.4]
  assign StickySelects_9_io_ins_1 = io_rPort_8_en_0 & _T_1811; // @[MemPrimitives.scala 122:60:@10270.4]
  assign StickySelects_9_io_ins_2 = io_rPort_15_en_0 & _T_1816; // @[MemPrimitives.scala 122:60:@10271.4]
  assign StickySelects_9_io_ins_3 = io_rPort_16_en_0 & _T_1821; // @[MemPrimitives.scala 122:60:@10272.4]
  assign StickySelects_10_clock = clock; // @[:@10319.4]
  assign StickySelects_10_reset = reset; // @[:@10320.4]
  assign StickySelects_10_io_ins_0 = io_rPort_3_en_0 & _T_1844; // @[MemPrimitives.scala 122:60:@10321.4]
  assign StickySelects_10_io_ins_1 = io_rPort_6_en_0 & _T_1849; // @[MemPrimitives.scala 122:60:@10322.4]
  assign StickySelects_10_io_ins_2 = io_rPort_9_en_0 & _T_1854; // @[MemPrimitives.scala 122:60:@10323.4]
  assign StickySelects_10_io_ins_3 = io_rPort_12_en_0 & _T_1859; // @[MemPrimitives.scala 122:60:@10324.4]
  assign StickySelects_10_io_ins_4 = io_rPort_13_en_0 & _T_1864; // @[MemPrimitives.scala 122:60:@10325.4]
  assign StickySelects_10_io_ins_5 = io_rPort_19_en_0 & _T_1869; // @[MemPrimitives.scala 122:60:@10326.4]
  assign StickySelects_10_io_ins_6 = io_rPort_20_en_0 & _T_1874; // @[MemPrimitives.scala 122:60:@10327.4]
  assign StickySelects_10_io_ins_7 = io_rPort_22_en_0 & _T_1879; // @[MemPrimitives.scala 122:60:@10328.4]
  assign StickySelects_11_clock = clock; // @[:@10391.4]
  assign StickySelects_11_reset = reset; // @[:@10392.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1918; // @[MemPrimitives.scala 122:60:@10393.4]
  assign StickySelects_11_io_ins_1 = io_rPort_5_en_0 & _T_1923; // @[MemPrimitives.scala 122:60:@10394.4]
  assign StickySelects_11_io_ins_2 = io_rPort_7_en_0 & _T_1928; // @[MemPrimitives.scala 122:60:@10395.4]
  assign StickySelects_11_io_ins_3 = io_rPort_11_en_0 & _T_1933; // @[MemPrimitives.scala 122:60:@10396.4]
  assign StickySelects_11_io_ins_4 = io_rPort_14_en_0 & _T_1938; // @[MemPrimitives.scala 122:60:@10397.4]
  assign StickySelects_11_io_ins_5 = io_rPort_17_en_0 & _T_1943; // @[MemPrimitives.scala 122:60:@10398.4]
  assign StickySelects_11_io_ins_6 = io_rPort_18_en_0 & _T_1948; // @[MemPrimitives.scala 122:60:@10399.4]
  assign StickySelects_11_io_ins_7 = io_rPort_21_en_0 & _T_1953; // @[MemPrimitives.scala 122:60:@10400.4]
  assign StickySelects_12_clock = clock; // @[:@10451.4]
  assign StickySelects_12_reset = reset; // @[:@10452.4]
  assign StickySelects_12_io_ins_0 = io_rPort_2_en_0 & _T_1992; // @[MemPrimitives.scala 122:60:@10453.4]
  assign StickySelects_12_io_ins_1 = io_rPort_4_en_0 & _T_1997; // @[MemPrimitives.scala 122:60:@10454.4]
  assign StickySelects_12_io_ins_2 = io_rPort_10_en_0 & _T_2002; // @[MemPrimitives.scala 122:60:@10455.4]
  assign StickySelects_12_io_ins_3 = io_rPort_23_en_0 & _T_2007; // @[MemPrimitives.scala 122:60:@10456.4]
  assign StickySelects_13_clock = clock; // @[:@10491.4]
  assign StickySelects_13_reset = reset; // @[:@10492.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_2030; // @[MemPrimitives.scala 122:60:@10493.4]
  assign StickySelects_13_io_ins_1 = io_rPort_8_en_0 & _T_2035; // @[MemPrimitives.scala 122:60:@10494.4]
  assign StickySelects_13_io_ins_2 = io_rPort_15_en_0 & _T_2040; // @[MemPrimitives.scala 122:60:@10495.4]
  assign StickySelects_13_io_ins_3 = io_rPort_16_en_0 & _T_2045; // @[MemPrimitives.scala 122:60:@10496.4]
  assign StickySelects_14_clock = clock; // @[:@10543.4]
  assign StickySelects_14_reset = reset; // @[:@10544.4]
  assign StickySelects_14_io_ins_0 = io_rPort_3_en_0 & _T_2068; // @[MemPrimitives.scala 122:60:@10545.4]
  assign StickySelects_14_io_ins_1 = io_rPort_6_en_0 & _T_2073; // @[MemPrimitives.scala 122:60:@10546.4]
  assign StickySelects_14_io_ins_2 = io_rPort_9_en_0 & _T_2078; // @[MemPrimitives.scala 122:60:@10547.4]
  assign StickySelects_14_io_ins_3 = io_rPort_12_en_0 & _T_2083; // @[MemPrimitives.scala 122:60:@10548.4]
  assign StickySelects_14_io_ins_4 = io_rPort_13_en_0 & _T_2088; // @[MemPrimitives.scala 122:60:@10549.4]
  assign StickySelects_14_io_ins_5 = io_rPort_19_en_0 & _T_2093; // @[MemPrimitives.scala 122:60:@10550.4]
  assign StickySelects_14_io_ins_6 = io_rPort_20_en_0 & _T_2098; // @[MemPrimitives.scala 122:60:@10551.4]
  assign StickySelects_14_io_ins_7 = io_rPort_22_en_0 & _T_2103; // @[MemPrimitives.scala 122:60:@10552.4]
  assign StickySelects_15_clock = clock; // @[:@10615.4]
  assign StickySelects_15_reset = reset; // @[:@10616.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_2142; // @[MemPrimitives.scala 122:60:@10617.4]
  assign StickySelects_15_io_ins_1 = io_rPort_5_en_0 & _T_2147; // @[MemPrimitives.scala 122:60:@10618.4]
  assign StickySelects_15_io_ins_2 = io_rPort_7_en_0 & _T_2152; // @[MemPrimitives.scala 122:60:@10619.4]
  assign StickySelects_15_io_ins_3 = io_rPort_11_en_0 & _T_2157; // @[MemPrimitives.scala 122:60:@10620.4]
  assign StickySelects_15_io_ins_4 = io_rPort_14_en_0 & _T_2162; // @[MemPrimitives.scala 122:60:@10621.4]
  assign StickySelects_15_io_ins_5 = io_rPort_17_en_0 & _T_2167; // @[MemPrimitives.scala 122:60:@10622.4]
  assign StickySelects_15_io_ins_6 = io_rPort_18_en_0 & _T_2172; // @[MemPrimitives.scala 122:60:@10623.4]
  assign StickySelects_15_io_ins_7 = io_rPort_21_en_0 & _T_2177; // @[MemPrimitives.scala 122:60:@10624.4]
  assign RetimeWrapper_clock = clock; // @[:@10676.4]
  assign RetimeWrapper_reset = reset; // @[:@10677.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10679.4]
  assign RetimeWrapper_io_in = _T_1358 & io_rPort_0_en_0; // @[package.scala 94:16:@10678.4]
  assign RetimeWrapper_1_clock = clock; // @[:@10684.4]
  assign RetimeWrapper_1_reset = reset; // @[:@10685.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10687.4]
  assign RetimeWrapper_1_io_in = _T_1582 & io_rPort_0_en_0; // @[package.scala 94:16:@10686.4]
  assign RetimeWrapper_2_clock = clock; // @[:@10692.4]
  assign RetimeWrapper_2_reset = reset; // @[:@10693.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10695.4]
  assign RetimeWrapper_2_io_in = _T_1806 & io_rPort_0_en_0; // @[package.scala 94:16:@10694.4]
  assign RetimeWrapper_3_clock = clock; // @[:@10700.4]
  assign RetimeWrapper_3_reset = reset; // @[:@10701.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@10703.4]
  assign RetimeWrapper_3_io_in = _T_2030 & io_rPort_0_en_0; // @[package.scala 94:16:@10702.4]
  assign RetimeWrapper_4_clock = clock; // @[:@10724.4]
  assign RetimeWrapper_4_reset = reset; // @[:@10725.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10727.4]
  assign RetimeWrapper_4_io_in = _T_1470 & io_rPort_1_en_0; // @[package.scala 94:16:@10726.4]
  assign RetimeWrapper_5_clock = clock; // @[:@10732.4]
  assign RetimeWrapper_5_reset = reset; // @[:@10733.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10735.4]
  assign RetimeWrapper_5_io_in = _T_1694 & io_rPort_1_en_0; // @[package.scala 94:16:@10734.4]
  assign RetimeWrapper_6_clock = clock; // @[:@10740.4]
  assign RetimeWrapper_6_reset = reset; // @[:@10741.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10743.4]
  assign RetimeWrapper_6_io_in = _T_1918 & io_rPort_1_en_0; // @[package.scala 94:16:@10742.4]
  assign RetimeWrapper_7_clock = clock; // @[:@10748.4]
  assign RetimeWrapper_7_reset = reset; // @[:@10749.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@10751.4]
  assign RetimeWrapper_7_io_in = _T_2142 & io_rPort_1_en_0; // @[package.scala 94:16:@10750.4]
  assign RetimeWrapper_8_clock = clock; // @[:@10772.4]
  assign RetimeWrapper_8_reset = reset; // @[:@10773.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10775.4]
  assign RetimeWrapper_8_io_in = _T_1320 & io_rPort_2_en_0; // @[package.scala 94:16:@10774.4]
  assign RetimeWrapper_9_clock = clock; // @[:@10780.4]
  assign RetimeWrapper_9_reset = reset; // @[:@10781.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10783.4]
  assign RetimeWrapper_9_io_in = _T_1544 & io_rPort_2_en_0; // @[package.scala 94:16:@10782.4]
  assign RetimeWrapper_10_clock = clock; // @[:@10788.4]
  assign RetimeWrapper_10_reset = reset; // @[:@10789.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10791.4]
  assign RetimeWrapper_10_io_in = _T_1768 & io_rPort_2_en_0; // @[package.scala 94:16:@10790.4]
  assign RetimeWrapper_11_clock = clock; // @[:@10796.4]
  assign RetimeWrapper_11_reset = reset; // @[:@10797.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@10799.4]
  assign RetimeWrapper_11_io_in = _T_1992 & io_rPort_2_en_0; // @[package.scala 94:16:@10798.4]
  assign RetimeWrapper_12_clock = clock; // @[:@10820.4]
  assign RetimeWrapper_12_reset = reset; // @[:@10821.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10823.4]
  assign RetimeWrapper_12_io_in = _T_1396 & io_rPort_3_en_0; // @[package.scala 94:16:@10822.4]
  assign RetimeWrapper_13_clock = clock; // @[:@10828.4]
  assign RetimeWrapper_13_reset = reset; // @[:@10829.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10831.4]
  assign RetimeWrapper_13_io_in = _T_1620 & io_rPort_3_en_0; // @[package.scala 94:16:@10830.4]
  assign RetimeWrapper_14_clock = clock; // @[:@10836.4]
  assign RetimeWrapper_14_reset = reset; // @[:@10837.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10839.4]
  assign RetimeWrapper_14_io_in = _T_1844 & io_rPort_3_en_0; // @[package.scala 94:16:@10838.4]
  assign RetimeWrapper_15_clock = clock; // @[:@10844.4]
  assign RetimeWrapper_15_reset = reset; // @[:@10845.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@10847.4]
  assign RetimeWrapper_15_io_in = _T_2068 & io_rPort_3_en_0; // @[package.scala 94:16:@10846.4]
  assign RetimeWrapper_16_clock = clock; // @[:@10868.4]
  assign RetimeWrapper_16_reset = reset; // @[:@10869.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10871.4]
  assign RetimeWrapper_16_io_in = _T_1325 & io_rPort_4_en_0; // @[package.scala 94:16:@10870.4]
  assign RetimeWrapper_17_clock = clock; // @[:@10876.4]
  assign RetimeWrapper_17_reset = reset; // @[:@10877.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10879.4]
  assign RetimeWrapper_17_io_in = _T_1549 & io_rPort_4_en_0; // @[package.scala 94:16:@10878.4]
  assign RetimeWrapper_18_clock = clock; // @[:@10884.4]
  assign RetimeWrapper_18_reset = reset; // @[:@10885.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10887.4]
  assign RetimeWrapper_18_io_in = _T_1773 & io_rPort_4_en_0; // @[package.scala 94:16:@10886.4]
  assign RetimeWrapper_19_clock = clock; // @[:@10892.4]
  assign RetimeWrapper_19_reset = reset; // @[:@10893.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@10895.4]
  assign RetimeWrapper_19_io_in = _T_1997 & io_rPort_4_en_0; // @[package.scala 94:16:@10894.4]
  assign RetimeWrapper_20_clock = clock; // @[:@10916.4]
  assign RetimeWrapper_20_reset = reset; // @[:@10917.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10919.4]
  assign RetimeWrapper_20_io_in = _T_1475 & io_rPort_5_en_0; // @[package.scala 94:16:@10918.4]
  assign RetimeWrapper_21_clock = clock; // @[:@10924.4]
  assign RetimeWrapper_21_reset = reset; // @[:@10925.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10927.4]
  assign RetimeWrapper_21_io_in = _T_1699 & io_rPort_5_en_0; // @[package.scala 94:16:@10926.4]
  assign RetimeWrapper_22_clock = clock; // @[:@10932.4]
  assign RetimeWrapper_22_reset = reset; // @[:@10933.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10935.4]
  assign RetimeWrapper_22_io_in = _T_1923 & io_rPort_5_en_0; // @[package.scala 94:16:@10934.4]
  assign RetimeWrapper_23_clock = clock; // @[:@10940.4]
  assign RetimeWrapper_23_reset = reset; // @[:@10941.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@10943.4]
  assign RetimeWrapper_23_io_in = _T_2147 & io_rPort_5_en_0; // @[package.scala 94:16:@10942.4]
  assign RetimeWrapper_24_clock = clock; // @[:@10964.4]
  assign RetimeWrapper_24_reset = reset; // @[:@10965.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10967.4]
  assign RetimeWrapper_24_io_in = _T_1401 & io_rPort_6_en_0; // @[package.scala 94:16:@10966.4]
  assign RetimeWrapper_25_clock = clock; // @[:@10972.4]
  assign RetimeWrapper_25_reset = reset; // @[:@10973.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10975.4]
  assign RetimeWrapper_25_io_in = _T_1625 & io_rPort_6_en_0; // @[package.scala 94:16:@10974.4]
  assign RetimeWrapper_26_clock = clock; // @[:@10980.4]
  assign RetimeWrapper_26_reset = reset; // @[:@10981.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10983.4]
  assign RetimeWrapper_26_io_in = _T_1849 & io_rPort_6_en_0; // @[package.scala 94:16:@10982.4]
  assign RetimeWrapper_27_clock = clock; // @[:@10988.4]
  assign RetimeWrapper_27_reset = reset; // @[:@10989.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@10991.4]
  assign RetimeWrapper_27_io_in = _T_2073 & io_rPort_6_en_0; // @[package.scala 94:16:@10990.4]
  assign RetimeWrapper_28_clock = clock; // @[:@11012.4]
  assign RetimeWrapper_28_reset = reset; // @[:@11013.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11015.4]
  assign RetimeWrapper_28_io_in = _T_1480 & io_rPort_7_en_0; // @[package.scala 94:16:@11014.4]
  assign RetimeWrapper_29_clock = clock; // @[:@11020.4]
  assign RetimeWrapper_29_reset = reset; // @[:@11021.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11023.4]
  assign RetimeWrapper_29_io_in = _T_1704 & io_rPort_7_en_0; // @[package.scala 94:16:@11022.4]
  assign RetimeWrapper_30_clock = clock; // @[:@11028.4]
  assign RetimeWrapper_30_reset = reset; // @[:@11029.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11031.4]
  assign RetimeWrapper_30_io_in = _T_1928 & io_rPort_7_en_0; // @[package.scala 94:16:@11030.4]
  assign RetimeWrapper_31_clock = clock; // @[:@11036.4]
  assign RetimeWrapper_31_reset = reset; // @[:@11037.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@11039.4]
  assign RetimeWrapper_31_io_in = _T_2152 & io_rPort_7_en_0; // @[package.scala 94:16:@11038.4]
  assign RetimeWrapper_32_clock = clock; // @[:@11060.4]
  assign RetimeWrapper_32_reset = reset; // @[:@11061.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11063.4]
  assign RetimeWrapper_32_io_in = _T_1363 & io_rPort_8_en_0; // @[package.scala 94:16:@11062.4]
  assign RetimeWrapper_33_clock = clock; // @[:@11068.4]
  assign RetimeWrapper_33_reset = reset; // @[:@11069.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11071.4]
  assign RetimeWrapper_33_io_in = _T_1587 & io_rPort_8_en_0; // @[package.scala 94:16:@11070.4]
  assign RetimeWrapper_34_clock = clock; // @[:@11076.4]
  assign RetimeWrapper_34_reset = reset; // @[:@11077.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11079.4]
  assign RetimeWrapper_34_io_in = _T_1811 & io_rPort_8_en_0; // @[package.scala 94:16:@11078.4]
  assign RetimeWrapper_35_clock = clock; // @[:@11084.4]
  assign RetimeWrapper_35_reset = reset; // @[:@11085.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@11087.4]
  assign RetimeWrapper_35_io_in = _T_2035 & io_rPort_8_en_0; // @[package.scala 94:16:@11086.4]
  assign RetimeWrapper_36_clock = clock; // @[:@11108.4]
  assign RetimeWrapper_36_reset = reset; // @[:@11109.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11111.4]
  assign RetimeWrapper_36_io_in = _T_1406 & io_rPort_9_en_0; // @[package.scala 94:16:@11110.4]
  assign RetimeWrapper_37_clock = clock; // @[:@11116.4]
  assign RetimeWrapper_37_reset = reset; // @[:@11117.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11119.4]
  assign RetimeWrapper_37_io_in = _T_1630 & io_rPort_9_en_0; // @[package.scala 94:16:@11118.4]
  assign RetimeWrapper_38_clock = clock; // @[:@11124.4]
  assign RetimeWrapper_38_reset = reset; // @[:@11125.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11127.4]
  assign RetimeWrapper_38_io_in = _T_1854 & io_rPort_9_en_0; // @[package.scala 94:16:@11126.4]
  assign RetimeWrapper_39_clock = clock; // @[:@11132.4]
  assign RetimeWrapper_39_reset = reset; // @[:@11133.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@11135.4]
  assign RetimeWrapper_39_io_in = _T_2078 & io_rPort_9_en_0; // @[package.scala 94:16:@11134.4]
  assign RetimeWrapper_40_clock = clock; // @[:@11156.4]
  assign RetimeWrapper_40_reset = reset; // @[:@11157.4]
  assign RetimeWrapper_40_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11159.4]
  assign RetimeWrapper_40_io_in = _T_1330 & io_rPort_10_en_0; // @[package.scala 94:16:@11158.4]
  assign RetimeWrapper_41_clock = clock; // @[:@11164.4]
  assign RetimeWrapper_41_reset = reset; // @[:@11165.4]
  assign RetimeWrapper_41_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11167.4]
  assign RetimeWrapper_41_io_in = _T_1554 & io_rPort_10_en_0; // @[package.scala 94:16:@11166.4]
  assign RetimeWrapper_42_clock = clock; // @[:@11172.4]
  assign RetimeWrapper_42_reset = reset; // @[:@11173.4]
  assign RetimeWrapper_42_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11175.4]
  assign RetimeWrapper_42_io_in = _T_1778 & io_rPort_10_en_0; // @[package.scala 94:16:@11174.4]
  assign RetimeWrapper_43_clock = clock; // @[:@11180.4]
  assign RetimeWrapper_43_reset = reset; // @[:@11181.4]
  assign RetimeWrapper_43_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@11183.4]
  assign RetimeWrapper_43_io_in = _T_2002 & io_rPort_10_en_0; // @[package.scala 94:16:@11182.4]
  assign RetimeWrapper_44_clock = clock; // @[:@11204.4]
  assign RetimeWrapper_44_reset = reset; // @[:@11205.4]
  assign RetimeWrapper_44_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11207.4]
  assign RetimeWrapper_44_io_in = _T_1485 & io_rPort_11_en_0; // @[package.scala 94:16:@11206.4]
  assign RetimeWrapper_45_clock = clock; // @[:@11212.4]
  assign RetimeWrapper_45_reset = reset; // @[:@11213.4]
  assign RetimeWrapper_45_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11215.4]
  assign RetimeWrapper_45_io_in = _T_1709 & io_rPort_11_en_0; // @[package.scala 94:16:@11214.4]
  assign RetimeWrapper_46_clock = clock; // @[:@11220.4]
  assign RetimeWrapper_46_reset = reset; // @[:@11221.4]
  assign RetimeWrapper_46_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11223.4]
  assign RetimeWrapper_46_io_in = _T_1933 & io_rPort_11_en_0; // @[package.scala 94:16:@11222.4]
  assign RetimeWrapper_47_clock = clock; // @[:@11228.4]
  assign RetimeWrapper_47_reset = reset; // @[:@11229.4]
  assign RetimeWrapper_47_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@11231.4]
  assign RetimeWrapper_47_io_in = _T_2157 & io_rPort_11_en_0; // @[package.scala 94:16:@11230.4]
  assign RetimeWrapper_48_clock = clock; // @[:@11252.4]
  assign RetimeWrapper_48_reset = reset; // @[:@11253.4]
  assign RetimeWrapper_48_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11255.4]
  assign RetimeWrapper_48_io_in = _T_1411 & io_rPort_12_en_0; // @[package.scala 94:16:@11254.4]
  assign RetimeWrapper_49_clock = clock; // @[:@11260.4]
  assign RetimeWrapper_49_reset = reset; // @[:@11261.4]
  assign RetimeWrapper_49_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11263.4]
  assign RetimeWrapper_49_io_in = _T_1635 & io_rPort_12_en_0; // @[package.scala 94:16:@11262.4]
  assign RetimeWrapper_50_clock = clock; // @[:@11268.4]
  assign RetimeWrapper_50_reset = reset; // @[:@11269.4]
  assign RetimeWrapper_50_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11271.4]
  assign RetimeWrapper_50_io_in = _T_1859 & io_rPort_12_en_0; // @[package.scala 94:16:@11270.4]
  assign RetimeWrapper_51_clock = clock; // @[:@11276.4]
  assign RetimeWrapper_51_reset = reset; // @[:@11277.4]
  assign RetimeWrapper_51_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@11279.4]
  assign RetimeWrapper_51_io_in = _T_2083 & io_rPort_12_en_0; // @[package.scala 94:16:@11278.4]
  assign RetimeWrapper_52_clock = clock; // @[:@11300.4]
  assign RetimeWrapper_52_reset = reset; // @[:@11301.4]
  assign RetimeWrapper_52_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11303.4]
  assign RetimeWrapper_52_io_in = _T_1416 & io_rPort_13_en_0; // @[package.scala 94:16:@11302.4]
  assign RetimeWrapper_53_clock = clock; // @[:@11308.4]
  assign RetimeWrapper_53_reset = reset; // @[:@11309.4]
  assign RetimeWrapper_53_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11311.4]
  assign RetimeWrapper_53_io_in = _T_1640 & io_rPort_13_en_0; // @[package.scala 94:16:@11310.4]
  assign RetimeWrapper_54_clock = clock; // @[:@11316.4]
  assign RetimeWrapper_54_reset = reset; // @[:@11317.4]
  assign RetimeWrapper_54_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11319.4]
  assign RetimeWrapper_54_io_in = _T_1864 & io_rPort_13_en_0; // @[package.scala 94:16:@11318.4]
  assign RetimeWrapper_55_clock = clock; // @[:@11324.4]
  assign RetimeWrapper_55_reset = reset; // @[:@11325.4]
  assign RetimeWrapper_55_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@11327.4]
  assign RetimeWrapper_55_io_in = _T_2088 & io_rPort_13_en_0; // @[package.scala 94:16:@11326.4]
  assign RetimeWrapper_56_clock = clock; // @[:@11348.4]
  assign RetimeWrapper_56_reset = reset; // @[:@11349.4]
  assign RetimeWrapper_56_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11351.4]
  assign RetimeWrapper_56_io_in = _T_1490 & io_rPort_14_en_0; // @[package.scala 94:16:@11350.4]
  assign RetimeWrapper_57_clock = clock; // @[:@11356.4]
  assign RetimeWrapper_57_reset = reset; // @[:@11357.4]
  assign RetimeWrapper_57_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11359.4]
  assign RetimeWrapper_57_io_in = _T_1714 & io_rPort_14_en_0; // @[package.scala 94:16:@11358.4]
  assign RetimeWrapper_58_clock = clock; // @[:@11364.4]
  assign RetimeWrapper_58_reset = reset; // @[:@11365.4]
  assign RetimeWrapper_58_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11367.4]
  assign RetimeWrapper_58_io_in = _T_1938 & io_rPort_14_en_0; // @[package.scala 94:16:@11366.4]
  assign RetimeWrapper_59_clock = clock; // @[:@11372.4]
  assign RetimeWrapper_59_reset = reset; // @[:@11373.4]
  assign RetimeWrapper_59_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@11375.4]
  assign RetimeWrapper_59_io_in = _T_2162 & io_rPort_14_en_0; // @[package.scala 94:16:@11374.4]
  assign RetimeWrapper_60_clock = clock; // @[:@11396.4]
  assign RetimeWrapper_60_reset = reset; // @[:@11397.4]
  assign RetimeWrapper_60_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11399.4]
  assign RetimeWrapper_60_io_in = _T_1368 & io_rPort_15_en_0; // @[package.scala 94:16:@11398.4]
  assign RetimeWrapper_61_clock = clock; // @[:@11404.4]
  assign RetimeWrapper_61_reset = reset; // @[:@11405.4]
  assign RetimeWrapper_61_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11407.4]
  assign RetimeWrapper_61_io_in = _T_1592 & io_rPort_15_en_0; // @[package.scala 94:16:@11406.4]
  assign RetimeWrapper_62_clock = clock; // @[:@11412.4]
  assign RetimeWrapper_62_reset = reset; // @[:@11413.4]
  assign RetimeWrapper_62_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11415.4]
  assign RetimeWrapper_62_io_in = _T_1816 & io_rPort_15_en_0; // @[package.scala 94:16:@11414.4]
  assign RetimeWrapper_63_clock = clock; // @[:@11420.4]
  assign RetimeWrapper_63_reset = reset; // @[:@11421.4]
  assign RetimeWrapper_63_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@11423.4]
  assign RetimeWrapper_63_io_in = _T_2040 & io_rPort_15_en_0; // @[package.scala 94:16:@11422.4]
  assign RetimeWrapper_64_clock = clock; // @[:@11444.4]
  assign RetimeWrapper_64_reset = reset; // @[:@11445.4]
  assign RetimeWrapper_64_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11447.4]
  assign RetimeWrapper_64_io_in = _T_1373 & io_rPort_16_en_0; // @[package.scala 94:16:@11446.4]
  assign RetimeWrapper_65_clock = clock; // @[:@11452.4]
  assign RetimeWrapper_65_reset = reset; // @[:@11453.4]
  assign RetimeWrapper_65_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11455.4]
  assign RetimeWrapper_65_io_in = _T_1597 & io_rPort_16_en_0; // @[package.scala 94:16:@11454.4]
  assign RetimeWrapper_66_clock = clock; // @[:@11460.4]
  assign RetimeWrapper_66_reset = reset; // @[:@11461.4]
  assign RetimeWrapper_66_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11463.4]
  assign RetimeWrapper_66_io_in = _T_1821 & io_rPort_16_en_0; // @[package.scala 94:16:@11462.4]
  assign RetimeWrapper_67_clock = clock; // @[:@11468.4]
  assign RetimeWrapper_67_reset = reset; // @[:@11469.4]
  assign RetimeWrapper_67_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@11471.4]
  assign RetimeWrapper_67_io_in = _T_2045 & io_rPort_16_en_0; // @[package.scala 94:16:@11470.4]
  assign RetimeWrapper_68_clock = clock; // @[:@11492.4]
  assign RetimeWrapper_68_reset = reset; // @[:@11493.4]
  assign RetimeWrapper_68_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11495.4]
  assign RetimeWrapper_68_io_in = _T_1495 & io_rPort_17_en_0; // @[package.scala 94:16:@11494.4]
  assign RetimeWrapper_69_clock = clock; // @[:@11500.4]
  assign RetimeWrapper_69_reset = reset; // @[:@11501.4]
  assign RetimeWrapper_69_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11503.4]
  assign RetimeWrapper_69_io_in = _T_1719 & io_rPort_17_en_0; // @[package.scala 94:16:@11502.4]
  assign RetimeWrapper_70_clock = clock; // @[:@11508.4]
  assign RetimeWrapper_70_reset = reset; // @[:@11509.4]
  assign RetimeWrapper_70_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11511.4]
  assign RetimeWrapper_70_io_in = _T_1943 & io_rPort_17_en_0; // @[package.scala 94:16:@11510.4]
  assign RetimeWrapper_71_clock = clock; // @[:@11516.4]
  assign RetimeWrapper_71_reset = reset; // @[:@11517.4]
  assign RetimeWrapper_71_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@11519.4]
  assign RetimeWrapper_71_io_in = _T_2167 & io_rPort_17_en_0; // @[package.scala 94:16:@11518.4]
  assign RetimeWrapper_72_clock = clock; // @[:@11540.4]
  assign RetimeWrapper_72_reset = reset; // @[:@11541.4]
  assign RetimeWrapper_72_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11543.4]
  assign RetimeWrapper_72_io_in = _T_1500 & io_rPort_18_en_0; // @[package.scala 94:16:@11542.4]
  assign RetimeWrapper_73_clock = clock; // @[:@11548.4]
  assign RetimeWrapper_73_reset = reset; // @[:@11549.4]
  assign RetimeWrapper_73_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11551.4]
  assign RetimeWrapper_73_io_in = _T_1724 & io_rPort_18_en_0; // @[package.scala 94:16:@11550.4]
  assign RetimeWrapper_74_clock = clock; // @[:@11556.4]
  assign RetimeWrapper_74_reset = reset; // @[:@11557.4]
  assign RetimeWrapper_74_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11559.4]
  assign RetimeWrapper_74_io_in = _T_1948 & io_rPort_18_en_0; // @[package.scala 94:16:@11558.4]
  assign RetimeWrapper_75_clock = clock; // @[:@11564.4]
  assign RetimeWrapper_75_reset = reset; // @[:@11565.4]
  assign RetimeWrapper_75_io_flow = io_rPort_18_backpressure; // @[package.scala 95:18:@11567.4]
  assign RetimeWrapper_75_io_in = _T_2172 & io_rPort_18_en_0; // @[package.scala 94:16:@11566.4]
  assign RetimeWrapper_76_clock = clock; // @[:@11588.4]
  assign RetimeWrapper_76_reset = reset; // @[:@11589.4]
  assign RetimeWrapper_76_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11591.4]
  assign RetimeWrapper_76_io_in = _T_1421 & io_rPort_19_en_0; // @[package.scala 94:16:@11590.4]
  assign RetimeWrapper_77_clock = clock; // @[:@11596.4]
  assign RetimeWrapper_77_reset = reset; // @[:@11597.4]
  assign RetimeWrapper_77_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11599.4]
  assign RetimeWrapper_77_io_in = _T_1645 & io_rPort_19_en_0; // @[package.scala 94:16:@11598.4]
  assign RetimeWrapper_78_clock = clock; // @[:@11604.4]
  assign RetimeWrapper_78_reset = reset; // @[:@11605.4]
  assign RetimeWrapper_78_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11607.4]
  assign RetimeWrapper_78_io_in = _T_1869 & io_rPort_19_en_0; // @[package.scala 94:16:@11606.4]
  assign RetimeWrapper_79_clock = clock; // @[:@11612.4]
  assign RetimeWrapper_79_reset = reset; // @[:@11613.4]
  assign RetimeWrapper_79_io_flow = io_rPort_19_backpressure; // @[package.scala 95:18:@11615.4]
  assign RetimeWrapper_79_io_in = _T_2093 & io_rPort_19_en_0; // @[package.scala 94:16:@11614.4]
  assign RetimeWrapper_80_clock = clock; // @[:@11636.4]
  assign RetimeWrapper_80_reset = reset; // @[:@11637.4]
  assign RetimeWrapper_80_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11639.4]
  assign RetimeWrapper_80_io_in = _T_1426 & io_rPort_20_en_0; // @[package.scala 94:16:@11638.4]
  assign RetimeWrapper_81_clock = clock; // @[:@11644.4]
  assign RetimeWrapper_81_reset = reset; // @[:@11645.4]
  assign RetimeWrapper_81_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11647.4]
  assign RetimeWrapper_81_io_in = _T_1650 & io_rPort_20_en_0; // @[package.scala 94:16:@11646.4]
  assign RetimeWrapper_82_clock = clock; // @[:@11652.4]
  assign RetimeWrapper_82_reset = reset; // @[:@11653.4]
  assign RetimeWrapper_82_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11655.4]
  assign RetimeWrapper_82_io_in = _T_1874 & io_rPort_20_en_0; // @[package.scala 94:16:@11654.4]
  assign RetimeWrapper_83_clock = clock; // @[:@11660.4]
  assign RetimeWrapper_83_reset = reset; // @[:@11661.4]
  assign RetimeWrapper_83_io_flow = io_rPort_20_backpressure; // @[package.scala 95:18:@11663.4]
  assign RetimeWrapper_83_io_in = _T_2098 & io_rPort_20_en_0; // @[package.scala 94:16:@11662.4]
  assign RetimeWrapper_84_clock = clock; // @[:@11684.4]
  assign RetimeWrapper_84_reset = reset; // @[:@11685.4]
  assign RetimeWrapper_84_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11687.4]
  assign RetimeWrapper_84_io_in = _T_1505 & io_rPort_21_en_0; // @[package.scala 94:16:@11686.4]
  assign RetimeWrapper_85_clock = clock; // @[:@11692.4]
  assign RetimeWrapper_85_reset = reset; // @[:@11693.4]
  assign RetimeWrapper_85_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11695.4]
  assign RetimeWrapper_85_io_in = _T_1729 & io_rPort_21_en_0; // @[package.scala 94:16:@11694.4]
  assign RetimeWrapper_86_clock = clock; // @[:@11700.4]
  assign RetimeWrapper_86_reset = reset; // @[:@11701.4]
  assign RetimeWrapper_86_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11703.4]
  assign RetimeWrapper_86_io_in = _T_1953 & io_rPort_21_en_0; // @[package.scala 94:16:@11702.4]
  assign RetimeWrapper_87_clock = clock; // @[:@11708.4]
  assign RetimeWrapper_87_reset = reset; // @[:@11709.4]
  assign RetimeWrapper_87_io_flow = io_rPort_21_backpressure; // @[package.scala 95:18:@11711.4]
  assign RetimeWrapper_87_io_in = _T_2177 & io_rPort_21_en_0; // @[package.scala 94:16:@11710.4]
  assign RetimeWrapper_88_clock = clock; // @[:@11732.4]
  assign RetimeWrapper_88_reset = reset; // @[:@11733.4]
  assign RetimeWrapper_88_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11735.4]
  assign RetimeWrapper_88_io_in = _T_1431 & io_rPort_22_en_0; // @[package.scala 94:16:@11734.4]
  assign RetimeWrapper_89_clock = clock; // @[:@11740.4]
  assign RetimeWrapper_89_reset = reset; // @[:@11741.4]
  assign RetimeWrapper_89_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11743.4]
  assign RetimeWrapper_89_io_in = _T_1655 & io_rPort_22_en_0; // @[package.scala 94:16:@11742.4]
  assign RetimeWrapper_90_clock = clock; // @[:@11748.4]
  assign RetimeWrapper_90_reset = reset; // @[:@11749.4]
  assign RetimeWrapper_90_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11751.4]
  assign RetimeWrapper_90_io_in = _T_1879 & io_rPort_22_en_0; // @[package.scala 94:16:@11750.4]
  assign RetimeWrapper_91_clock = clock; // @[:@11756.4]
  assign RetimeWrapper_91_reset = reset; // @[:@11757.4]
  assign RetimeWrapper_91_io_flow = io_rPort_22_backpressure; // @[package.scala 95:18:@11759.4]
  assign RetimeWrapper_91_io_in = _T_2103 & io_rPort_22_en_0; // @[package.scala 94:16:@11758.4]
  assign RetimeWrapper_92_clock = clock; // @[:@11780.4]
  assign RetimeWrapper_92_reset = reset; // @[:@11781.4]
  assign RetimeWrapper_92_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11783.4]
  assign RetimeWrapper_92_io_in = _T_1335 & io_rPort_23_en_0; // @[package.scala 94:16:@11782.4]
  assign RetimeWrapper_93_clock = clock; // @[:@11788.4]
  assign RetimeWrapper_93_reset = reset; // @[:@11789.4]
  assign RetimeWrapper_93_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11791.4]
  assign RetimeWrapper_93_io_in = _T_1559 & io_rPort_23_en_0; // @[package.scala 94:16:@11790.4]
  assign RetimeWrapper_94_clock = clock; // @[:@11796.4]
  assign RetimeWrapper_94_reset = reset; // @[:@11797.4]
  assign RetimeWrapper_94_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11799.4]
  assign RetimeWrapper_94_io_in = _T_1783 & io_rPort_23_en_0; // @[package.scala 94:16:@11798.4]
  assign RetimeWrapper_95_clock = clock; // @[:@11804.4]
  assign RetimeWrapper_95_reset = reset; // @[:@11805.4]
  assign RetimeWrapper_95_io_flow = io_rPort_23_backpressure; // @[package.scala 95:18:@11807.4]
  assign RetimeWrapper_95_io_in = _T_2007 & io_rPort_23_en_0; // @[package.scala 94:16:@11806.4]
endmodule
module RetimeWrapper_148( // @[:@11827.2]
  input         clock, // @[:@11828.4]
  input         reset, // @[:@11829.4]
  input         io_flow, // @[:@11830.4]
  input  [63:0] io_in, // @[:@11830.4]
  output [63:0] io_out // @[:@11830.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11832.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11832.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11845.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11844.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@11843.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11842.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11841.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11839.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@11847.2]
  input  [31:0] io_a, // @[:@11850.4]
  output [32:0] io_b // @[:@11850.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@11857.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@11857.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@11862.4]
endmodule
module __2( // @[:@11864.2]
  input  [31:0] io_b, // @[:@11867.4]
  output [32:0] io_result // @[:@11867.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@11872.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@11872.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@11872.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@11885.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@11880.4]
endmodule
module RetimeWrapper_149( // @[:@11939.2]
  input         clock, // @[:@11940.4]
  input         reset, // @[:@11941.4]
  input         io_flow, // @[:@11942.4]
  input  [31:0] io_in, // @[:@11942.4]
  output [31:0] io_out // @[:@11942.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@11944.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@11944.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@11957.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@11956.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@11955.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@11954.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@11953.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@11951.4]
endmodule
module fix2fixBox( // @[:@11959.2]
  input         clock, // @[:@11960.4]
  input         reset, // @[:@11961.4]
  input  [32:0] io_a, // @[:@11962.4]
  input         io_flow, // @[:@11962.4]
  output [31:0] io_b // @[:@11962.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@11972.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@11972.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@11972.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@11972.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@11972.4]
  RetimeWrapper_149 RetimeWrapper ( // @[package.scala 93:22:@11972.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@11979.4]
  assign RetimeWrapper_clock = clock; // @[:@11973.4]
  assign RetimeWrapper_reset = reset; // @[:@11974.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@11976.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@11975.4]
endmodule
module x553_sum( // @[:@11981.2]
  input         clock, // @[:@11982.4]
  input         reset, // @[:@11983.4]
  input  [31:0] io_a, // @[:@11984.4]
  input  [31:0] io_b, // @[:@11984.4]
  input         io_flow, // @[:@11984.4]
  output [31:0] io_result // @[:@11984.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@11992.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@11992.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@11999.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@11999.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@12017.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@12017.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@12017.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@12017.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@12017.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@11997.4 Math.scala 713:14:@11998.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@12004.4 Math.scala 713:14:@12005.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@12006.4]
  __2 _ ( // @[Math.scala 709:24:@11992.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@11999.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@12017.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@11997.4 Math.scala 713:14:@11998.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@12004.4 Math.scala 713:14:@12005.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@12006.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@12025.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@11995.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@12002.4]
  assign fix2fixBox_clock = clock; // @[:@12018.4]
  assign fix2fixBox_reset = reset; // @[:@12019.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@12020.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@12023.4]
endmodule
module RetimeWrapper_150( // @[:@12039.2]
  input   clock, // @[:@12040.4]
  input   reset, // @[:@12041.4]
  input   io_flow, // @[:@12042.4]
  input   io_in, // @[:@12042.4]
  output  io_out // @[:@12042.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12044.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@12044.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12057.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12056.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@12055.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12054.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12053.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12051.4]
endmodule
module RetimeWrapper_152( // @[:@12103.2]
  input         clock, // @[:@12104.4]
  input         reset, // @[:@12105.4]
  input         io_flow, // @[:@12106.4]
  input  [31:0] io_in, // @[:@12106.4]
  output [31:0] io_out // @[:@12106.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12108.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@12108.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12121.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12120.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12119.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12118.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12117.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12115.4]
endmodule
module RetimeWrapper_153( // @[:@12135.2]
  input        clock, // @[:@12136.4]
  input        reset, // @[:@12137.4]
  input        io_flow, // @[:@12138.4]
  input  [7:0] io_in, // @[:@12138.4]
  output [7:0] io_out // @[:@12138.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12140.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@12140.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12153.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12152.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@12151.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12150.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12149.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12147.4]
endmodule
module RetimeWrapper_154( // @[:@12167.2]
  input         clock, // @[:@12168.4]
  input         reset, // @[:@12169.4]
  input         io_flow, // @[:@12170.4]
  input  [31:0] io_in, // @[:@12170.4]
  output [31:0] io_out // @[:@12170.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12172.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12172.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12172.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12172.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12172.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12172.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@12172.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12185.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12184.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12183.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12182.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12181.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12179.4]
endmodule
module RetimeWrapper_159( // @[:@12623.2]
  input         clock, // @[:@12624.4]
  input         reset, // @[:@12625.4]
  input         io_flow, // @[:@12626.4]
  input  [31:0] io_in, // @[:@12626.4]
  output [31:0] io_out // @[:@12626.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@12628.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@12628.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@12628.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@12628.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@12628.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@12628.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@12628.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@12641.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@12640.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@12639.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@12638.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@12637.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@12635.4]
endmodule
module RetimeWrapper_191( // @[:@14979.2]
  input         clock, // @[:@14980.4]
  input         reset, // @[:@14981.4]
  input         io_flow, // @[:@14982.4]
  input  [31:0] io_in, // @[:@14982.4]
  output [31:0] io_out // @[:@14982.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14984.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@14984.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14997.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14996.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14995.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14994.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14993.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14991.4]
endmodule
module RetimeWrapper_195( // @[:@15255.2]
  input   clock, // @[:@15256.4]
  input   reset, // @[:@15257.4]
  input   io_flow, // @[:@15258.4]
  input   io_in, // @[:@15258.4]
  output  io_out // @[:@15258.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15260.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15260.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15260.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15260.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15260.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15260.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@15260.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15273.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15272.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15271.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15270.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15269.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15267.4]
endmodule
module RetimeWrapper_212( // @[:@16095.2]
  input         clock, // @[:@16096.4]
  input         reset, // @[:@16097.4]
  input         io_flow, // @[:@16098.4]
  input  [31:0] io_in, // @[:@16098.4]
  output [31:0] io_out // @[:@16098.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16100.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@16100.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16113.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16112.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16111.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16110.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16109.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16107.4]
endmodule
module RetimeWrapper_229( // @[:@17527.2]
  input         clock, // @[:@17528.4]
  input         reset, // @[:@17529.4]
  input         io_flow, // @[:@17530.4]
  input  [31:0] io_in, // @[:@17530.4]
  output [31:0] io_out // @[:@17530.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17532.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@17532.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17545.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17544.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17543.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17542.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17541.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17539.4]
endmodule
module SimBlackBoxesfix2fixBox_82( // @[:@22215.2]
  input  [7:0] io_a, // @[:@22218.4]
  output [8:0] io_b // @[:@22218.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@22229.4]
endmodule
module __82( // @[:@22231.2]
  input  [7:0] io_b, // @[:@22234.4]
  output [8:0] io_result // @[:@22234.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@22239.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@22239.4]
  SimBlackBoxesfix2fixBox_82 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@22239.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@22252.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@22247.4]
endmodule
module fix2fixBox_40( // @[:@22325.2]
  input        clock, // @[:@22326.4]
  input        reset, // @[:@22327.4]
  input  [8:0] io_a, // @[:@22328.4]
  input        io_flow, // @[:@22328.4]
  output [7:0] io_b // @[:@22328.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22338.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22338.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22338.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@22338.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@22338.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@22338.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@22345.4]
  assign RetimeWrapper_clock = clock; // @[:@22339.4]
  assign RetimeWrapper_reset = reset; // @[:@22340.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@22342.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@22341.4]
endmodule
module x825_x17( // @[:@22347.2]
  input        clock, // @[:@22348.4]
  input        reset, // @[:@22349.4]
  input  [7:0] io_a, // @[:@22350.4]
  input  [7:0] io_b, // @[:@22350.4]
  input        io_flow, // @[:@22350.4]
  output [7:0] io_result // @[:@22350.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22358.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22358.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22365.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22365.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@22375.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@22375.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22375.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@22375.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22375.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22363.4 Math.scala 713:14:@22364.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22370.4 Math.scala 713:14:@22371.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22372.4]
  __82 _ ( // @[Math.scala 709:24:@22358.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@22365.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_40 fix2fixBox ( // @[Math.scala 141:30:@22375.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22363.4 Math.scala 713:14:@22364.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22370.4 Math.scala 713:14:@22371.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22372.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22383.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22361.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22368.4]
  assign fix2fixBox_clock = clock; // @[:@22376.4]
  assign fix2fixBox_reset = reset; // @[:@22377.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22378.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@22381.4]
endmodule
module fix2fixBox_44( // @[:@22973.2]
  input  [8:0] io_a, // @[:@22976.4]
  output [7:0] io_b // @[:@22976.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@22986.4]
endmodule
module x829_x17( // @[:@22988.2]
  input  [7:0] io_a, // @[:@22991.4]
  input  [7:0] io_b, // @[:@22991.4]
  output [7:0] io_result // @[:@22991.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22999.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22999.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@23006.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@23006.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@23016.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@23016.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@23004.4 Math.scala 713:14:@23005.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@23011.4 Math.scala 713:14:@23012.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@23013.4]
  __82 _ ( // @[Math.scala 709:24:@22999.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@23006.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_44 fix2fixBox ( // @[Math.scala 141:30:@23016.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@23004.4 Math.scala 713:14:@23005.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@23011.4 Math.scala 713:14:@23012.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@23013.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@23024.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@23002.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@23009.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@23019.4]
endmodule
module RetimeWrapper_294( // @[:@23495.2]
  input        clock, // @[:@23496.4]
  input        reset, // @[:@23497.4]
  input        io_flow, // @[:@23498.4]
  input  [7:0] io_in, // @[:@23498.4]
  output [7:0] io_out // @[:@23498.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23500.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23500.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23500.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23500.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23500.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23500.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@23500.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23513.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23512.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@23511.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23510.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23509.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23507.4]
endmodule
module x834_sub( // @[:@23608.2]
  input  [7:0] io_a, // @[:@23611.4]
  input  [7:0] io_b, // @[:@23611.4]
  output [7:0] io_result // @[:@23611.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@23619.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@23619.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@23626.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@23626.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 182:30:@23637.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 182:30:@23637.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@23624.4 Math.scala 713:14:@23625.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@23631.4 Math.scala 713:14:@23632.4]
  wire [9:0] _T_21; // @[Math.scala 177:37:@23633.4]
  wire [9:0] _T_22; // @[Math.scala 177:37:@23634.4]
  __82 _ ( // @[Math.scala 709:24:@23619.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __82 __1 ( // @[Math.scala 709:24:@23626.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_44 fix2fixBox ( // @[Math.scala 182:30:@23637.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@23624.4 Math.scala 713:14:@23625.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@23631.4 Math.scala 713:14:@23632.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@23633.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@23634.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@23645.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@23622.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@23629.4]
  assign fix2fixBox_io_a = _T_22[8:0]; // @[Math.scala 183:23:@23640.4]
endmodule
module RetimeWrapper_296( // @[:@23691.2]
  input        clock, // @[:@23692.4]
  input        reset, // @[:@23693.4]
  input        io_flow, // @[:@23694.4]
  input  [7:0] io_in, // @[:@23694.4]
  output [7:0] io_out // @[:@23694.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23696.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23696.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23696.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23696.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23696.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23696.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@23696.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23709.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23708.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@23707.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23706.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23705.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23703.4]
endmodule
module SimBlackBoxesfix2fixBox_100( // @[:@23711.2]
  input  [7:0] io_a, // @[:@23714.4]
  output [7:0] io_b // @[:@23714.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@23724.4]
endmodule
module __100( // @[:@23726.2]
  input  [7:0] io_b, // @[:@23729.4]
  output [7:0] io_result // @[:@23729.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@23734.4]
  wire [7:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@23734.4]
  SimBlackBoxesfix2fixBox_100 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@23734.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@23747.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@23742.4]
endmodule
module x838_div( // @[:@23749.2]
  input        clock, // @[:@23750.4]
  input        reset, // @[:@23751.4]
  input  [7:0] io_a, // @[:@23752.4]
  input        io_flow, // @[:@23752.4]
  output [7:0] io_result // @[:@23752.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23759.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23759.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23759.4]
  wire [7:0] __io_b; // @[Math.scala 709:24:@23769.4]
  wire [7:0] __io_result; // @[Math.scala 709:24:@23769.4]
  RetimeWrapper_296 RetimeWrapper ( // @[package.scala 93:22:@23759.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  __100 _ ( // @[Math.scala 709:24:@23769.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign io_result = __io_result; // @[Math.scala 291:34:@23777.4]
  assign RetimeWrapper_clock = clock; // @[:@23760.4]
  assign RetimeWrapper_reset = reset; // @[:@23761.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@23763.4]
  assign RetimeWrapper_io_in = io_a / 8'h5; // @[package.scala 94:16:@23762.4]
  assign __io_b = RetimeWrapper_io_out; // @[Math.scala 710:17:@23772.4]
endmodule
module RetimeWrapper_297( // @[:@23791.2]
  input        clock, // @[:@23792.4]
  input        reset, // @[:@23793.4]
  input        io_flow, // @[:@23794.4]
  input  [7:0] io_in, // @[:@23794.4]
  output [7:0] io_out // @[:@23794.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23796.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23796.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23796.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23796.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23796.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23796.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@23796.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23809.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23808.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@23807.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23806.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23805.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23803.4]
endmodule
module RetimeWrapper_298( // @[:@23954.2]
  input        clock, // @[:@23955.4]
  input        reset, // @[:@23956.4]
  input        io_flow, // @[:@23957.4]
  input  [7:0] io_in, // @[:@23957.4]
  output [7:0] io_out // @[:@23957.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23959.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23959.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23959.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23959.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23959.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23959.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@23959.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23972.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23971.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@23970.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23969.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23968.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23966.4]
endmodule
module RetimeWrapper_299( // @[:@23986.2]
  input   clock, // @[:@23987.4]
  input   reset, // @[:@23988.4]
  input   io_flow, // @[:@23989.4]
  input   io_in, // @[:@23989.4]
  output  io_out // @[:@23989.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@23991.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@23991.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@23991.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23991.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23991.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23991.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@23991.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24004.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24003.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@24002.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24001.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24000.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23998.4]
endmodule
module RetimeWrapper_384( // @[:@36555.2]
  input         clock, // @[:@36556.4]
  input         reset, // @[:@36557.4]
  input         io_flow, // @[:@36558.4]
  input  [63:0] io_in, // @[:@36558.4]
  output [63:0] io_out // @[:@36558.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36560.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36560.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36560.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36560.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36560.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36560.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@36560.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36573.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36572.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@36571.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36570.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36569.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36567.4]
endmodule
module x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@36671.2]
  input          clock, // @[:@36672.4]
  input          reset, // @[:@36673.4]
  output         io_in_x527_TVALID, // @[:@36674.4]
  input          io_in_x527_TREADY, // @[:@36674.4]
  output [255:0] io_in_x527_TDATA, // @[:@36674.4]
  output         io_in_x526_TREADY, // @[:@36674.4]
  input  [255:0] io_in_x526_TDATA, // @[:@36674.4]
  input  [7:0]   io_in_x526_TID, // @[:@36674.4]
  input  [7:0]   io_in_x526_TDEST, // @[:@36674.4]
  input          io_sigsIn_backpressure, // @[:@36674.4]
  input          io_sigsIn_datapathEn, // @[:@36674.4]
  input          io_sigsIn_break, // @[:@36674.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@36674.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@36674.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@36674.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@36674.4]
  input          io_rr // @[:@36674.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@36688.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@36688.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@36700.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@36700.4]
  wire  x539_lb_0_clock; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_reset; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_23_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_23_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_23_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_23_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_23_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_22_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_22_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_22_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_22_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_22_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_21_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_21_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_21_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_21_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_21_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_20_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_20_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_20_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_20_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_20_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_19_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_19_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_19_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_19_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_19_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_18_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_18_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_18_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_18_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_18_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_17_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_17_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_17_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_17_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_17_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_16_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_16_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_16_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_16_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_16_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_15_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_15_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_15_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_15_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_15_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_14_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_14_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_14_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_14_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_14_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_13_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_13_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_13_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_13_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_13_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_12_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_12_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_12_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_12_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_12_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_11_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_11_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_11_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_11_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_11_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_10_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_10_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_10_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_10_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_10_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_9_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_9_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_9_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_9_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_9_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_8_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_8_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_8_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_8_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_8_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_7_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_7_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_7_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_7_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_7_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_6_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_6_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_6_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_6_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_6_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_5_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_5_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_5_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_5_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_5_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_4_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_4_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_4_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_4_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_4_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_3_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_3_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_3_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_3_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_3_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_2_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_2_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_2_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_2_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_2_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_1_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_1_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_1_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_1_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_1_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_rPort_0_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_0_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_0_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_rPort_0_backpressure; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_rPort_0_output_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_7_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_7_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_7_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_7_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_6_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_6_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_6_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_6_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_5_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_5_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_5_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_5_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_4_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_4_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_4_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_4_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_3_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_3_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_3_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_3_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_2_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_2_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_2_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_2_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_1_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_1_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_1_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_1_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [2:0] x539_lb_0_io_wPort_0_banks_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_0_ofs_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire [7:0] x539_lb_0_io_wPort_0_data_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  x539_lb_0_io_wPort_0_en_0; // @[m_x539_lb_0.scala 57:17:@36710.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36936.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36936.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36936.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@36936.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@36936.4]
  wire  x553_sum_1_clock; // @[Math.scala 150:24:@37044.4]
  wire  x553_sum_1_reset; // @[Math.scala 150:24:@37044.4]
  wire [31:0] x553_sum_1_io_a; // @[Math.scala 150:24:@37044.4]
  wire [31:0] x553_sum_1_io_b; // @[Math.scala 150:24:@37044.4]
  wire  x553_sum_1_io_flow; // @[Math.scala 150:24:@37044.4]
  wire [31:0] x553_sum_1_io_result; // @[Math.scala 150:24:@37044.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37054.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37054.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37054.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37054.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37054.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@37063.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@37063.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@37063.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@37063.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@37063.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@37072.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@37072.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@37072.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@37072.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@37072.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@37081.4]
  wire [7:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@37081.4]
  wire [7:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@37081.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@37090.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@37090.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@37090.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@37090.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@37090.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@37103.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@37103.4]
  wire  x559_rdcol_1_clock; // @[Math.scala 150:24:@37126.4]
  wire  x559_rdcol_1_reset; // @[Math.scala 150:24:@37126.4]
  wire [31:0] x559_rdcol_1_io_a; // @[Math.scala 150:24:@37126.4]
  wire [31:0] x559_rdcol_1_io_b; // @[Math.scala 150:24:@37126.4]
  wire  x559_rdcol_1_io_flow; // @[Math.scala 150:24:@37126.4]
  wire [31:0] x559_rdcol_1_io_result; // @[Math.scala 150:24:@37126.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@37147.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@37147.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@37147.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@37147.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@37147.4]
  wire  x563_sum_1_clock; // @[Math.scala 150:24:@37156.4]
  wire  x563_sum_1_reset; // @[Math.scala 150:24:@37156.4]
  wire [31:0] x563_sum_1_io_a; // @[Math.scala 150:24:@37156.4]
  wire [31:0] x563_sum_1_io_b; // @[Math.scala 150:24:@37156.4]
  wire  x563_sum_1_io_flow; // @[Math.scala 150:24:@37156.4]
  wire [31:0] x563_sum_1_io_result; // @[Math.scala 150:24:@37156.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@37166.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@37166.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@37166.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@37166.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@37166.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@37175.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@37175.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@37175.4]
  wire [7:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@37175.4]
  wire [7:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@37175.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@37188.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@37188.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@37188.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@37188.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@37188.4]
  wire  x568_rdcol_1_clock; // @[Math.scala 150:24:@37211.4]
  wire  x568_rdcol_1_reset; // @[Math.scala 150:24:@37211.4]
  wire [31:0] x568_rdcol_1_io_a; // @[Math.scala 150:24:@37211.4]
  wire [31:0] x568_rdcol_1_io_b; // @[Math.scala 150:24:@37211.4]
  wire  x568_rdcol_1_io_flow; // @[Math.scala 150:24:@37211.4]
  wire [31:0] x568_rdcol_1_io_result; // @[Math.scala 150:24:@37211.4]
  wire  x572_sum_1_clock; // @[Math.scala 150:24:@37232.4]
  wire  x572_sum_1_reset; // @[Math.scala 150:24:@37232.4]
  wire [31:0] x572_sum_1_io_a; // @[Math.scala 150:24:@37232.4]
  wire [31:0] x572_sum_1_io_b; // @[Math.scala 150:24:@37232.4]
  wire  x572_sum_1_io_flow; // @[Math.scala 150:24:@37232.4]
  wire [31:0] x572_sum_1_io_result; // @[Math.scala 150:24:@37232.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@37242.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@37242.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@37242.4]
  wire [7:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@37242.4]
  wire [7:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@37242.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@37251.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@37251.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@37251.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@37251.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@37251.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@37264.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@37264.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@37264.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@37264.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@37264.4]
  wire  x577_rdcol_1_clock; // @[Math.scala 150:24:@37287.4]
  wire  x577_rdcol_1_reset; // @[Math.scala 150:24:@37287.4]
  wire [31:0] x577_rdcol_1_io_a; // @[Math.scala 150:24:@37287.4]
  wire [31:0] x577_rdcol_1_io_b; // @[Math.scala 150:24:@37287.4]
  wire  x577_rdcol_1_io_flow; // @[Math.scala 150:24:@37287.4]
  wire [31:0] x577_rdcol_1_io_result; // @[Math.scala 150:24:@37287.4]
  wire  x581_sum_1_clock; // @[Math.scala 150:24:@37308.4]
  wire  x581_sum_1_reset; // @[Math.scala 150:24:@37308.4]
  wire [31:0] x581_sum_1_io_a; // @[Math.scala 150:24:@37308.4]
  wire [31:0] x581_sum_1_io_b; // @[Math.scala 150:24:@37308.4]
  wire  x581_sum_1_io_flow; // @[Math.scala 150:24:@37308.4]
  wire [31:0] x581_sum_1_io_result; // @[Math.scala 150:24:@37308.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@37318.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@37318.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@37318.4]
  wire [7:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@37318.4]
  wire [7:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@37318.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@37327.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@37327.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@37327.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@37327.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@37327.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@37340.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@37340.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@37340.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@37340.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@37340.4]
  wire  x586_rdrow_1_clock; // @[Math.scala 150:24:@37363.4]
  wire  x586_rdrow_1_reset; // @[Math.scala 150:24:@37363.4]
  wire [31:0] x586_rdrow_1_io_a; // @[Math.scala 150:24:@37363.4]
  wire [31:0] x586_rdrow_1_io_b; // @[Math.scala 150:24:@37363.4]
  wire  x586_rdrow_1_io_flow; // @[Math.scala 150:24:@37363.4]
  wire [31:0] x586_rdrow_1_io_result; // @[Math.scala 150:24:@37363.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@37444.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@37444.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@37444.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@37444.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@37444.4]
  wire  x595_sum_1_clock; // @[Math.scala 150:24:@37453.4]
  wire  x595_sum_1_reset; // @[Math.scala 150:24:@37453.4]
  wire [31:0] x595_sum_1_io_a; // @[Math.scala 150:24:@37453.4]
  wire [31:0] x595_sum_1_io_b; // @[Math.scala 150:24:@37453.4]
  wire  x595_sum_1_io_flow; // @[Math.scala 150:24:@37453.4]
  wire [31:0] x595_sum_1_io_result; // @[Math.scala 150:24:@37453.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@37463.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@37463.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@37463.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@37463.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@37463.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@37472.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@37472.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@37472.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@37472.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@37472.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@37481.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@37481.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@37481.4]
  wire [7:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@37481.4]
  wire [7:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@37481.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@37494.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@37494.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@37494.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@37494.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@37494.4]
  wire  x601_sum_1_clock; // @[Math.scala 150:24:@37517.4]
  wire  x601_sum_1_reset; // @[Math.scala 150:24:@37517.4]
  wire [31:0] x601_sum_1_io_a; // @[Math.scala 150:24:@37517.4]
  wire [31:0] x601_sum_1_io_b; // @[Math.scala 150:24:@37517.4]
  wire  x601_sum_1_io_flow; // @[Math.scala 150:24:@37517.4]
  wire [31:0] x601_sum_1_io_result; // @[Math.scala 150:24:@37517.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@37527.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@37527.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@37527.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@37527.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@37527.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@37536.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@37536.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@37536.4]
  wire [7:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@37536.4]
  wire [7:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@37536.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@37549.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@37549.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@37549.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@37549.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@37549.4]
  wire  x606_sum_1_clock; // @[Math.scala 150:24:@37572.4]
  wire  x606_sum_1_reset; // @[Math.scala 150:24:@37572.4]
  wire [31:0] x606_sum_1_io_a; // @[Math.scala 150:24:@37572.4]
  wire [31:0] x606_sum_1_io_b; // @[Math.scala 150:24:@37572.4]
  wire  x606_sum_1_io_flow; // @[Math.scala 150:24:@37572.4]
  wire [31:0] x606_sum_1_io_result; // @[Math.scala 150:24:@37572.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@37582.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@37582.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@37582.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@37582.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@37582.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@37591.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@37591.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@37591.4]
  wire [7:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@37591.4]
  wire [7:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@37591.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@37604.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@37604.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@37604.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@37604.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@37604.4]
  wire  x611_sum_1_clock; // @[Math.scala 150:24:@37627.4]
  wire  x611_sum_1_reset; // @[Math.scala 150:24:@37627.4]
  wire [31:0] x611_sum_1_io_a; // @[Math.scala 150:24:@37627.4]
  wire [31:0] x611_sum_1_io_b; // @[Math.scala 150:24:@37627.4]
  wire  x611_sum_1_io_flow; // @[Math.scala 150:24:@37627.4]
  wire [31:0] x611_sum_1_io_result; // @[Math.scala 150:24:@37627.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@37637.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@37637.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@37637.4]
  wire [7:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@37637.4]
  wire [7:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@37637.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@37646.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@37646.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@37646.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@37646.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@37646.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@37659.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@37680.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@37680.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@37680.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@37680.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@37680.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@37707.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@37707.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@37749.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@37749.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@37749.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@37749.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@37749.4]
  wire  x623_sum_1_clock; // @[Math.scala 150:24:@37758.4]
  wire  x623_sum_1_reset; // @[Math.scala 150:24:@37758.4]
  wire [31:0] x623_sum_1_io_a; // @[Math.scala 150:24:@37758.4]
  wire [31:0] x623_sum_1_io_b; // @[Math.scala 150:24:@37758.4]
  wire  x623_sum_1_io_flow; // @[Math.scala 150:24:@37758.4]
  wire [31:0] x623_sum_1_io_result; // @[Math.scala 150:24:@37758.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@37768.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@37768.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@37768.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@37768.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@37768.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@37777.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@37777.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@37777.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@37777.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@37777.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@37786.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@37786.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@37786.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@37786.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@37786.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@37795.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@37795.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@37795.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@37795.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@37795.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@37809.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@37809.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@37809.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@37809.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@37809.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@37830.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@37830.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@37830.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@37830.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@37830.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@37852.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@37852.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@37852.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@37852.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@37852.4]
  wire  x632_sum_1_clock; // @[Math.scala 150:24:@37861.4]
  wire  x632_sum_1_reset; // @[Math.scala 150:24:@37861.4]
  wire [31:0] x632_sum_1_io_a; // @[Math.scala 150:24:@37861.4]
  wire [31:0] x632_sum_1_io_b; // @[Math.scala 150:24:@37861.4]
  wire  x632_sum_1_io_flow; // @[Math.scala 150:24:@37861.4]
  wire [31:0] x632_sum_1_io_result; // @[Math.scala 150:24:@37861.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@37871.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@37871.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@37871.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@37871.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@37871.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@37885.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@37885.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@37885.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@37885.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@37885.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@37906.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@37906.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@37906.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@37906.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@37906.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@37930.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@37930.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@37930.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@37930.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@37930.4]
  wire  x640_sum_1_clock; // @[Math.scala 150:24:@37939.4]
  wire  x640_sum_1_reset; // @[Math.scala 150:24:@37939.4]
  wire [31:0] x640_sum_1_io_a; // @[Math.scala 150:24:@37939.4]
  wire [31:0] x640_sum_1_io_b; // @[Math.scala 150:24:@37939.4]
  wire  x640_sum_1_io_flow; // @[Math.scala 150:24:@37939.4]
  wire [31:0] x640_sum_1_io_result; // @[Math.scala 150:24:@37939.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@37949.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@37949.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@37949.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@37949.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@37949.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@37963.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@37963.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@37963.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@37963.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@37963.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@37984.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@37984.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@37984.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@37984.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@37984.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@38000.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@38000.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@38000.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@38000.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@38000.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@38015.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@38015.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@38015.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@38015.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@38015.4]
  wire  x648_sum_1_clock; // @[Math.scala 150:24:@38024.4]
  wire  x648_sum_1_reset; // @[Math.scala 150:24:@38024.4]
  wire [31:0] x648_sum_1_io_a; // @[Math.scala 150:24:@38024.4]
  wire [31:0] x648_sum_1_io_b; // @[Math.scala 150:24:@38024.4]
  wire  x648_sum_1_io_flow; // @[Math.scala 150:24:@38024.4]
  wire [31:0] x648_sum_1_io_result; // @[Math.scala 150:24:@38024.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@38034.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@38034.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@38034.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@38034.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@38034.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@38048.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@38048.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@38048.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@38048.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@38048.4]
  wire  x653_rdcol_1_clock; // @[Math.scala 150:24:@38071.4]
  wire  x653_rdcol_1_reset; // @[Math.scala 150:24:@38071.4]
  wire [31:0] x653_rdcol_1_io_a; // @[Math.scala 150:24:@38071.4]
  wire [31:0] x653_rdcol_1_io_b; // @[Math.scala 150:24:@38071.4]
  wire  x653_rdcol_1_io_flow; // @[Math.scala 150:24:@38071.4]
  wire [31:0] x653_rdcol_1_io_result; // @[Math.scala 150:24:@38071.4]
  wire  x659_sum_1_clock; // @[Math.scala 150:24:@38103.4]
  wire  x659_sum_1_reset; // @[Math.scala 150:24:@38103.4]
  wire [31:0] x659_sum_1_io_a; // @[Math.scala 150:24:@38103.4]
  wire [31:0] x659_sum_1_io_b; // @[Math.scala 150:24:@38103.4]
  wire  x659_sum_1_io_flow; // @[Math.scala 150:24:@38103.4]
  wire [31:0] x659_sum_1_io_result; // @[Math.scala 150:24:@38103.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@38113.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@38113.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@38113.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@38113.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@38113.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@38127.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@38127.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@38127.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@38127.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@38127.4]
  wire  x665_rdcol_1_clock; // @[Math.scala 150:24:@38150.4]
  wire  x665_rdcol_1_reset; // @[Math.scala 150:24:@38150.4]
  wire [31:0] x665_rdcol_1_io_a; // @[Math.scala 150:24:@38150.4]
  wire [31:0] x665_rdcol_1_io_b; // @[Math.scala 150:24:@38150.4]
  wire  x665_rdcol_1_io_flow; // @[Math.scala 150:24:@38150.4]
  wire [31:0] x665_rdcol_1_io_result; // @[Math.scala 150:24:@38150.4]
  wire  x671_sum_1_clock; // @[Math.scala 150:24:@38182.4]
  wire  x671_sum_1_reset; // @[Math.scala 150:24:@38182.4]
  wire [31:0] x671_sum_1_io_a; // @[Math.scala 150:24:@38182.4]
  wire [31:0] x671_sum_1_io_b; // @[Math.scala 150:24:@38182.4]
  wire  x671_sum_1_io_flow; // @[Math.scala 150:24:@38182.4]
  wire [31:0] x671_sum_1_io_result; // @[Math.scala 150:24:@38182.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@38192.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@38192.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@38192.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@38192.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@38192.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@38206.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@38227.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@38227.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@38227.4]
  wire [31:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@38227.4]
  wire [31:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@38227.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@38254.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@38254.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@38254.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@38254.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@38254.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@38289.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@38289.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@38289.4]
  wire [31:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@38289.4]
  wire [31:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@38289.4]
  wire  x683_sum_1_clock; // @[Math.scala 150:24:@38298.4]
  wire  x683_sum_1_reset; // @[Math.scala 150:24:@38298.4]
  wire [31:0] x683_sum_1_io_a; // @[Math.scala 150:24:@38298.4]
  wire [31:0] x683_sum_1_io_b; // @[Math.scala 150:24:@38298.4]
  wire  x683_sum_1_io_flow; // @[Math.scala 150:24:@38298.4]
  wire [31:0] x683_sum_1_io_result; // @[Math.scala 150:24:@38298.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@38308.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@38308.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@38308.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@38308.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@38308.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@38317.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@38317.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@38317.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@38317.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@38317.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@38331.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@38331.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@38331.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@38331.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@38331.4]
  wire  x691_sum_1_clock; // @[Math.scala 150:24:@38360.4]
  wire  x691_sum_1_reset; // @[Math.scala 150:24:@38360.4]
  wire [31:0] x691_sum_1_io_a; // @[Math.scala 150:24:@38360.4]
  wire [31:0] x691_sum_1_io_b; // @[Math.scala 150:24:@38360.4]
  wire  x691_sum_1_io_flow; // @[Math.scala 150:24:@38360.4]
  wire [31:0] x691_sum_1_io_result; // @[Math.scala 150:24:@38360.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@38370.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@38370.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@38370.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@38370.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@38370.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@38384.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@38384.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@38384.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@38384.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@38384.4]
  wire  x698_sum_1_clock; // @[Math.scala 150:24:@38411.4]
  wire  x698_sum_1_reset; // @[Math.scala 150:24:@38411.4]
  wire [31:0] x698_sum_1_io_a; // @[Math.scala 150:24:@38411.4]
  wire [31:0] x698_sum_1_io_b; // @[Math.scala 150:24:@38411.4]
  wire  x698_sum_1_io_flow; // @[Math.scala 150:24:@38411.4]
  wire [31:0] x698_sum_1_io_result; // @[Math.scala 150:24:@38411.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@38421.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@38421.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@38421.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@38421.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@38421.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@38435.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@38435.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@38435.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@38435.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@38435.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@38462.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@38462.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@38462.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@38462.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@38462.4]
  wire  x705_sum_1_clock; // @[Math.scala 150:24:@38471.4]
  wire  x705_sum_1_reset; // @[Math.scala 150:24:@38471.4]
  wire [31:0] x705_sum_1_io_a; // @[Math.scala 150:24:@38471.4]
  wire [31:0] x705_sum_1_io_b; // @[Math.scala 150:24:@38471.4]
  wire  x705_sum_1_io_flow; // @[Math.scala 150:24:@38471.4]
  wire [31:0] x705_sum_1_io_result; // @[Math.scala 150:24:@38471.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@38481.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@38481.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@38481.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@38481.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@38481.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@38490.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@38490.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@38490.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@38490.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@38490.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@38504.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@38504.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@38504.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@38504.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@38504.4]
  wire  x712_sum_1_clock; // @[Math.scala 150:24:@38531.4]
  wire  x712_sum_1_reset; // @[Math.scala 150:24:@38531.4]
  wire [31:0] x712_sum_1_io_a; // @[Math.scala 150:24:@38531.4]
  wire [31:0] x712_sum_1_io_b; // @[Math.scala 150:24:@38531.4]
  wire  x712_sum_1_io_flow; // @[Math.scala 150:24:@38531.4]
  wire [31:0] x712_sum_1_io_result; // @[Math.scala 150:24:@38531.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@38541.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@38541.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@38541.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@38541.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@38541.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@38555.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@38555.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@38555.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@38555.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@38555.4]
  wire  x719_sum_1_clock; // @[Math.scala 150:24:@38582.4]
  wire  x719_sum_1_reset; // @[Math.scala 150:24:@38582.4]
  wire [31:0] x719_sum_1_io_a; // @[Math.scala 150:24:@38582.4]
  wire [31:0] x719_sum_1_io_b; // @[Math.scala 150:24:@38582.4]
  wire  x719_sum_1_io_flow; // @[Math.scala 150:24:@38582.4]
  wire [31:0] x719_sum_1_io_result; // @[Math.scala 150:24:@38582.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@38592.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@38592.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@38592.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@38592.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@38592.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@38606.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@38606.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@38606.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@38606.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@38606.4]
  wire  x724_rdrow_1_clock; // @[Math.scala 150:24:@38629.4]
  wire  x724_rdrow_1_reset; // @[Math.scala 150:24:@38629.4]
  wire [31:0] x724_rdrow_1_io_a; // @[Math.scala 150:24:@38629.4]
  wire [31:0] x724_rdrow_1_io_b; // @[Math.scala 150:24:@38629.4]
  wire  x724_rdrow_1_io_flow; // @[Math.scala 150:24:@38629.4]
  wire [31:0] x724_rdrow_1_io_result; // @[Math.scala 150:24:@38629.4]
  wire  x731_sum_1_clock; // @[Math.scala 150:24:@38683.4]
  wire  x731_sum_1_reset; // @[Math.scala 150:24:@38683.4]
  wire [31:0] x731_sum_1_io_a; // @[Math.scala 150:24:@38683.4]
  wire [31:0] x731_sum_1_io_b; // @[Math.scala 150:24:@38683.4]
  wire  x731_sum_1_io_flow; // @[Math.scala 150:24:@38683.4]
  wire [31:0] x731_sum_1_io_result; // @[Math.scala 150:24:@38683.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@38693.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@38693.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@38693.4]
  wire [31:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@38693.4]
  wire [31:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@38693.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@38702.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@38702.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@38702.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@38702.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@38702.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@38716.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@38716.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@38716.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@38716.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@38716.4]
  wire  x739_sum_1_clock; // @[Math.scala 150:24:@38745.4]
  wire  x739_sum_1_reset; // @[Math.scala 150:24:@38745.4]
  wire [31:0] x739_sum_1_io_a; // @[Math.scala 150:24:@38745.4]
  wire [31:0] x739_sum_1_io_b; // @[Math.scala 150:24:@38745.4]
  wire  x739_sum_1_io_flow; // @[Math.scala 150:24:@38745.4]
  wire [31:0] x739_sum_1_io_result; // @[Math.scala 150:24:@38745.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@38755.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@38755.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@38755.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@38755.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@38755.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@38769.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@38769.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@38769.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@38769.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@38769.4]
  wire  x746_sum_1_clock; // @[Math.scala 150:24:@38796.4]
  wire  x746_sum_1_reset; // @[Math.scala 150:24:@38796.4]
  wire [31:0] x746_sum_1_io_a; // @[Math.scala 150:24:@38796.4]
  wire [31:0] x746_sum_1_io_b; // @[Math.scala 150:24:@38796.4]
  wire  x746_sum_1_io_flow; // @[Math.scala 150:24:@38796.4]
  wire [31:0] x746_sum_1_io_result; // @[Math.scala 150:24:@38796.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@38806.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@38806.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@38806.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@38806.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@38806.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@38820.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@38820.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@38820.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@38820.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@38820.4]
  wire  x753_sum_1_clock; // @[Math.scala 150:24:@38847.4]
  wire  x753_sum_1_reset; // @[Math.scala 150:24:@38847.4]
  wire [31:0] x753_sum_1_io_a; // @[Math.scala 150:24:@38847.4]
  wire [31:0] x753_sum_1_io_b; // @[Math.scala 150:24:@38847.4]
  wire  x753_sum_1_io_flow; // @[Math.scala 150:24:@38847.4]
  wire [31:0] x753_sum_1_io_result; // @[Math.scala 150:24:@38847.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@38857.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@38857.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@38857.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@38857.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@38857.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@38871.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@38871.4]
  wire  x760_sum_1_clock; // @[Math.scala 150:24:@38898.4]
  wire  x760_sum_1_reset; // @[Math.scala 150:24:@38898.4]
  wire [31:0] x760_sum_1_io_a; // @[Math.scala 150:24:@38898.4]
  wire [31:0] x760_sum_1_io_b; // @[Math.scala 150:24:@38898.4]
  wire  x760_sum_1_io_flow; // @[Math.scala 150:24:@38898.4]
  wire [31:0] x760_sum_1_io_result; // @[Math.scala 150:24:@38898.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@38908.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@38922.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@38922.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@38922.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@38922.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@38922.4]
  wire  x767_sum_1_clock; // @[Math.scala 150:24:@38949.4]
  wire  x767_sum_1_reset; // @[Math.scala 150:24:@38949.4]
  wire [31:0] x767_sum_1_io_a; // @[Math.scala 150:24:@38949.4]
  wire [31:0] x767_sum_1_io_b; // @[Math.scala 150:24:@38949.4]
  wire  x767_sum_1_io_flow; // @[Math.scala 150:24:@38949.4]
  wire [31:0] x767_sum_1_io_result; // @[Math.scala 150:24:@38949.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@38959.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@38959.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@38959.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@38959.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@38959.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@38973.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@38973.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@38973.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@38973.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@38973.4]
  wire  x772_rdrow_1_clock; // @[Math.scala 150:24:@38996.4]
  wire  x772_rdrow_1_reset; // @[Math.scala 150:24:@38996.4]
  wire [31:0] x772_rdrow_1_io_a; // @[Math.scala 150:24:@38996.4]
  wire [31:0] x772_rdrow_1_io_b; // @[Math.scala 150:24:@38996.4]
  wire  x772_rdrow_1_io_flow; // @[Math.scala 150:24:@38996.4]
  wire [31:0] x772_rdrow_1_io_result; // @[Math.scala 150:24:@38996.4]
  wire  x779_sum_1_clock; // @[Math.scala 150:24:@39050.4]
  wire  x779_sum_1_reset; // @[Math.scala 150:24:@39050.4]
  wire [31:0] x779_sum_1_io_a; // @[Math.scala 150:24:@39050.4]
  wire [31:0] x779_sum_1_io_b; // @[Math.scala 150:24:@39050.4]
  wire  x779_sum_1_io_flow; // @[Math.scala 150:24:@39050.4]
  wire [31:0] x779_sum_1_io_result; // @[Math.scala 150:24:@39050.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@39060.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@39060.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@39060.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@39060.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@39060.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@39069.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@39069.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@39069.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@39069.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@39069.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@39083.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@39083.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@39083.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@39083.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@39083.4]
  wire  x787_sum_1_clock; // @[Math.scala 150:24:@39110.4]
  wire  x787_sum_1_reset; // @[Math.scala 150:24:@39110.4]
  wire [31:0] x787_sum_1_io_a; // @[Math.scala 150:24:@39110.4]
  wire [31:0] x787_sum_1_io_b; // @[Math.scala 150:24:@39110.4]
  wire  x787_sum_1_io_flow; // @[Math.scala 150:24:@39110.4]
  wire [31:0] x787_sum_1_io_result; // @[Math.scala 150:24:@39110.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@39120.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@39120.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@39120.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@39120.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@39120.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@39134.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@39134.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@39134.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@39134.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@39134.4]
  wire  x794_sum_1_clock; // @[Math.scala 150:24:@39163.4]
  wire  x794_sum_1_reset; // @[Math.scala 150:24:@39163.4]
  wire [31:0] x794_sum_1_io_a; // @[Math.scala 150:24:@39163.4]
  wire [31:0] x794_sum_1_io_b; // @[Math.scala 150:24:@39163.4]
  wire  x794_sum_1_io_flow; // @[Math.scala 150:24:@39163.4]
  wire [31:0] x794_sum_1_io_result; // @[Math.scala 150:24:@39163.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@39173.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@39173.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@39173.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@39173.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@39173.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@39187.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@39187.4]
  wire  x801_sum_1_clock; // @[Math.scala 150:24:@39214.4]
  wire  x801_sum_1_reset; // @[Math.scala 150:24:@39214.4]
  wire [31:0] x801_sum_1_io_a; // @[Math.scala 150:24:@39214.4]
  wire [31:0] x801_sum_1_io_b; // @[Math.scala 150:24:@39214.4]
  wire  x801_sum_1_io_flow; // @[Math.scala 150:24:@39214.4]
  wire [31:0] x801_sum_1_io_result; // @[Math.scala 150:24:@39214.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@39224.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@39224.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@39224.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@39224.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@39224.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@39238.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@39238.4]
  wire  x808_sum_1_clock; // @[Math.scala 150:24:@39265.4]
  wire  x808_sum_1_reset; // @[Math.scala 150:24:@39265.4]
  wire [31:0] x808_sum_1_io_a; // @[Math.scala 150:24:@39265.4]
  wire [31:0] x808_sum_1_io_b; // @[Math.scala 150:24:@39265.4]
  wire  x808_sum_1_io_flow; // @[Math.scala 150:24:@39265.4]
  wire [31:0] x808_sum_1_io_result; // @[Math.scala 150:24:@39265.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@39275.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@39275.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@39275.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@39275.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@39275.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@39289.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@39289.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@39289.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@39289.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@39289.4]
  wire  x815_sum_1_clock; // @[Math.scala 150:24:@39316.4]
  wire  x815_sum_1_reset; // @[Math.scala 150:24:@39316.4]
  wire [31:0] x815_sum_1_io_a; // @[Math.scala 150:24:@39316.4]
  wire [31:0] x815_sum_1_io_b; // @[Math.scala 150:24:@39316.4]
  wire  x815_sum_1_io_flow; // @[Math.scala 150:24:@39316.4]
  wire [31:0] x815_sum_1_io_result; // @[Math.scala 150:24:@39316.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@39326.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@39326.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@39326.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@39326.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@39326.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@39340.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@39340.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@39340.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@39340.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@39340.4]
  wire  x825_x17_1_clock; // @[Math.scala 150:24:@39386.4]
  wire  x825_x17_1_reset; // @[Math.scala 150:24:@39386.4]
  wire [7:0] x825_x17_1_io_a; // @[Math.scala 150:24:@39386.4]
  wire [7:0] x825_x17_1_io_b; // @[Math.scala 150:24:@39386.4]
  wire  x825_x17_1_io_flow; // @[Math.scala 150:24:@39386.4]
  wire [7:0] x825_x17_1_io_result; // @[Math.scala 150:24:@39386.4]
  wire  x826_x18_1_clock; // @[Math.scala 150:24:@39396.4]
  wire  x826_x18_1_reset; // @[Math.scala 150:24:@39396.4]
  wire [7:0] x826_x18_1_io_a; // @[Math.scala 150:24:@39396.4]
  wire [7:0] x826_x18_1_io_b; // @[Math.scala 150:24:@39396.4]
  wire  x826_x18_1_io_flow; // @[Math.scala 150:24:@39396.4]
  wire [7:0] x826_x18_1_io_result; // @[Math.scala 150:24:@39396.4]
  wire  x827_x17_1_clock; // @[Math.scala 150:24:@39406.4]
  wire  x827_x17_1_reset; // @[Math.scala 150:24:@39406.4]
  wire [7:0] x827_x17_1_io_a; // @[Math.scala 150:24:@39406.4]
  wire [7:0] x827_x17_1_io_b; // @[Math.scala 150:24:@39406.4]
  wire  x827_x17_1_io_flow; // @[Math.scala 150:24:@39406.4]
  wire [7:0] x827_x17_1_io_result; // @[Math.scala 150:24:@39406.4]
  wire  x828_x18_1_clock; // @[Math.scala 150:24:@39416.4]
  wire  x828_x18_1_reset; // @[Math.scala 150:24:@39416.4]
  wire [7:0] x828_x18_1_io_a; // @[Math.scala 150:24:@39416.4]
  wire [7:0] x828_x18_1_io_b; // @[Math.scala 150:24:@39416.4]
  wire  x828_x18_1_io_flow; // @[Math.scala 150:24:@39416.4]
  wire [7:0] x828_x18_1_io_result; // @[Math.scala 150:24:@39416.4]
  wire [7:0] x829_x17_1_io_a; // @[Math.scala 150:24:@39426.4]
  wire [7:0] x829_x17_1_io_b; // @[Math.scala 150:24:@39426.4]
  wire [7:0] x829_x17_1_io_result; // @[Math.scala 150:24:@39426.4]
  wire [7:0] x830_x18_1_io_a; // @[Math.scala 150:24:@39436.4]
  wire [7:0] x830_x18_1_io_b; // @[Math.scala 150:24:@39436.4]
  wire [7:0] x830_x18_1_io_result; // @[Math.scala 150:24:@39436.4]
  wire [7:0] x831_x17_1_io_a; // @[Math.scala 150:24:@39446.4]
  wire [7:0] x831_x17_1_io_b; // @[Math.scala 150:24:@39446.4]
  wire [7:0] x831_x17_1_io_result; // @[Math.scala 150:24:@39446.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@39456.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@39456.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@39456.4]
  wire [7:0] RetimeWrapper_100_io_in; // @[package.scala 93:22:@39456.4]
  wire [7:0] RetimeWrapper_100_io_out; // @[package.scala 93:22:@39456.4]
  wire [7:0] x832_sum_1_io_a; // @[Math.scala 150:24:@39465.4]
  wire [7:0] x832_sum_1_io_b; // @[Math.scala 150:24:@39465.4]
  wire [7:0] x832_sum_1_io_result; // @[Math.scala 150:24:@39465.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@39479.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@39479.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@39479.4]
  wire [7:0] RetimeWrapper_101_io_in; // @[package.scala 93:22:@39479.4]
  wire [7:0] RetimeWrapper_101_io_out; // @[package.scala 93:22:@39479.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@39489.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@39489.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@39489.4]
  wire [7:0] RetimeWrapper_102_io_in; // @[package.scala 93:22:@39489.4]
  wire [7:0] RetimeWrapper_102_io_out; // @[package.scala 93:22:@39489.4]
  wire [7:0] x834_sub_1_io_a; // @[Math.scala 191:24:@39498.4]
  wire [7:0] x834_sub_1_io_b; // @[Math.scala 191:24:@39498.4]
  wire [7:0] x834_sub_1_io_result; // @[Math.scala 191:24:@39498.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@39523.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@39523.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@39523.4]
  wire [7:0] RetimeWrapper_103_io_in; // @[package.scala 93:22:@39523.4]
  wire [7:0] RetimeWrapper_103_io_out; // @[package.scala 93:22:@39523.4]
  wire  x838_div_1_clock; // @[Math.scala 327:24:@39534.4]
  wire  x838_div_1_reset; // @[Math.scala 327:24:@39534.4]
  wire [7:0] x838_div_1_io_a; // @[Math.scala 327:24:@39534.4]
  wire  x838_div_1_io_flow; // @[Math.scala 327:24:@39534.4]
  wire [7:0] x838_div_1_io_result; // @[Math.scala 327:24:@39534.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@39544.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@39544.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@39544.4]
  wire [7:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@39544.4]
  wire [7:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@39544.4]
  wire [7:0] x839_sum_1_io_a; // @[Math.scala 150:24:@39553.4]
  wire [7:0] x839_sum_1_io_b; // @[Math.scala 150:24:@39553.4]
  wire [7:0] x839_sum_1_io_result; // @[Math.scala 150:24:@39553.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@39563.4]
  wire [7:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@39563.4]
  wire [7:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@39563.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@39572.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@39572.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@39572.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@39572.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@39572.4]
  wire  x846_x17_1_clock; // @[Math.scala 150:24:@39611.4]
  wire  x846_x17_1_reset; // @[Math.scala 150:24:@39611.4]
  wire [7:0] x846_x17_1_io_a; // @[Math.scala 150:24:@39611.4]
  wire [7:0] x846_x17_1_io_b; // @[Math.scala 150:24:@39611.4]
  wire  x846_x17_1_io_flow; // @[Math.scala 150:24:@39611.4]
  wire [7:0] x846_x17_1_io_result; // @[Math.scala 150:24:@39611.4]
  wire  x847_x18_1_clock; // @[Math.scala 150:24:@39621.4]
  wire  x847_x18_1_reset; // @[Math.scala 150:24:@39621.4]
  wire [7:0] x847_x18_1_io_a; // @[Math.scala 150:24:@39621.4]
  wire [7:0] x847_x18_1_io_b; // @[Math.scala 150:24:@39621.4]
  wire  x847_x18_1_io_flow; // @[Math.scala 150:24:@39621.4]
  wire [7:0] x847_x18_1_io_result; // @[Math.scala 150:24:@39621.4]
  wire  x848_x17_1_clock; // @[Math.scala 150:24:@39631.4]
  wire  x848_x17_1_reset; // @[Math.scala 150:24:@39631.4]
  wire [7:0] x848_x17_1_io_a; // @[Math.scala 150:24:@39631.4]
  wire [7:0] x848_x17_1_io_b; // @[Math.scala 150:24:@39631.4]
  wire  x848_x17_1_io_flow; // @[Math.scala 150:24:@39631.4]
  wire [7:0] x848_x17_1_io_result; // @[Math.scala 150:24:@39631.4]
  wire  x849_x18_1_clock; // @[Math.scala 150:24:@39641.4]
  wire  x849_x18_1_reset; // @[Math.scala 150:24:@39641.4]
  wire [7:0] x849_x18_1_io_a; // @[Math.scala 150:24:@39641.4]
  wire [7:0] x849_x18_1_io_b; // @[Math.scala 150:24:@39641.4]
  wire  x849_x18_1_io_flow; // @[Math.scala 150:24:@39641.4]
  wire [7:0] x849_x18_1_io_result; // @[Math.scala 150:24:@39641.4]
  wire [7:0] x850_x17_1_io_a; // @[Math.scala 150:24:@39651.4]
  wire [7:0] x850_x17_1_io_b; // @[Math.scala 150:24:@39651.4]
  wire [7:0] x850_x17_1_io_result; // @[Math.scala 150:24:@39651.4]
  wire [7:0] x851_x18_1_io_a; // @[Math.scala 150:24:@39661.4]
  wire [7:0] x851_x18_1_io_b; // @[Math.scala 150:24:@39661.4]
  wire [7:0] x851_x18_1_io_result; // @[Math.scala 150:24:@39661.4]
  wire [7:0] x852_x17_1_io_a; // @[Math.scala 150:24:@39671.4]
  wire [7:0] x852_x17_1_io_b; // @[Math.scala 150:24:@39671.4]
  wire [7:0] x852_x17_1_io_result; // @[Math.scala 150:24:@39671.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@39681.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@39681.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@39681.4]
  wire [7:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@39681.4]
  wire [7:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@39681.4]
  wire [7:0] x853_sum_1_io_a; // @[Math.scala 150:24:@39690.4]
  wire [7:0] x853_sum_1_io_b; // @[Math.scala 150:24:@39690.4]
  wire [7:0] x853_sum_1_io_result; // @[Math.scala 150:24:@39690.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@39704.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@39704.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@39704.4]
  wire [7:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@39704.4]
  wire [7:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@39704.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@39714.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@39714.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@39714.4]
  wire [7:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@39714.4]
  wire [7:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@39714.4]
  wire [7:0] x855_sub_1_io_a; // @[Math.scala 191:24:@39723.4]
  wire [7:0] x855_sub_1_io_b; // @[Math.scala 191:24:@39723.4]
  wire [7:0] x855_sub_1_io_result; // @[Math.scala 191:24:@39723.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@39748.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@39748.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@39748.4]
  wire [7:0] RetimeWrapper_110_io_in; // @[package.scala 93:22:@39748.4]
  wire [7:0] RetimeWrapper_110_io_out; // @[package.scala 93:22:@39748.4]
  wire  x859_div_1_clock; // @[Math.scala 327:24:@39759.4]
  wire  x859_div_1_reset; // @[Math.scala 327:24:@39759.4]
  wire [7:0] x859_div_1_io_a; // @[Math.scala 327:24:@39759.4]
  wire  x859_div_1_io_flow; // @[Math.scala 327:24:@39759.4]
  wire [7:0] x859_div_1_io_result; // @[Math.scala 327:24:@39759.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@39769.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@39769.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@39769.4]
  wire [7:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@39769.4]
  wire [7:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@39769.4]
  wire [7:0] x860_sum_1_io_a; // @[Math.scala 150:24:@39778.4]
  wire [7:0] x860_sum_1_io_b; // @[Math.scala 150:24:@39778.4]
  wire [7:0] x860_sum_1_io_result; // @[Math.scala 150:24:@39778.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@39788.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@39788.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@39788.4]
  wire [7:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@39788.4]
  wire [7:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@39788.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@39797.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@39797.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@39797.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@39797.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@39797.4]
  wire  x866_x17_1_clock; // @[Math.scala 150:24:@39829.4]
  wire  x866_x17_1_reset; // @[Math.scala 150:24:@39829.4]
  wire [7:0] x866_x17_1_io_a; // @[Math.scala 150:24:@39829.4]
  wire [7:0] x866_x17_1_io_b; // @[Math.scala 150:24:@39829.4]
  wire  x866_x17_1_io_flow; // @[Math.scala 150:24:@39829.4]
  wire [7:0] x866_x17_1_io_result; // @[Math.scala 150:24:@39829.4]
  wire  x867_x18_1_clock; // @[Math.scala 150:24:@39839.4]
  wire  x867_x18_1_reset; // @[Math.scala 150:24:@39839.4]
  wire [7:0] x867_x18_1_io_a; // @[Math.scala 150:24:@39839.4]
  wire [7:0] x867_x18_1_io_b; // @[Math.scala 150:24:@39839.4]
  wire  x867_x18_1_io_flow; // @[Math.scala 150:24:@39839.4]
  wire [7:0] x867_x18_1_io_result; // @[Math.scala 150:24:@39839.4]
  wire  x868_x17_1_clock; // @[Math.scala 150:24:@39849.4]
  wire  x868_x17_1_reset; // @[Math.scala 150:24:@39849.4]
  wire [7:0] x868_x17_1_io_a; // @[Math.scala 150:24:@39849.4]
  wire [7:0] x868_x17_1_io_b; // @[Math.scala 150:24:@39849.4]
  wire  x868_x17_1_io_flow; // @[Math.scala 150:24:@39849.4]
  wire [7:0] x868_x17_1_io_result; // @[Math.scala 150:24:@39849.4]
  wire  x869_x18_1_clock; // @[Math.scala 150:24:@39859.4]
  wire  x869_x18_1_reset; // @[Math.scala 150:24:@39859.4]
  wire [7:0] x869_x18_1_io_a; // @[Math.scala 150:24:@39859.4]
  wire [7:0] x869_x18_1_io_b; // @[Math.scala 150:24:@39859.4]
  wire  x869_x18_1_io_flow; // @[Math.scala 150:24:@39859.4]
  wire [7:0] x869_x18_1_io_result; // @[Math.scala 150:24:@39859.4]
  wire [7:0] x870_x17_1_io_a; // @[Math.scala 150:24:@39869.4]
  wire [7:0] x870_x17_1_io_b; // @[Math.scala 150:24:@39869.4]
  wire [7:0] x870_x17_1_io_result; // @[Math.scala 150:24:@39869.4]
  wire [7:0] x871_x18_1_io_a; // @[Math.scala 150:24:@39879.4]
  wire [7:0] x871_x18_1_io_b; // @[Math.scala 150:24:@39879.4]
  wire [7:0] x871_x18_1_io_result; // @[Math.scala 150:24:@39879.4]
  wire [7:0] x872_x17_1_io_a; // @[Math.scala 150:24:@39889.4]
  wire [7:0] x872_x17_1_io_b; // @[Math.scala 150:24:@39889.4]
  wire [7:0] x872_x17_1_io_result; // @[Math.scala 150:24:@39889.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@39899.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@39899.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@39899.4]
  wire [7:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@39899.4]
  wire [7:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@39899.4]
  wire [7:0] x873_sum_1_io_a; // @[Math.scala 150:24:@39908.4]
  wire [7:0] x873_sum_1_io_b; // @[Math.scala 150:24:@39908.4]
  wire [7:0] x873_sum_1_io_result; // @[Math.scala 150:24:@39908.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@39922.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@39922.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@39922.4]
  wire [7:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@39922.4]
  wire [7:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@39922.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@39932.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@39932.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@39932.4]
  wire [7:0] RetimeWrapper_116_io_in; // @[package.scala 93:22:@39932.4]
  wire [7:0] RetimeWrapper_116_io_out; // @[package.scala 93:22:@39932.4]
  wire [7:0] x875_sub_1_io_a; // @[Math.scala 191:24:@39941.4]
  wire [7:0] x875_sub_1_io_b; // @[Math.scala 191:24:@39941.4]
  wire [7:0] x875_sub_1_io_result; // @[Math.scala 191:24:@39941.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@39966.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@39966.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@39966.4]
  wire [7:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@39966.4]
  wire [7:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@39966.4]
  wire  x879_div_1_clock; // @[Math.scala 327:24:@39977.4]
  wire  x879_div_1_reset; // @[Math.scala 327:24:@39977.4]
  wire [7:0] x879_div_1_io_a; // @[Math.scala 327:24:@39977.4]
  wire  x879_div_1_io_flow; // @[Math.scala 327:24:@39977.4]
  wire [7:0] x879_div_1_io_result; // @[Math.scala 327:24:@39977.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@39987.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@39987.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@39987.4]
  wire [7:0] RetimeWrapper_118_io_in; // @[package.scala 93:22:@39987.4]
  wire [7:0] RetimeWrapper_118_io_out; // @[package.scala 93:22:@39987.4]
  wire [7:0] x880_sum_1_io_a; // @[Math.scala 150:24:@39998.4]
  wire [7:0] x880_sum_1_io_b; // @[Math.scala 150:24:@39998.4]
  wire [7:0] x880_sum_1_io_result; // @[Math.scala 150:24:@39998.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@40008.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@40008.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@40008.4]
  wire [7:0] RetimeWrapper_119_io_in; // @[package.scala 93:22:@40008.4]
  wire [7:0] RetimeWrapper_119_io_out; // @[package.scala 93:22:@40008.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@40017.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@40017.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@40017.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@40017.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@40017.4]
  wire  x886_x17_1_clock; // @[Math.scala 150:24:@40049.4]
  wire  x886_x17_1_reset; // @[Math.scala 150:24:@40049.4]
  wire [7:0] x886_x17_1_io_a; // @[Math.scala 150:24:@40049.4]
  wire [7:0] x886_x17_1_io_b; // @[Math.scala 150:24:@40049.4]
  wire  x886_x17_1_io_flow; // @[Math.scala 150:24:@40049.4]
  wire [7:0] x886_x17_1_io_result; // @[Math.scala 150:24:@40049.4]
  wire  x887_x18_1_clock; // @[Math.scala 150:24:@40059.4]
  wire  x887_x18_1_reset; // @[Math.scala 150:24:@40059.4]
  wire [7:0] x887_x18_1_io_a; // @[Math.scala 150:24:@40059.4]
  wire [7:0] x887_x18_1_io_b; // @[Math.scala 150:24:@40059.4]
  wire  x887_x18_1_io_flow; // @[Math.scala 150:24:@40059.4]
  wire [7:0] x887_x18_1_io_result; // @[Math.scala 150:24:@40059.4]
  wire  x888_x17_1_clock; // @[Math.scala 150:24:@40069.4]
  wire  x888_x17_1_reset; // @[Math.scala 150:24:@40069.4]
  wire [7:0] x888_x17_1_io_a; // @[Math.scala 150:24:@40069.4]
  wire [7:0] x888_x17_1_io_b; // @[Math.scala 150:24:@40069.4]
  wire  x888_x17_1_io_flow; // @[Math.scala 150:24:@40069.4]
  wire [7:0] x888_x17_1_io_result; // @[Math.scala 150:24:@40069.4]
  wire  x889_x18_1_clock; // @[Math.scala 150:24:@40079.4]
  wire  x889_x18_1_reset; // @[Math.scala 150:24:@40079.4]
  wire [7:0] x889_x18_1_io_a; // @[Math.scala 150:24:@40079.4]
  wire [7:0] x889_x18_1_io_b; // @[Math.scala 150:24:@40079.4]
  wire  x889_x18_1_io_flow; // @[Math.scala 150:24:@40079.4]
  wire [7:0] x889_x18_1_io_result; // @[Math.scala 150:24:@40079.4]
  wire [7:0] x890_x17_1_io_a; // @[Math.scala 150:24:@40089.4]
  wire [7:0] x890_x17_1_io_b; // @[Math.scala 150:24:@40089.4]
  wire [7:0] x890_x17_1_io_result; // @[Math.scala 150:24:@40089.4]
  wire [7:0] x891_x18_1_io_a; // @[Math.scala 150:24:@40099.4]
  wire [7:0] x891_x18_1_io_b; // @[Math.scala 150:24:@40099.4]
  wire [7:0] x891_x18_1_io_result; // @[Math.scala 150:24:@40099.4]
  wire [7:0] x892_x17_1_io_a; // @[Math.scala 150:24:@40109.4]
  wire [7:0] x892_x17_1_io_b; // @[Math.scala 150:24:@40109.4]
  wire [7:0] x892_x17_1_io_result; // @[Math.scala 150:24:@40109.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@40119.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@40119.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@40119.4]
  wire [7:0] RetimeWrapper_121_io_in; // @[package.scala 93:22:@40119.4]
  wire [7:0] RetimeWrapper_121_io_out; // @[package.scala 93:22:@40119.4]
  wire [7:0] x893_sum_1_io_a; // @[Math.scala 150:24:@40128.4]
  wire [7:0] x893_sum_1_io_b; // @[Math.scala 150:24:@40128.4]
  wire [7:0] x893_sum_1_io_result; // @[Math.scala 150:24:@40128.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@40142.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@40142.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@40142.4]
  wire [7:0] RetimeWrapper_122_io_in; // @[package.scala 93:22:@40142.4]
  wire [7:0] RetimeWrapper_122_io_out; // @[package.scala 93:22:@40142.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@40152.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@40152.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@40152.4]
  wire [7:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@40152.4]
  wire [7:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@40152.4]
  wire [7:0] x895_sub_1_io_a; // @[Math.scala 191:24:@40161.4]
  wire [7:0] x895_sub_1_io_b; // @[Math.scala 191:24:@40161.4]
  wire [7:0] x895_sub_1_io_result; // @[Math.scala 191:24:@40161.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@40186.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@40186.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@40186.4]
  wire [7:0] RetimeWrapper_124_io_in; // @[package.scala 93:22:@40186.4]
  wire [7:0] RetimeWrapper_124_io_out; // @[package.scala 93:22:@40186.4]
  wire  x899_div_1_clock; // @[Math.scala 327:24:@40197.4]
  wire  x899_div_1_reset; // @[Math.scala 327:24:@40197.4]
  wire [7:0] x899_div_1_io_a; // @[Math.scala 327:24:@40197.4]
  wire  x899_div_1_io_flow; // @[Math.scala 327:24:@40197.4]
  wire [7:0] x899_div_1_io_result; // @[Math.scala 327:24:@40197.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@40207.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@40207.4]
  wire [7:0] RetimeWrapper_125_io_in; // @[package.scala 93:22:@40207.4]
  wire [7:0] RetimeWrapper_125_io_out; // @[package.scala 93:22:@40207.4]
  wire [7:0] x900_sum_1_io_a; // @[Math.scala 150:24:@40216.4]
  wire [7:0] x900_sum_1_io_b; // @[Math.scala 150:24:@40216.4]
  wire [7:0] x900_sum_1_io_result; // @[Math.scala 150:24:@40216.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@40226.4]
  wire [7:0] RetimeWrapper_126_io_in; // @[package.scala 93:22:@40226.4]
  wire [7:0] RetimeWrapper_126_io_out; // @[package.scala 93:22:@40226.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@40235.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@40235.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@40235.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@40235.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@40235.4]
  wire  x905_x17_1_clock; // @[Math.scala 150:24:@40262.4]
  wire  x905_x17_1_reset; // @[Math.scala 150:24:@40262.4]
  wire [7:0] x905_x17_1_io_a; // @[Math.scala 150:24:@40262.4]
  wire [7:0] x905_x17_1_io_b; // @[Math.scala 150:24:@40262.4]
  wire  x905_x17_1_io_flow; // @[Math.scala 150:24:@40262.4]
  wire [7:0] x905_x17_1_io_result; // @[Math.scala 150:24:@40262.4]
  wire  x906_x18_1_clock; // @[Math.scala 150:24:@40272.4]
  wire  x906_x18_1_reset; // @[Math.scala 150:24:@40272.4]
  wire [7:0] x906_x18_1_io_a; // @[Math.scala 150:24:@40272.4]
  wire [7:0] x906_x18_1_io_b; // @[Math.scala 150:24:@40272.4]
  wire  x906_x18_1_io_flow; // @[Math.scala 150:24:@40272.4]
  wire [7:0] x906_x18_1_io_result; // @[Math.scala 150:24:@40272.4]
  wire  x907_x17_1_clock; // @[Math.scala 150:24:@40282.4]
  wire  x907_x17_1_reset; // @[Math.scala 150:24:@40282.4]
  wire [7:0] x907_x17_1_io_a; // @[Math.scala 150:24:@40282.4]
  wire [7:0] x907_x17_1_io_b; // @[Math.scala 150:24:@40282.4]
  wire  x907_x17_1_io_flow; // @[Math.scala 150:24:@40282.4]
  wire [7:0] x907_x17_1_io_result; // @[Math.scala 150:24:@40282.4]
  wire  x908_x18_1_clock; // @[Math.scala 150:24:@40292.4]
  wire  x908_x18_1_reset; // @[Math.scala 150:24:@40292.4]
  wire [7:0] x908_x18_1_io_a; // @[Math.scala 150:24:@40292.4]
  wire [7:0] x908_x18_1_io_b; // @[Math.scala 150:24:@40292.4]
  wire  x908_x18_1_io_flow; // @[Math.scala 150:24:@40292.4]
  wire [7:0] x908_x18_1_io_result; // @[Math.scala 150:24:@40292.4]
  wire [7:0] x909_x17_1_io_a; // @[Math.scala 150:24:@40302.4]
  wire [7:0] x909_x17_1_io_b; // @[Math.scala 150:24:@40302.4]
  wire [7:0] x909_x17_1_io_result; // @[Math.scala 150:24:@40302.4]
  wire [7:0] x910_x18_1_io_a; // @[Math.scala 150:24:@40312.4]
  wire [7:0] x910_x18_1_io_b; // @[Math.scala 150:24:@40312.4]
  wire [7:0] x910_x18_1_io_result; // @[Math.scala 150:24:@40312.4]
  wire [7:0] x911_x17_1_io_a; // @[Math.scala 150:24:@40322.4]
  wire [7:0] x911_x17_1_io_b; // @[Math.scala 150:24:@40322.4]
  wire [7:0] x911_x17_1_io_result; // @[Math.scala 150:24:@40322.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@40332.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@40332.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@40332.4]
  wire [7:0] RetimeWrapper_128_io_in; // @[package.scala 93:22:@40332.4]
  wire [7:0] RetimeWrapper_128_io_out; // @[package.scala 93:22:@40332.4]
  wire [7:0] x912_sum_1_io_a; // @[Math.scala 150:24:@40341.4]
  wire [7:0] x912_sum_1_io_b; // @[Math.scala 150:24:@40341.4]
  wire [7:0] x912_sum_1_io_result; // @[Math.scala 150:24:@40341.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@40355.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@40355.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@40355.4]
  wire [7:0] RetimeWrapper_129_io_in; // @[package.scala 93:22:@40355.4]
  wire [7:0] RetimeWrapper_129_io_out; // @[package.scala 93:22:@40355.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@40365.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@40365.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@40365.4]
  wire [7:0] RetimeWrapper_130_io_in; // @[package.scala 93:22:@40365.4]
  wire [7:0] RetimeWrapper_130_io_out; // @[package.scala 93:22:@40365.4]
  wire [7:0] x914_sub_1_io_a; // @[Math.scala 191:24:@40374.4]
  wire [7:0] x914_sub_1_io_b; // @[Math.scala 191:24:@40374.4]
  wire [7:0] x914_sub_1_io_result; // @[Math.scala 191:24:@40374.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@40399.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@40399.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@40399.4]
  wire [7:0] RetimeWrapper_131_io_in; // @[package.scala 93:22:@40399.4]
  wire [7:0] RetimeWrapper_131_io_out; // @[package.scala 93:22:@40399.4]
  wire  x918_div_1_clock; // @[Math.scala 327:24:@40412.4]
  wire  x918_div_1_reset; // @[Math.scala 327:24:@40412.4]
  wire [7:0] x918_div_1_io_a; // @[Math.scala 327:24:@40412.4]
  wire  x918_div_1_io_flow; // @[Math.scala 327:24:@40412.4]
  wire [7:0] x918_div_1_io_result; // @[Math.scala 327:24:@40412.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@40422.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@40422.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@40422.4]
  wire [7:0] RetimeWrapper_132_io_in; // @[package.scala 93:22:@40422.4]
  wire [7:0] RetimeWrapper_132_io_out; // @[package.scala 93:22:@40422.4]
  wire [7:0] x919_sum_1_io_a; // @[Math.scala 150:24:@40431.4]
  wire [7:0] x919_sum_1_io_b; // @[Math.scala 150:24:@40431.4]
  wire [7:0] x919_sum_1_io_result; // @[Math.scala 150:24:@40431.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@40441.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@40441.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@40441.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@40441.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@40441.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@40450.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@40450.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@40450.4]
  wire [7:0] RetimeWrapper_134_io_in; // @[package.scala 93:22:@40450.4]
  wire [7:0] RetimeWrapper_134_io_out; // @[package.scala 93:22:@40450.4]
  wire  x923_x17_1_clock; // @[Math.scala 150:24:@40472.4]
  wire  x923_x17_1_reset; // @[Math.scala 150:24:@40472.4]
  wire [7:0] x923_x17_1_io_a; // @[Math.scala 150:24:@40472.4]
  wire [7:0] x923_x17_1_io_b; // @[Math.scala 150:24:@40472.4]
  wire  x923_x17_1_io_flow; // @[Math.scala 150:24:@40472.4]
  wire [7:0] x923_x17_1_io_result; // @[Math.scala 150:24:@40472.4]
  wire  x924_x18_1_clock; // @[Math.scala 150:24:@40482.4]
  wire  x924_x18_1_reset; // @[Math.scala 150:24:@40482.4]
  wire [7:0] x924_x18_1_io_a; // @[Math.scala 150:24:@40482.4]
  wire [7:0] x924_x18_1_io_b; // @[Math.scala 150:24:@40482.4]
  wire  x924_x18_1_io_flow; // @[Math.scala 150:24:@40482.4]
  wire [7:0] x924_x18_1_io_result; // @[Math.scala 150:24:@40482.4]
  wire  x925_x17_1_clock; // @[Math.scala 150:24:@40492.4]
  wire  x925_x17_1_reset; // @[Math.scala 150:24:@40492.4]
  wire [7:0] x925_x17_1_io_a; // @[Math.scala 150:24:@40492.4]
  wire [7:0] x925_x17_1_io_b; // @[Math.scala 150:24:@40492.4]
  wire  x925_x17_1_io_flow; // @[Math.scala 150:24:@40492.4]
  wire [7:0] x925_x17_1_io_result; // @[Math.scala 150:24:@40492.4]
  wire  x926_x18_1_clock; // @[Math.scala 150:24:@40502.4]
  wire  x926_x18_1_reset; // @[Math.scala 150:24:@40502.4]
  wire [7:0] x926_x18_1_io_a; // @[Math.scala 150:24:@40502.4]
  wire [7:0] x926_x18_1_io_b; // @[Math.scala 150:24:@40502.4]
  wire  x926_x18_1_io_flow; // @[Math.scala 150:24:@40502.4]
  wire [7:0] x926_x18_1_io_result; // @[Math.scala 150:24:@40502.4]
  wire [7:0] x927_x17_1_io_a; // @[Math.scala 150:24:@40512.4]
  wire [7:0] x927_x17_1_io_b; // @[Math.scala 150:24:@40512.4]
  wire [7:0] x927_x17_1_io_result; // @[Math.scala 150:24:@40512.4]
  wire [7:0] x928_x18_1_io_a; // @[Math.scala 150:24:@40522.4]
  wire [7:0] x928_x18_1_io_b; // @[Math.scala 150:24:@40522.4]
  wire [7:0] x928_x18_1_io_result; // @[Math.scala 150:24:@40522.4]
  wire [7:0] x929_x17_1_io_a; // @[Math.scala 150:24:@40532.4]
  wire [7:0] x929_x17_1_io_b; // @[Math.scala 150:24:@40532.4]
  wire [7:0] x929_x17_1_io_result; // @[Math.scala 150:24:@40532.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@40542.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@40542.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@40542.4]
  wire [7:0] RetimeWrapper_135_io_in; // @[package.scala 93:22:@40542.4]
  wire [7:0] RetimeWrapper_135_io_out; // @[package.scala 93:22:@40542.4]
  wire [7:0] x930_sum_1_io_a; // @[Math.scala 150:24:@40551.4]
  wire [7:0] x930_sum_1_io_b; // @[Math.scala 150:24:@40551.4]
  wire [7:0] x930_sum_1_io_result; // @[Math.scala 150:24:@40551.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@40565.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@40565.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@40565.4]
  wire [7:0] RetimeWrapper_136_io_in; // @[package.scala 93:22:@40565.4]
  wire [7:0] RetimeWrapper_136_io_out; // @[package.scala 93:22:@40565.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@40575.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@40575.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@40575.4]
  wire [7:0] RetimeWrapper_137_io_in; // @[package.scala 93:22:@40575.4]
  wire [7:0] RetimeWrapper_137_io_out; // @[package.scala 93:22:@40575.4]
  wire [7:0] x932_sub_1_io_a; // @[Math.scala 191:24:@40584.4]
  wire [7:0] x932_sub_1_io_b; // @[Math.scala 191:24:@40584.4]
  wire [7:0] x932_sub_1_io_result; // @[Math.scala 191:24:@40584.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@40609.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@40609.4]
  wire [7:0] RetimeWrapper_138_io_in; // @[package.scala 93:22:@40609.4]
  wire [7:0] RetimeWrapper_138_io_out; // @[package.scala 93:22:@40609.4]
  wire  x936_div_1_clock; // @[Math.scala 327:24:@40620.4]
  wire  x936_div_1_reset; // @[Math.scala 327:24:@40620.4]
  wire [7:0] x936_div_1_io_a; // @[Math.scala 327:24:@40620.4]
  wire  x936_div_1_io_flow; // @[Math.scala 327:24:@40620.4]
  wire [7:0] x936_div_1_io_result; // @[Math.scala 327:24:@40620.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@40630.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@40630.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@40630.4]
  wire [7:0] RetimeWrapper_139_io_in; // @[package.scala 93:22:@40630.4]
  wire [7:0] RetimeWrapper_139_io_out; // @[package.scala 93:22:@40630.4]
  wire [7:0] x937_sum_1_io_a; // @[Math.scala 150:24:@40639.4]
  wire [7:0] x937_sum_1_io_b; // @[Math.scala 150:24:@40639.4]
  wire [7:0] x937_sum_1_io_result; // @[Math.scala 150:24:@40639.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@40649.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@40649.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@40649.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@40649.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@40649.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@40658.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@40658.4]
  wire [7:0] RetimeWrapper_141_io_in; // @[package.scala 93:22:@40658.4]
  wire [7:0] RetimeWrapper_141_io_out; // @[package.scala 93:22:@40658.4]
  wire  x941_x17_1_clock; // @[Math.scala 150:24:@40680.4]
  wire  x941_x17_1_reset; // @[Math.scala 150:24:@40680.4]
  wire [7:0] x941_x17_1_io_a; // @[Math.scala 150:24:@40680.4]
  wire [7:0] x941_x17_1_io_b; // @[Math.scala 150:24:@40680.4]
  wire  x941_x17_1_io_flow; // @[Math.scala 150:24:@40680.4]
  wire [7:0] x941_x17_1_io_result; // @[Math.scala 150:24:@40680.4]
  wire  x942_x18_1_clock; // @[Math.scala 150:24:@40690.4]
  wire  x942_x18_1_reset; // @[Math.scala 150:24:@40690.4]
  wire [7:0] x942_x18_1_io_a; // @[Math.scala 150:24:@40690.4]
  wire [7:0] x942_x18_1_io_b; // @[Math.scala 150:24:@40690.4]
  wire  x942_x18_1_io_flow; // @[Math.scala 150:24:@40690.4]
  wire [7:0] x942_x18_1_io_result; // @[Math.scala 150:24:@40690.4]
  wire  x943_x17_1_clock; // @[Math.scala 150:24:@40700.4]
  wire  x943_x17_1_reset; // @[Math.scala 150:24:@40700.4]
  wire [7:0] x943_x17_1_io_a; // @[Math.scala 150:24:@40700.4]
  wire [7:0] x943_x17_1_io_b; // @[Math.scala 150:24:@40700.4]
  wire  x943_x17_1_io_flow; // @[Math.scala 150:24:@40700.4]
  wire [7:0] x943_x17_1_io_result; // @[Math.scala 150:24:@40700.4]
  wire  x944_x18_1_clock; // @[Math.scala 150:24:@40710.4]
  wire  x944_x18_1_reset; // @[Math.scala 150:24:@40710.4]
  wire [7:0] x944_x18_1_io_a; // @[Math.scala 150:24:@40710.4]
  wire [7:0] x944_x18_1_io_b; // @[Math.scala 150:24:@40710.4]
  wire  x944_x18_1_io_flow; // @[Math.scala 150:24:@40710.4]
  wire [7:0] x944_x18_1_io_result; // @[Math.scala 150:24:@40710.4]
  wire [7:0] x945_x17_1_io_a; // @[Math.scala 150:24:@40720.4]
  wire [7:0] x945_x17_1_io_b; // @[Math.scala 150:24:@40720.4]
  wire [7:0] x945_x17_1_io_result; // @[Math.scala 150:24:@40720.4]
  wire [7:0] x946_x18_1_io_a; // @[Math.scala 150:24:@40730.4]
  wire [7:0] x946_x18_1_io_b; // @[Math.scala 150:24:@40730.4]
  wire [7:0] x946_x18_1_io_result; // @[Math.scala 150:24:@40730.4]
  wire [7:0] x947_x17_1_io_a; // @[Math.scala 150:24:@40740.4]
  wire [7:0] x947_x17_1_io_b; // @[Math.scala 150:24:@40740.4]
  wire [7:0] x947_x17_1_io_result; // @[Math.scala 150:24:@40740.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@40750.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@40750.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@40750.4]
  wire [7:0] RetimeWrapper_142_io_in; // @[package.scala 93:22:@40750.4]
  wire [7:0] RetimeWrapper_142_io_out; // @[package.scala 93:22:@40750.4]
  wire [7:0] x948_sum_1_io_a; // @[Math.scala 150:24:@40759.4]
  wire [7:0] x948_sum_1_io_b; // @[Math.scala 150:24:@40759.4]
  wire [7:0] x948_sum_1_io_result; // @[Math.scala 150:24:@40759.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@40773.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@40773.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@40773.4]
  wire [7:0] RetimeWrapper_143_io_in; // @[package.scala 93:22:@40773.4]
  wire [7:0] RetimeWrapper_143_io_out; // @[package.scala 93:22:@40773.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@40783.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@40783.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@40783.4]
  wire [7:0] RetimeWrapper_144_io_in; // @[package.scala 93:22:@40783.4]
  wire [7:0] RetimeWrapper_144_io_out; // @[package.scala 93:22:@40783.4]
  wire [7:0] x950_sub_1_io_a; // @[Math.scala 191:24:@40792.4]
  wire [7:0] x950_sub_1_io_b; // @[Math.scala 191:24:@40792.4]
  wire [7:0] x950_sub_1_io_result; // @[Math.scala 191:24:@40792.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@40817.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@40817.4]
  wire [7:0] RetimeWrapper_145_io_in; // @[package.scala 93:22:@40817.4]
  wire [7:0] RetimeWrapper_145_io_out; // @[package.scala 93:22:@40817.4]
  wire  x954_div_1_clock; // @[Math.scala 327:24:@40828.4]
  wire  x954_div_1_reset; // @[Math.scala 327:24:@40828.4]
  wire [7:0] x954_div_1_io_a; // @[Math.scala 327:24:@40828.4]
  wire  x954_div_1_io_flow; // @[Math.scala 327:24:@40828.4]
  wire [7:0] x954_div_1_io_result; // @[Math.scala 327:24:@40828.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@40838.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@40838.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@40838.4]
  wire [7:0] RetimeWrapper_146_io_in; // @[package.scala 93:22:@40838.4]
  wire [7:0] RetimeWrapper_146_io_out; // @[package.scala 93:22:@40838.4]
  wire [7:0] x955_sum_1_io_a; // @[Math.scala 150:24:@40849.4]
  wire [7:0] x955_sum_1_io_b; // @[Math.scala 150:24:@40849.4]
  wire [7:0] x955_sum_1_io_result; // @[Math.scala 150:24:@40849.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@40859.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@40859.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@40859.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@40859.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@40859.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@40868.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@40868.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@40868.4]
  wire [7:0] RetimeWrapper_148_io_in; // @[package.scala 93:22:@40868.4]
  wire [7:0] RetimeWrapper_148_io_out; // @[package.scala 93:22:@40868.4]
  wire  x960_x17_1_clock; // @[Math.scala 150:24:@40895.4]
  wire  x960_x17_1_reset; // @[Math.scala 150:24:@40895.4]
  wire [7:0] x960_x17_1_io_a; // @[Math.scala 150:24:@40895.4]
  wire [7:0] x960_x17_1_io_b; // @[Math.scala 150:24:@40895.4]
  wire  x960_x17_1_io_flow; // @[Math.scala 150:24:@40895.4]
  wire [7:0] x960_x17_1_io_result; // @[Math.scala 150:24:@40895.4]
  wire  x961_x18_1_clock; // @[Math.scala 150:24:@40905.4]
  wire  x961_x18_1_reset; // @[Math.scala 150:24:@40905.4]
  wire [7:0] x961_x18_1_io_a; // @[Math.scala 150:24:@40905.4]
  wire [7:0] x961_x18_1_io_b; // @[Math.scala 150:24:@40905.4]
  wire  x961_x18_1_io_flow; // @[Math.scala 150:24:@40905.4]
  wire [7:0] x961_x18_1_io_result; // @[Math.scala 150:24:@40905.4]
  wire  x962_x17_1_clock; // @[Math.scala 150:24:@40915.4]
  wire  x962_x17_1_reset; // @[Math.scala 150:24:@40915.4]
  wire [7:0] x962_x17_1_io_a; // @[Math.scala 150:24:@40915.4]
  wire [7:0] x962_x17_1_io_b; // @[Math.scala 150:24:@40915.4]
  wire  x962_x17_1_io_flow; // @[Math.scala 150:24:@40915.4]
  wire [7:0] x962_x17_1_io_result; // @[Math.scala 150:24:@40915.4]
  wire  x963_x18_1_clock; // @[Math.scala 150:24:@40925.4]
  wire  x963_x18_1_reset; // @[Math.scala 150:24:@40925.4]
  wire [7:0] x963_x18_1_io_a; // @[Math.scala 150:24:@40925.4]
  wire [7:0] x963_x18_1_io_b; // @[Math.scala 150:24:@40925.4]
  wire  x963_x18_1_io_flow; // @[Math.scala 150:24:@40925.4]
  wire [7:0] x963_x18_1_io_result; // @[Math.scala 150:24:@40925.4]
  wire [7:0] x964_x17_1_io_a; // @[Math.scala 150:24:@40935.4]
  wire [7:0] x964_x17_1_io_b; // @[Math.scala 150:24:@40935.4]
  wire [7:0] x964_x17_1_io_result; // @[Math.scala 150:24:@40935.4]
  wire [7:0] x965_x18_1_io_a; // @[Math.scala 150:24:@40945.4]
  wire [7:0] x965_x18_1_io_b; // @[Math.scala 150:24:@40945.4]
  wire [7:0] x965_x18_1_io_result; // @[Math.scala 150:24:@40945.4]
  wire [7:0] x966_x17_1_io_a; // @[Math.scala 150:24:@40955.4]
  wire [7:0] x966_x17_1_io_b; // @[Math.scala 150:24:@40955.4]
  wire [7:0] x966_x17_1_io_result; // @[Math.scala 150:24:@40955.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@40965.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@40965.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@40965.4]
  wire [7:0] RetimeWrapper_149_io_in; // @[package.scala 93:22:@40965.4]
  wire [7:0] RetimeWrapper_149_io_out; // @[package.scala 93:22:@40965.4]
  wire [7:0] x967_sum_1_io_a; // @[Math.scala 150:24:@40974.4]
  wire [7:0] x967_sum_1_io_b; // @[Math.scala 150:24:@40974.4]
  wire [7:0] x967_sum_1_io_result; // @[Math.scala 150:24:@40974.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@40988.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@40988.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@40988.4]
  wire [7:0] RetimeWrapper_150_io_in; // @[package.scala 93:22:@40988.4]
  wire [7:0] RetimeWrapper_150_io_out; // @[package.scala 93:22:@40988.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@40998.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@40998.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@40998.4]
  wire [7:0] RetimeWrapper_151_io_in; // @[package.scala 93:22:@40998.4]
  wire [7:0] RetimeWrapper_151_io_out; // @[package.scala 93:22:@40998.4]
  wire [7:0] x969_sub_1_io_a; // @[Math.scala 191:24:@41007.4]
  wire [7:0] x969_sub_1_io_b; // @[Math.scala 191:24:@41007.4]
  wire [7:0] x969_sub_1_io_result; // @[Math.scala 191:24:@41007.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@41032.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@41032.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@41032.4]
  wire [7:0] RetimeWrapper_152_io_in; // @[package.scala 93:22:@41032.4]
  wire [7:0] RetimeWrapper_152_io_out; // @[package.scala 93:22:@41032.4]
  wire  x973_div_1_clock; // @[Math.scala 327:24:@41043.4]
  wire  x973_div_1_reset; // @[Math.scala 327:24:@41043.4]
  wire [7:0] x973_div_1_io_a; // @[Math.scala 327:24:@41043.4]
  wire  x973_div_1_io_flow; // @[Math.scala 327:24:@41043.4]
  wire [7:0] x973_div_1_io_result; // @[Math.scala 327:24:@41043.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@41053.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@41053.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@41053.4]
  wire [7:0] RetimeWrapper_153_io_in; // @[package.scala 93:22:@41053.4]
  wire [7:0] RetimeWrapper_153_io_out; // @[package.scala 93:22:@41053.4]
  wire [7:0] x974_sum_1_io_a; // @[Math.scala 150:24:@41062.4]
  wire [7:0] x974_sum_1_io_b; // @[Math.scala 150:24:@41062.4]
  wire [7:0] x974_sum_1_io_result; // @[Math.scala 150:24:@41062.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@41072.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@41072.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@41072.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@41072.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@41072.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@41081.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@41081.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@41081.4]
  wire [7:0] RetimeWrapper_155_io_in; // @[package.scala 93:22:@41081.4]
  wire [7:0] RetimeWrapper_155_io_out; // @[package.scala 93:22:@41081.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@41111.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@41111.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@41111.4]
  wire [63:0] RetimeWrapper_156_io_in; // @[package.scala 93:22:@41111.4]
  wire [63:0] RetimeWrapper_156_io_out; // @[package.scala 93:22:@41111.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@41120.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@41120.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@41120.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@41120.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@41120.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@41129.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@41129.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@41129.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@41129.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@41129.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@41138.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@41138.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@41138.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@41138.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@41138.4]
  wire  b537; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 62:18:@36708.4]
  wire  b538; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 63:18:@36709.4]
  wire  _T_206; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 68:30:@36924.4]
  wire  _T_207; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 68:37:@36925.4]
  wire  _T_211; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:76:@36930.4]
  wire  _T_212; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:62:@36931.4]
  wire  _T_214; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:101:@36932.4]
  wire [63:0] x1058_x540_D1_0_number; // @[package.scala 96:25:@36941.4 package.scala 96:25:@36942.4]
  wire [31:0] b535_number; // @[Math.scala 712:22:@36693.4 Math.scala 713:14:@36694.4]
  wire [31:0] _T_254; // @[Math.scala 499:52:@36969.4]
  wire  x544; // @[Math.scala 499:44:@36977.4]
  wire  x545; // @[Math.scala 499:44:@36984.4]
  wire  x546; // @[Math.scala 499:44:@36991.4]
  wire [31:0] _T_301; // @[Mux.scala 19:72:@37003.4]
  wire [31:0] _T_303; // @[Mux.scala 19:72:@37004.4]
  wire [31:0] _T_305; // @[Mux.scala 19:72:@37005.4]
  wire [31:0] _T_307; // @[Mux.scala 19:72:@37007.4]
  wire [31:0] x547_number; // @[Mux.scala 19:72:@37008.4]
  wire [31:0] _T_319; // @[Math.scala 406:49:@37018.4]
  wire [31:0] _T_321; // @[Math.scala 406:56:@37020.4]
  wire [31:0] _T_322; // @[Math.scala 406:56:@37021.4]
  wire  _T_327; // @[FixedPoint.scala 50:25:@37027.4]
  wire [1:0] _T_331; // @[Bitwise.scala 72:12:@37029.4]
  wire [29:0] _T_332; // @[FixedPoint.scala 18:52:@37030.4]
  wire [31:0] b536_number; // @[Math.scala 712:22:@36705.4 Math.scala 713:14:@36706.4]
  wire  _T_337; // @[FixedPoint.scala 50:25:@37036.4]
  wire [1:0] _T_341; // @[Bitwise.scala 72:12:@37038.4]
  wire [29:0] _T_342; // @[FixedPoint.scala 18:52:@37039.4]
  wire  _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:101:@37100.4]
  wire  _T_371; // @[package.scala 96:25:@37108.4 package.scala 96:25:@37109.4]
  wire  _T_373; // @[implicits.scala 55:10:@37110.4]
  wire  _T_374; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:118:@37111.4]
  wire  _T_376; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:205:@37113.4]
  wire  _T_377; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:224:@37114.4]
  wire  x1060_b537_D8; // @[package.scala 96:25:@37068.4 package.scala 96:25:@37069.4]
  wire  _T_378; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:250:@37115.4]
  wire  x1059_b538_D8; // @[package.scala 96:25:@37059.4 package.scala 96:25:@37060.4]
  wire [31:0] x559_rdcol_number; // @[Math.scala 154:22:@37132.4 Math.scala 155:14:@37133.4]
  wire  _T_391; // @[FixedPoint.scala 50:25:@37139.4]
  wire [1:0] _T_395; // @[Bitwise.scala 72:12:@37141.4]
  wire [29:0] _T_396; // @[FixedPoint.scala 18:52:@37142.4]
  wire  _T_419; // @[package.scala 96:25:@37193.4 package.scala 96:25:@37194.4]
  wire  _T_421; // @[implicits.scala 55:10:@37195.4]
  wire  _T_422; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:118:@37196.4]
  wire  _T_424; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:205:@37198.4]
  wire  _T_425; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:224:@37199.4]
  wire  _T_426; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:250:@37200.4]
  wire [31:0] x568_rdcol_number; // @[Math.scala 154:22:@37217.4 Math.scala 155:14:@37218.4]
  wire  _T_439; // @[FixedPoint.scala 50:25:@37224.4]
  wire [1:0] _T_443; // @[Bitwise.scala 72:12:@37226.4]
  wire [29:0] _T_444; // @[FixedPoint.scala 18:52:@37227.4]
  wire  _T_464; // @[package.scala 96:25:@37269.4 package.scala 96:25:@37270.4]
  wire  _T_466; // @[implicits.scala 55:10:@37271.4]
  wire  _T_467; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:118:@37272.4]
  wire  _T_469; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:205:@37274.4]
  wire  _T_470; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:224:@37275.4]
  wire  _T_471; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:250:@37276.4]
  wire [31:0] x577_rdcol_number; // @[Math.scala 154:22:@37293.4 Math.scala 155:14:@37294.4]
  wire  _T_484; // @[FixedPoint.scala 50:25:@37300.4]
  wire [1:0] _T_488; // @[Bitwise.scala 72:12:@37302.4]
  wire [29:0] _T_489; // @[FixedPoint.scala 18:52:@37303.4]
  wire  _T_509; // @[package.scala 96:25:@37345.4 package.scala 96:25:@37346.4]
  wire  _T_511; // @[implicits.scala 55:10:@37347.4]
  wire  _T_512; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:118:@37348.4]
  wire  _T_514; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:205:@37350.4]
  wire  _T_515; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:224:@37351.4]
  wire  _T_516; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:250:@37352.4]
  wire [31:0] x586_rdrow_number; // @[Math.scala 154:22:@37369.4 Math.scala 155:14:@37370.4]
  wire [31:0] _T_531; // @[Math.scala 499:52:@37376.4]
  wire  x588; // @[Math.scala 499:44:@37384.4]
  wire  x589; // @[Math.scala 499:44:@37391.4]
  wire  x590; // @[Math.scala 499:44:@37398.4]
  wire [31:0] _T_578; // @[Mux.scala 19:72:@37410.4]
  wire [31:0] _T_580; // @[Mux.scala 19:72:@37411.4]
  wire [31:0] _T_582; // @[Mux.scala 19:72:@37412.4]
  wire [31:0] _T_584; // @[Mux.scala 19:72:@37414.4]
  wire [31:0] x591_number; // @[Mux.scala 19:72:@37415.4]
  wire [31:0] _T_598; // @[Math.scala 406:49:@37427.4]
  wire [31:0] _T_600; // @[Math.scala 406:56:@37429.4]
  wire [31:0] _T_601; // @[Math.scala 406:56:@37430.4]
  wire  _T_606; // @[FixedPoint.scala 50:25:@37436.4]
  wire [1:0] _T_610; // @[Bitwise.scala 72:12:@37438.4]
  wire [29:0] _T_611; // @[FixedPoint.scala 18:52:@37439.4]
  wire  _T_637; // @[package.scala 96:25:@37499.4 package.scala 96:25:@37500.4]
  wire  _T_639; // @[implicits.scala 55:10:@37501.4]
  wire  _T_640; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:166:@37502.4]
  wire  _T_642; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:253:@37504.4]
  wire  _T_643; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:272:@37505.4]
  wire  _T_644; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:298:@37506.4]
  wire  _T_665; // @[package.scala 96:25:@37554.4 package.scala 96:25:@37555.4]
  wire  _T_667; // @[implicits.scala 55:10:@37556.4]
  wire  _T_668; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:166:@37557.4]
  wire  _T_670; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:253:@37559.4]
  wire  _T_671; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:272:@37560.4]
  wire  _T_672; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:298:@37561.4]
  wire  _T_693; // @[package.scala 96:25:@37609.4 package.scala 96:25:@37610.4]
  wire  _T_695; // @[implicits.scala 55:10:@37611.4]
  wire  _T_696; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:166:@37612.4]
  wire  _T_698; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:253:@37614.4]
  wire  _T_699; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:272:@37615.4]
  wire  _T_700; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:298:@37616.4]
  wire  _T_721; // @[package.scala 96:25:@37664.4 package.scala 96:25:@37665.4]
  wire  _T_723; // @[implicits.scala 55:10:@37666.4]
  wire  _T_724; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:166:@37667.4]
  wire  _T_726; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:253:@37669.4]
  wire  _T_727; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:272:@37670.4]
  wire  _T_728; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:298:@37671.4]
  wire [31:0] x1081_x586_rdrow_D11_number; // @[package.scala 96:25:@37685.4 package.scala 96:25:@37686.4]
  wire [31:0] _T_740; // @[Math.scala 406:49:@37692.4]
  wire [31:0] _T_742; // @[Math.scala 406:56:@37694.4]
  wire [31:0] _T_743; // @[Math.scala 406:56:@37695.4]
  wire [31:0] x1050_number; // @[implicits.scala 133:21:@37696.4]
  wire  x617; // @[Math.scala 465:44:@37704.4]
  wire [31:0] x1082_x577_rdcol_D11_number; // @[package.scala 96:25:@37712.4 package.scala 96:25:@37713.4]
  wire [31:0] _T_761; // @[Math.scala 465:37:@37718.4]
  wire  x618; // @[Math.scala 465:44:@37720.4]
  wire  x619; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 259:24:@37723.4]
  wire [31:0] _T_775; // @[Math.scala 406:49:@37732.4]
  wire [31:0] _T_777; // @[Math.scala 406:56:@37734.4]
  wire [31:0] _T_778; // @[Math.scala 406:56:@37735.4]
  wire  _T_783; // @[FixedPoint.scala 50:25:@37741.4]
  wire [1:0] _T_787; // @[Bitwise.scala 72:12:@37743.4]
  wire [29:0] _T_788; // @[FixedPoint.scala 18:52:@37744.4]
  wire  _T_823; // @[package.scala 96:25:@37814.4 package.scala 96:25:@37815.4]
  wire  _T_825; // @[implicits.scala 55:10:@37816.4]
  wire  _T_826; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 282:194:@37817.4]
  wire  x1087_x620_D1; // @[package.scala 96:25:@37800.4 package.scala 96:25:@37801.4]
  wire  _T_827; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 282:282:@37818.4]
  wire  x1086_b537_D13; // @[package.scala 96:25:@37791.4 package.scala 96:25:@37792.4]
  wire  _T_828; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 282:291:@37819.4]
  wire  x1084_b538_D13; // @[package.scala 96:25:@37773.4 package.scala 96:25:@37774.4]
  wire [31:0] x1088_x568_rdcol_D11_number; // @[package.scala 96:25:@37835.4 package.scala 96:25:@37836.4]
  wire [31:0] _T_839; // @[Math.scala 465:37:@37841.4]
  wire  x629; // @[Math.scala 465:44:@37843.4]
  wire  x630; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 290:24:@37846.4]
  wire  _T_870; // @[package.scala 96:25:@37890.4 package.scala 96:25:@37891.4]
  wire  _T_872; // @[implicits.scala 55:10:@37892.4]
  wire  _T_873; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:194:@37893.4]
  wire  x1090_x631_D1; // @[package.scala 96:25:@37876.4 package.scala 96:25:@37877.4]
  wire  _T_874; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:282:@37894.4]
  wire  _T_875; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:326:@37895.4]
  wire [31:0] x1091_x559_rdcol_D11_number; // @[package.scala 96:25:@37911.4 package.scala 96:25:@37912.4]
  wire [31:0] _T_888; // @[Math.scala 465:37:@37919.4]
  wire  x637; // @[Math.scala 465:44:@37921.4]
  wire  x638; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 319:59:@37924.4]
  wire  _T_919; // @[package.scala 96:25:@37968.4 package.scala 96:25:@37969.4]
  wire  _T_921; // @[implicits.scala 55:10:@37970.4]
  wire  _T_922; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:194:@37971.4]
  wire  x1093_x639_D1; // @[package.scala 96:25:@37954.4 package.scala 96:25:@37955.4]
  wire  _T_923; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:282:@37972.4]
  wire  _T_924; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:291:@37973.4]
  wire [31:0] x1094_b536_D11_number; // @[package.scala 96:25:@37989.4 package.scala 96:25:@37990.4]
  wire [31:0] _T_935; // @[Math.scala 465:37:@37995.4]
  wire  x645; // @[Math.scala 465:44:@37997.4]
  wire  x1095_x645_D1; // @[package.scala 96:25:@38005.4 package.scala 96:25:@38006.4]
  wire  x646; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 342:59:@38009.4]
  wire  _T_969; // @[package.scala 96:25:@38053.4 package.scala 96:25:@38054.4]
  wire  _T_971; // @[implicits.scala 55:10:@38055.4]
  wire  _T_972; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:194:@38056.4]
  wire  x1097_x647_D1; // @[package.scala 96:25:@38039.4 package.scala 96:25:@38040.4]
  wire  _T_973; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:282:@38057.4]
  wire  _T_974; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:291:@38058.4]
  wire [31:0] x653_rdcol_number; // @[Math.scala 154:22:@38077.4 Math.scala 155:14:@38078.4]
  wire [31:0] _T_989; // @[Math.scala 465:37:@38083.4]
  wire  x654; // @[Math.scala 465:44:@38085.4]
  wire  x655; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 363:59:@38088.4]
  wire  _T_999; // @[FixedPoint.scala 50:25:@38095.4]
  wire [1:0] _T_1003; // @[Bitwise.scala 72:12:@38097.4]
  wire [29:0] _T_1004; // @[FixedPoint.scala 18:52:@38098.4]
  wire  _T_1027; // @[package.scala 96:25:@38132.4 package.scala 96:25:@38133.4]
  wire  _T_1029; // @[implicits.scala 55:10:@38134.4]
  wire  _T_1030; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:194:@38135.4]
  wire  x1098_x656_D1; // @[package.scala 96:25:@38118.4 package.scala 96:25:@38119.4]
  wire  _T_1031; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:282:@38136.4]
  wire  _T_1032; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:291:@38137.4]
  wire [31:0] x665_rdcol_number; // @[Math.scala 154:22:@38156.4 Math.scala 155:14:@38157.4]
  wire [31:0] _T_1047; // @[Math.scala 465:37:@38162.4]
  wire  x666; // @[Math.scala 465:44:@38164.4]
  wire  x667; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 384:59:@38167.4]
  wire  _T_1057; // @[FixedPoint.scala 50:25:@38174.4]
  wire [1:0] _T_1061; // @[Bitwise.scala 72:12:@38176.4]
  wire [29:0] _T_1062; // @[FixedPoint.scala 18:52:@38177.4]
  wire  _T_1085; // @[package.scala 96:25:@38211.4 package.scala 96:25:@38212.4]
  wire  _T_1087; // @[implicits.scala 55:10:@38213.4]
  wire  _T_1088; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 397:194:@38214.4]
  wire  x1099_x668_D1; // @[package.scala 96:25:@38197.4 package.scala 96:25:@38198.4]
  wire  _T_1089; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 397:282:@38215.4]
  wire  _T_1090; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 397:291:@38216.4]
  wire [31:0] x1100_b535_D11_number; // @[package.scala 96:25:@38232.4 package.scala 96:25:@38233.4]
  wire [31:0] _T_1103; // @[Math.scala 406:49:@38239.4]
  wire [31:0] _T_1105; // @[Math.scala 406:56:@38241.4]
  wire [31:0] _T_1106; // @[Math.scala 406:56:@38242.4]
  wire [31:0] x1052_number; // @[implicits.scala 133:21:@38243.4]
  wire  x678; // @[Math.scala 465:44:@38251.4]
  wire  x1101_x678_D1; // @[package.scala 96:25:@38259.4 package.scala 96:25:@38260.4]
  wire  x679; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 409:25:@38263.4]
  wire [31:0] _T_1130; // @[Math.scala 406:49:@38272.4]
  wire [31:0] _T_1132; // @[Math.scala 406:56:@38274.4]
  wire [31:0] _T_1133; // @[Math.scala 406:56:@38275.4]
  wire  _T_1138; // @[FixedPoint.scala 50:25:@38281.4]
  wire [1:0] _T_1142; // @[Bitwise.scala 72:12:@38283.4]
  wire [29:0] _T_1143; // @[FixedPoint.scala 18:52:@38284.4]
  wire  _T_1172; // @[package.scala 96:25:@38336.4 package.scala 96:25:@38337.4]
  wire  _T_1174; // @[implicits.scala 55:10:@38338.4]
  wire  _T_1175; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:194:@38339.4]
  wire  x1103_x680_D1; // @[package.scala 96:25:@38313.4 package.scala 96:25:@38314.4]
  wire  _T_1176; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:282:@38340.4]
  wire  _T_1177; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:291:@38341.4]
  wire  x689; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 438:60:@38352.4]
  wire  _T_1207; // @[package.scala 96:25:@38389.4 package.scala 96:25:@38390.4]
  wire  _T_1209; // @[implicits.scala 55:10:@38391.4]
  wire  _T_1210; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:194:@38392.4]
  wire  x1105_x690_D1; // @[package.scala 96:25:@38375.4 package.scala 96:25:@38376.4]
  wire  _T_1211; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:282:@38393.4]
  wire  _T_1212; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:291:@38394.4]
  wire  x696; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 455:60:@38405.4]
  wire  _T_1240; // @[package.scala 96:25:@38440.4 package.scala 96:25:@38441.4]
  wire  _T_1242; // @[implicits.scala 55:10:@38442.4]
  wire  _T_1243; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:194:@38443.4]
  wire  x1106_x697_D1; // @[package.scala 96:25:@38426.4 package.scala 96:25:@38427.4]
  wire  _T_1244; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:282:@38444.4]
  wire  _T_1245; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:291:@38445.4]
  wire  x703; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 470:59:@38456.4]
  wire  _T_1279; // @[package.scala 96:25:@38509.4 package.scala 96:25:@38510.4]
  wire  _T_1281; // @[implicits.scala 55:10:@38511.4]
  wire  _T_1282; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:194:@38512.4]
  wire  x1108_x704_D2; // @[package.scala 96:25:@38486.4 package.scala 96:25:@38487.4]
  wire  _T_1283; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:282:@38513.4]
  wire  _T_1284; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:291:@38514.4]
  wire  x710; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 489:60:@38525.4]
  wire  _T_1312; // @[package.scala 96:25:@38560.4 package.scala 96:25:@38561.4]
  wire  _T_1314; // @[implicits.scala 55:10:@38562.4]
  wire  _T_1315; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:194:@38563.4]
  wire  x1110_x711_D1; // @[package.scala 96:25:@38546.4 package.scala 96:25:@38547.4]
  wire  _T_1316; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:282:@38564.4]
  wire  _T_1317; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:291:@38565.4]
  wire  x717; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 504:60:@38576.4]
  wire  _T_1345; // @[package.scala 96:25:@38611.4 package.scala 96:25:@38612.4]
  wire  _T_1347; // @[implicits.scala 55:10:@38613.4]
  wire  _T_1348; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:194:@38614.4]
  wire  x1111_x718_D1; // @[package.scala 96:25:@38597.4 package.scala 96:25:@38598.4]
  wire  _T_1349; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:282:@38615.4]
  wire  _T_1350; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:291:@38616.4]
  wire [31:0] x724_rdrow_number; // @[Math.scala 154:22:@38635.4 Math.scala 155:14:@38636.4]
  wire [31:0] _T_1367; // @[Math.scala 406:49:@38642.4]
  wire [31:0] _T_1369; // @[Math.scala 406:56:@38644.4]
  wire [31:0] _T_1370; // @[Math.scala 406:56:@38645.4]
  wire [31:0] x1054_number; // @[implicits.scala 133:21:@38646.4]
  wire  x726; // @[Math.scala 465:44:@38654.4]
  wire  x727; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 525:24:@38657.4]
  wire [31:0] _T_1391; // @[Math.scala 406:49:@38666.4]
  wire [31:0] _T_1393; // @[Math.scala 406:56:@38668.4]
  wire [31:0] _T_1394; // @[Math.scala 406:56:@38669.4]
  wire  _T_1399; // @[FixedPoint.scala 50:25:@38675.4]
  wire [1:0] _T_1403; // @[Bitwise.scala 72:12:@38677.4]
  wire [29:0] _T_1404; // @[FixedPoint.scala 18:52:@38678.4]
  wire  _T_1430; // @[package.scala 96:25:@38721.4 package.scala 96:25:@38722.4]
  wire  _T_1432; // @[implicits.scala 55:10:@38723.4]
  wire  _T_1433; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:194:@38724.4]
  wire  x1113_x728_D1; // @[package.scala 96:25:@38707.4 package.scala 96:25:@38708.4]
  wire  _T_1434; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:282:@38725.4]
  wire  _T_1435; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:291:@38726.4]
  wire  x737; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 546:24:@38737.4]
  wire  _T_1465; // @[package.scala 96:25:@38774.4 package.scala 96:25:@38775.4]
  wire  _T_1467; // @[implicits.scala 55:10:@38776.4]
  wire  _T_1468; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:194:@38777.4]
  wire  x1114_x738_D1; // @[package.scala 96:25:@38760.4 package.scala 96:25:@38761.4]
  wire  _T_1469; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:282:@38778.4]
  wire  _T_1470; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:291:@38779.4]
  wire  x744; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 569:59:@38790.4]
  wire  _T_1498; // @[package.scala 96:25:@38825.4 package.scala 96:25:@38826.4]
  wire  _T_1500; // @[implicits.scala 55:10:@38827.4]
  wire  _T_1501; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:194:@38828.4]
  wire  x1115_x745_D1; // @[package.scala 96:25:@38811.4 package.scala 96:25:@38812.4]
  wire  _T_1502; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:282:@38829.4]
  wire  _T_1503; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:291:@38830.4]
  wire  x751; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 584:59:@38841.4]
  wire  _T_1531; // @[package.scala 96:25:@38876.4 package.scala 96:25:@38877.4]
  wire  _T_1533; // @[implicits.scala 55:10:@38878.4]
  wire  _T_1534; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:194:@38879.4]
  wire  x1116_x752_D1; // @[package.scala 96:25:@38862.4 package.scala 96:25:@38863.4]
  wire  _T_1535; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:282:@38880.4]
  wire  _T_1536; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:291:@38881.4]
  wire  x758; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 599:59:@38892.4]
  wire  _T_1564; // @[package.scala 96:25:@38927.4 package.scala 96:25:@38928.4]
  wire  _T_1566; // @[implicits.scala 55:10:@38929.4]
  wire  _T_1567; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:194:@38930.4]
  wire  x1117_x759_D1; // @[package.scala 96:25:@38913.4 package.scala 96:25:@38914.4]
  wire  _T_1568; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:282:@38931.4]
  wire  _T_1569; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:291:@38932.4]
  wire  x765; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 614:59:@38943.4]
  wire  _T_1597; // @[package.scala 96:25:@38978.4 package.scala 96:25:@38979.4]
  wire  _T_1599; // @[implicits.scala 55:10:@38980.4]
  wire  _T_1600; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:194:@38981.4]
  wire  x1118_x766_D1; // @[package.scala 96:25:@38964.4 package.scala 96:25:@38965.4]
  wire  _T_1601; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:282:@38982.4]
  wire  _T_1602; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:291:@38983.4]
  wire [31:0] x772_rdrow_number; // @[Math.scala 154:22:@39002.4 Math.scala 155:14:@39003.4]
  wire [31:0] _T_1619; // @[Math.scala 406:49:@39009.4]
  wire [31:0] _T_1621; // @[Math.scala 406:56:@39011.4]
  wire [31:0] _T_1622; // @[Math.scala 406:56:@39012.4]
  wire [31:0] x1056_number; // @[implicits.scala 133:21:@39013.4]
  wire  x774; // @[Math.scala 465:44:@39021.4]
  wire  x775; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 635:24:@39024.4]
  wire [31:0] _T_1643; // @[Math.scala 406:49:@39033.4]
  wire [31:0] _T_1645; // @[Math.scala 406:56:@39035.4]
  wire [31:0] _T_1646; // @[Math.scala 406:56:@39036.4]
  wire  _T_1651; // @[FixedPoint.scala 50:25:@39042.4]
  wire [1:0] _T_1655; // @[Bitwise.scala 72:12:@39044.4]
  wire [29:0] _T_1656; // @[FixedPoint.scala 18:52:@39045.4]
  wire  _T_1682; // @[package.scala 96:25:@39088.4 package.scala 96:25:@39089.4]
  wire  _T_1684; // @[implicits.scala 55:10:@39090.4]
  wire  _T_1685; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 652:194:@39091.4]
  wire  x1120_x776_D1; // @[package.scala 96:25:@39074.4 package.scala 96:25:@39075.4]
  wire  _T_1686; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 652:282:@39092.4]
  wire  _T_1687; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 652:291:@39093.4]
  wire  x785; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 656:24:@39104.4]
  wire  _T_1715; // @[package.scala 96:25:@39139.4 package.scala 96:25:@39140.4]
  wire  _T_1717; // @[implicits.scala 55:10:@39141.4]
  wire  _T_1718; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:194:@39142.4]
  wire  x1121_x786_D1; // @[package.scala 96:25:@39125.4 package.scala 96:25:@39126.4]
  wire  _T_1719; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:282:@39143.4]
  wire  _T_1720; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:291:@39144.4]
  wire  x792; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 671:24:@39155.4]
  wire  _T_1750; // @[package.scala 96:25:@39192.4 package.scala 96:25:@39193.4]
  wire  _T_1752; // @[implicits.scala 55:10:@39194.4]
  wire  _T_1753; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:194:@39195.4]
  wire  x1122_x793_D1; // @[package.scala 96:25:@39178.4 package.scala 96:25:@39179.4]
  wire  _T_1754; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:282:@39196.4]
  wire  _T_1755; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:291:@39197.4]
  wire  x799; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 694:59:@39208.4]
  wire  _T_1783; // @[package.scala 96:25:@39243.4 package.scala 96:25:@39244.4]
  wire  _T_1785; // @[implicits.scala 55:10:@39245.4]
  wire  _T_1786; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:194:@39246.4]
  wire  x1123_x800_D1; // @[package.scala 96:25:@39229.4 package.scala 96:25:@39230.4]
  wire  _T_1787; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:282:@39247.4]
  wire  _T_1788; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:291:@39248.4]
  wire  x806; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 709:59:@39259.4]
  wire  _T_1816; // @[package.scala 96:25:@39294.4 package.scala 96:25:@39295.4]
  wire  _T_1818; // @[implicits.scala 55:10:@39296.4]
  wire  _T_1819; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:194:@39297.4]
  wire  x1124_x807_D1; // @[package.scala 96:25:@39280.4 package.scala 96:25:@39281.4]
  wire  _T_1820; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:282:@39298.4]
  wire  _T_1821; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:291:@39299.4]
  wire  x813; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 724:59:@39310.4]
  wire  _T_1849; // @[package.scala 96:25:@39345.4 package.scala 96:25:@39346.4]
  wire  _T_1851; // @[implicits.scala 55:10:@39347.4]
  wire  _T_1852; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 735:194:@39348.4]
  wire  x1125_x814_D1; // @[package.scala 96:25:@39331.4 package.scala 96:25:@39332.4]
  wire  _T_1853; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 735:282:@39349.4]
  wire  _T_1854; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 735:291:@39350.4]
  wire [7:0] x635_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 305:29:@37879.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:445:@37902.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@39362.4]
  wire [8:0] _T_1860; // @[Math.scala 450:32:@39362.4]
  wire [7:0] x687_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 430:29:@38325.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:410:@38348.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@39367.4]
  wire [8:0] _T_1864; // @[Math.scala 450:32:@39367.4]
  wire [7:0] x694_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 447:29:@38378.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:410:@38401.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@39372.4]
  wire [9:0] _T_1868; // @[Math.scala 450:32:@39372.4]
  wire [7:0] x701_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 462:29:@38429.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:410:@38452.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@39377.4]
  wire [8:0] _T_1872; // @[Math.scala 450:32:@39377.4]
  wire [7:0] x742_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 561:29:@38763.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:410:@38786.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@39382.4]
  wire [8:0] _T_1876; // @[Math.scala 450:32:@39382.4]
  wire [7:0] x832_sum_number; // @[Math.scala 154:22:@39471.4 Math.scala 155:14:@39472.4]
  wire [3:0] _T_1912; // @[FixedPoint.scala 18:52:@39477.4]
  wire [7:0] x834_sub_number; // @[Math.scala 195:22:@39504.4 Math.scala 196:14:@39505.4]
  wire  x835; // @[Math.scala 466:37:@39510.4]
  wire [7:0] x833_number; // @[package.scala 96:25:@39484.4 package.scala 96:25:@39485.4]
  wire  x1131_x837_D6; // @[package.scala 96:25:@39577.4 package.scala 96:25:@39578.4]
  wire [7:0] x1130_x833_D6_number; // @[package.scala 96:25:@39568.4 package.scala 96:25:@39569.4]
  wire [7:0] x839_sum_number; // @[Math.scala 154:22:@39559.4 Math.scala 155:14:@39560.4]
  wire [7:0] x840_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 791:24:@39581.4]
  wire [7:0] x643_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 328:29:@37957.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:410:@37980.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@39587.4]
  wire [8:0] _T_1969; // @[Math.scala 450:32:@39587.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@39592.4]
  wire [8:0] _T_1973; // @[Math.scala 450:32:@39592.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@39597.4]
  wire [9:0] _T_1977; // @[Math.scala 450:32:@39597.4]
  wire [7:0] x708_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 481:29:@38498.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:410:@38521.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@39602.4]
  wire [8:0] _T_1981; // @[Math.scala 450:32:@39602.4]
  wire [7:0] x749_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 576:29:@38814.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:410:@38837.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@39607.4]
  wire [8:0] _T_1985; // @[Math.scala 450:32:@39607.4]
  wire [7:0] x853_sum_number; // @[Math.scala 154:22:@39696.4 Math.scala 155:14:@39697.4]
  wire [3:0] _T_2021; // @[FixedPoint.scala 18:52:@39702.4]
  wire [7:0] x855_sub_number; // @[Math.scala 195:22:@39729.4 Math.scala 196:14:@39730.4]
  wire  x856; // @[Math.scala 466:37:@39735.4]
  wire [7:0] x854_number; // @[package.scala 96:25:@39709.4 package.scala 96:25:@39710.4]
  wire  x1137_x858_D6; // @[package.scala 96:25:@39802.4 package.scala 96:25:@39803.4]
  wire [7:0] x1136_x854_D6_number; // @[package.scala 96:25:@39793.4 package.scala 96:25:@39794.4]
  wire [7:0] x860_sum_number; // @[Math.scala 154:22:@39784.4 Math.scala 155:14:@39785.4]
  wire [7:0] x861_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 853:24:@39806.4]
  wire [7:0] x651_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 351:29:@38042.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:410:@38065.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@39810.4]
  wire [8:0] _T_2076; // @[Math.scala 450:32:@39810.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@39815.4]
  wire [9:0] _T_2080; // @[Math.scala 450:32:@39815.4]
  wire [7:0] x715_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 496:29:@38549.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:410:@38572.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@39820.4]
  wire [8:0] _T_2084; // @[Math.scala 450:32:@39820.4]
  wire [7:0] x756_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 591:29:@38865.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:410:@38888.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@39825.4]
  wire [8:0] _T_2088; // @[Math.scala 450:32:@39825.4]
  wire [7:0] x873_sum_number; // @[Math.scala 154:22:@39914.4 Math.scala 155:14:@39915.4]
  wire [3:0] _T_2124; // @[FixedPoint.scala 18:52:@39920.4]
  wire [7:0] x875_sub_number; // @[Math.scala 195:22:@39947.4 Math.scala 196:14:@39948.4]
  wire  x876; // @[Math.scala 466:37:@39953.4]
  wire [7:0] x874_number; // @[package.scala 96:25:@39927.4 package.scala 96:25:@39928.4]
  wire  x1143_x878_D6; // @[package.scala 96:25:@40022.4 package.scala 96:25:@40023.4]
  wire [7:0] x1142_x874_D6_number; // @[package.scala 96:25:@40013.4 package.scala 96:25:@40014.4]
  wire [7:0] x880_sum_number; // @[Math.scala 154:22:@40004.4 Math.scala 155:14:@40005.4]
  wire [7:0] x881_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 913:24:@40026.4]
  wire [7:0] x663_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 372:29:@38121.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:410:@38144.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@40030.4]
  wire [8:0] _T_2181; // @[Math.scala 450:32:@40030.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@40035.4]
  wire [9:0] _T_2185; // @[Math.scala 450:32:@40035.4]
  wire [7:0] x722_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 511:29:@38600.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:410:@38623.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@40040.4]
  wire [8:0] _T_2189; // @[Math.scala 450:32:@40040.4]
  wire [7:0] x763_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 606:29:@38916.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:410:@38939.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@40045.4]
  wire [8:0] _T_2193; // @[Math.scala 450:32:@40045.4]
  wire [7:0] x893_sum_number; // @[Math.scala 154:22:@40134.4 Math.scala 155:14:@40135.4]
  wire [3:0] _T_2229; // @[FixedPoint.scala 18:52:@40140.4]
  wire [7:0] x895_sub_number; // @[Math.scala 195:22:@40167.4 Math.scala 196:14:@40168.4]
  wire  x896; // @[Math.scala 466:37:@40173.4]
  wire [7:0] x894_number; // @[package.scala 96:25:@40147.4 package.scala 96:25:@40148.4]
  wire  x1149_x898_D6; // @[package.scala 96:25:@40240.4 package.scala 96:25:@40241.4]
  wire [7:0] x1148_x894_D6_number; // @[package.scala 96:25:@40231.4 package.scala 96:25:@40232.4]
  wire [7:0] x900_sum_number; // @[Math.scala 154:22:@40222.4 Math.scala 155:14:@40223.4]
  wire [7:0] x901_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 965:24:@40244.4]
  wire [7:0] x735_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 538:29:@38710.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:410:@38733.4]
  wire [8:0] _GEN_18; // @[Math.scala 450:32:@40248.4]
  wire [8:0] _T_2284; // @[Math.scala 450:32:@40248.4]
  wire [9:0] _GEN_19; // @[Math.scala 450:32:@40253.4]
  wire [9:0] _T_2288; // @[Math.scala 450:32:@40253.4]
  wire [7:0] x790_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 663:29:@39128.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:410:@39151.4]
  wire [8:0] _GEN_20; // @[Math.scala 450:32:@40258.4]
  wire [8:0] _T_2292; // @[Math.scala 450:32:@40258.4]
  wire [7:0] x912_sum_number; // @[Math.scala 154:22:@40347.4 Math.scala 155:14:@40348.4]
  wire [3:0] _T_2328; // @[FixedPoint.scala 18:52:@40353.4]
  wire [7:0] x914_sub_number; // @[Math.scala 195:22:@40380.4 Math.scala 196:14:@40381.4]
  wire  x915; // @[Math.scala 466:37:@40386.4]
  wire [7:0] x913_number; // @[package.scala 96:25:@40360.4 package.scala 96:25:@40361.4]
  wire  x1154_x917_D6; // @[package.scala 96:25:@40446.4 package.scala 96:25:@40447.4]
  wire [7:0] x1155_x913_D6_number; // @[package.scala 96:25:@40455.4 package.scala 96:25:@40456.4]
  wire [7:0] x919_sum_number; // @[Math.scala 154:22:@40437.4 Math.scala 155:14:@40438.4]
  wire [7:0] x920_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1023:24:@40459.4]
  wire [9:0] _GEN_21; // @[Math.scala 450:32:@40463.4]
  wire [9:0] _T_2385; // @[Math.scala 450:32:@40463.4]
  wire [7:0] x797_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 686:29:@39181.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:410:@39204.4]
  wire [8:0] _GEN_22; // @[Math.scala 450:32:@40468.4]
  wire [8:0] _T_2389; // @[Math.scala 450:32:@40468.4]
  wire [7:0] x930_sum_number; // @[Math.scala 154:22:@40557.4 Math.scala 155:14:@40558.4]
  wire [3:0] _T_2425; // @[FixedPoint.scala 18:52:@40563.4]
  wire [7:0] x932_sub_number; // @[Math.scala 195:22:@40590.4 Math.scala 196:14:@40591.4]
  wire  x933; // @[Math.scala 466:37:@40596.4]
  wire [7:0] x931_number; // @[package.scala 96:25:@40570.4 package.scala 96:25:@40571.4]
  wire  x1160_x935_D6; // @[package.scala 96:25:@40654.4 package.scala 96:25:@40655.4]
  wire [7:0] x1161_x931_D6_number; // @[package.scala 96:25:@40663.4 package.scala 96:25:@40664.4]
  wire [7:0] x937_sum_number; // @[Math.scala 154:22:@40645.4 Math.scala 155:14:@40646.4]
  wire [7:0] x938_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1071:24:@40667.4]
  wire [9:0] _GEN_23; // @[Math.scala 450:32:@40671.4]
  wire [9:0] _T_2480; // @[Math.scala 450:32:@40671.4]
  wire [7:0] x804_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 701:29:@39232.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:410:@39255.4]
  wire [8:0] _GEN_24; // @[Math.scala 450:32:@40676.4]
  wire [8:0] _T_2484; // @[Math.scala 450:32:@40676.4]
  wire [7:0] x948_sum_number; // @[Math.scala 154:22:@40765.4 Math.scala 155:14:@40766.4]
  wire [3:0] _T_2520; // @[FixedPoint.scala 18:52:@40771.4]
  wire [7:0] x950_sub_number; // @[Math.scala 195:22:@40798.4 Math.scala 196:14:@40799.4]
  wire  x951; // @[Math.scala 466:37:@40804.4]
  wire [7:0] x949_number; // @[package.scala 96:25:@40778.4 package.scala 96:25:@40779.4]
  wire  x1166_x953_D6; // @[package.scala 96:25:@40864.4 package.scala 96:25:@40865.4]
  wire [7:0] x1167_x949_D6_number; // @[package.scala 96:25:@40873.4 package.scala 96:25:@40874.4]
  wire [7:0] x955_sum_number; // @[Math.scala 154:22:@40855.4 Math.scala 155:14:@40856.4]
  wire [7:0] x956_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1127:24:@40877.4]
  wire [9:0] _GEN_25; // @[Math.scala 450:32:@40881.4]
  wire [9:0] _T_2577; // @[Math.scala 450:32:@40881.4]
  wire [7:0] x770_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 621:29:@38967.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:410:@38990.4]
  wire [8:0] _GEN_26; // @[Math.scala 450:32:@40886.4]
  wire [8:0] _T_2581; // @[Math.scala 450:32:@40886.4]
  wire [7:0] x811_rd_0_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 716:29:@39283.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:410:@39306.4]
  wire [8:0] _GEN_27; // @[Math.scala 450:32:@40891.4]
  wire [8:0] _T_2585; // @[Math.scala 450:32:@40891.4]
  wire [7:0] x967_sum_number; // @[Math.scala 154:22:@40980.4 Math.scala 155:14:@40981.4]
  wire [3:0] _T_2621; // @[FixedPoint.scala 18:52:@40986.4]
  wire [7:0] x969_sub_number; // @[Math.scala 195:22:@41013.4 Math.scala 196:14:@41014.4]
  wire  x970; // @[Math.scala 466:37:@41019.4]
  wire [7:0] x968_number; // @[package.scala 96:25:@40993.4 package.scala 96:25:@40994.4]
  wire  x1172_x972_D6; // @[package.scala 96:25:@41077.4 package.scala 96:25:@41078.4]
  wire [7:0] x1173_x968_D6_number; // @[package.scala 96:25:@41086.4 package.scala 96:25:@41087.4]
  wire [7:0] x974_sum_number; // @[Math.scala 154:22:@41068.4 Math.scala 155:14:@41069.4]
  wire [7:0] x975_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1177:24:@41090.4]
  wire [31:0] _T_2690; // @[Cat.scala 30:58:@41104.4]
  wire [31:0] _T_2693; // @[Cat.scala 30:58:@41107.4]
  wire  _T_2706; // @[package.scala 96:25:@41143.4 package.scala 96:25:@41144.4]
  wire  _T_2708; // @[implicits.scala 55:10:@41145.4]
  wire  x1174_b537_D26; // @[package.scala 96:25:@41125.4 package.scala 96:25:@41126.4]
  wire  _T_2709; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1187:116:@41146.4]
  wire  x1175_b538_D26; // @[package.scala 96:25:@41134.4 package.scala 96:25:@41135.4]
  wire  _T_2710; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1187:123:@41147.4]
  wire [31:0] x1061_x1048_D8_number; // @[package.scala 96:25:@37077.4 package.scala 96:25:@37078.4]
  wire [31:0] x1063_x553_sum_D7_number; // @[package.scala 96:25:@37095.4 package.scala 96:25:@37096.4]
  wire [31:0] x1065_x563_sum_D6_number; // @[package.scala 96:25:@37171.4 package.scala 96:25:@37172.4]
  wire [31:0] x1068_x572_sum_D6_number; // @[package.scala 96:25:@37256.4 package.scala 96:25:@37257.4]
  wire [31:0] x1070_x581_sum_D6_number; // @[package.scala 96:25:@37332.4 package.scala 96:25:@37333.4]
  wire [31:0] x1072_x1049_D7_number; // @[package.scala 96:25:@37468.4 package.scala 96:25:@37469.4]
  wire [31:0] x1073_x595_sum_D6_number; // @[package.scala 96:25:@37477.4 package.scala 96:25:@37478.4]
  wire [31:0] x1075_x601_sum_D6_number; // @[package.scala 96:25:@37532.4 package.scala 96:25:@37533.4]
  wire [31:0] x1077_x606_sum_D6_number; // @[package.scala 96:25:@37587.4 package.scala 96:25:@37588.4]
  wire [31:0] x1080_x611_sum_D6_number; // @[package.scala 96:25:@37651.4 package.scala 96:25:@37652.4]
  wire [31:0] x623_sum_number; // @[Math.scala 154:22:@37764.4 Math.scala 155:14:@37765.4]
  wire [31:0] x1085_x1051_D1_number; // @[package.scala 96:25:@37782.4 package.scala 96:25:@37783.4]
  wire [31:0] x632_sum_number; // @[Math.scala 154:22:@37867.4 Math.scala 155:14:@37868.4]
  wire [31:0] x640_sum_number; // @[Math.scala 154:22:@37945.4 Math.scala 155:14:@37946.4]
  wire [31:0] x648_sum_number; // @[Math.scala 154:22:@38030.4 Math.scala 155:14:@38031.4]
  wire [31:0] x659_sum_number; // @[Math.scala 154:22:@38109.4 Math.scala 155:14:@38110.4]
  wire [31:0] x671_sum_number; // @[Math.scala 154:22:@38188.4 Math.scala 155:14:@38189.4]
  wire [31:0] x683_sum_number; // @[Math.scala 154:22:@38304.4 Math.scala 155:14:@38305.4]
  wire [31:0] x1104_x1053_D2_number; // @[package.scala 96:25:@38322.4 package.scala 96:25:@38323.4]
  wire [31:0] x691_sum_number; // @[Math.scala 154:22:@38366.4 Math.scala 155:14:@38367.4]
  wire [31:0] x698_sum_number; // @[Math.scala 154:22:@38417.4 Math.scala 155:14:@38418.4]
  wire [31:0] x1109_x705_sum_D1_number; // @[package.scala 96:25:@38495.4 package.scala 96:25:@38496.4]
  wire [31:0] x712_sum_number; // @[Math.scala 154:22:@38537.4 Math.scala 155:14:@38538.4]
  wire [31:0] x719_sum_number; // @[Math.scala 154:22:@38588.4 Math.scala 155:14:@38589.4]
  wire [31:0] x731_sum_number; // @[Math.scala 154:22:@38689.4 Math.scala 155:14:@38690.4]
  wire [31:0] x1112_x1055_D1_number; // @[package.scala 96:25:@38698.4 package.scala 96:25:@38699.4]
  wire [31:0] x739_sum_number; // @[Math.scala 154:22:@38751.4 Math.scala 155:14:@38752.4]
  wire [31:0] x746_sum_number; // @[Math.scala 154:22:@38802.4 Math.scala 155:14:@38803.4]
  wire [31:0] x753_sum_number; // @[Math.scala 154:22:@38853.4 Math.scala 155:14:@38854.4]
  wire [31:0] x760_sum_number; // @[Math.scala 154:22:@38904.4 Math.scala 155:14:@38905.4]
  wire [31:0] x767_sum_number; // @[Math.scala 154:22:@38955.4 Math.scala 155:14:@38956.4]
  wire [31:0] x779_sum_number; // @[Math.scala 154:22:@39056.4 Math.scala 155:14:@39057.4]
  wire [31:0] x1119_x1057_D1_number; // @[package.scala 96:25:@39065.4 package.scala 96:25:@39066.4]
  wire [31:0] x787_sum_number; // @[Math.scala 154:22:@39116.4 Math.scala 155:14:@39117.4]
  wire [31:0] x794_sum_number; // @[Math.scala 154:22:@39169.4 Math.scala 155:14:@39170.4]
  wire [31:0] x801_sum_number; // @[Math.scala 154:22:@39220.4 Math.scala 155:14:@39221.4]
  wire [31:0] x808_sum_number; // @[Math.scala 154:22:@39271.4 Math.scala 155:14:@39272.4]
  wire [31:0] x815_sum_number; // @[Math.scala 154:22:@39322.4 Math.scala 155:14:@39323.4]
  _ _ ( // @[Math.scala 709:24:@36688.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@36700.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x539_lb_0 x539_lb_0 ( // @[m_x539_lb_0.scala 57:17:@36710.4]
    .clock(x539_lb_0_clock),
    .reset(x539_lb_0_reset),
    .io_rPort_23_banks_0(x539_lb_0_io_rPort_23_banks_0),
    .io_rPort_23_ofs_0(x539_lb_0_io_rPort_23_ofs_0),
    .io_rPort_23_en_0(x539_lb_0_io_rPort_23_en_0),
    .io_rPort_23_backpressure(x539_lb_0_io_rPort_23_backpressure),
    .io_rPort_23_output_0(x539_lb_0_io_rPort_23_output_0),
    .io_rPort_22_banks_0(x539_lb_0_io_rPort_22_banks_0),
    .io_rPort_22_ofs_0(x539_lb_0_io_rPort_22_ofs_0),
    .io_rPort_22_en_0(x539_lb_0_io_rPort_22_en_0),
    .io_rPort_22_backpressure(x539_lb_0_io_rPort_22_backpressure),
    .io_rPort_22_output_0(x539_lb_0_io_rPort_22_output_0),
    .io_rPort_21_banks_0(x539_lb_0_io_rPort_21_banks_0),
    .io_rPort_21_ofs_0(x539_lb_0_io_rPort_21_ofs_0),
    .io_rPort_21_en_0(x539_lb_0_io_rPort_21_en_0),
    .io_rPort_21_backpressure(x539_lb_0_io_rPort_21_backpressure),
    .io_rPort_21_output_0(x539_lb_0_io_rPort_21_output_0),
    .io_rPort_20_banks_0(x539_lb_0_io_rPort_20_banks_0),
    .io_rPort_20_ofs_0(x539_lb_0_io_rPort_20_ofs_0),
    .io_rPort_20_en_0(x539_lb_0_io_rPort_20_en_0),
    .io_rPort_20_backpressure(x539_lb_0_io_rPort_20_backpressure),
    .io_rPort_20_output_0(x539_lb_0_io_rPort_20_output_0),
    .io_rPort_19_banks_0(x539_lb_0_io_rPort_19_banks_0),
    .io_rPort_19_ofs_0(x539_lb_0_io_rPort_19_ofs_0),
    .io_rPort_19_en_0(x539_lb_0_io_rPort_19_en_0),
    .io_rPort_19_backpressure(x539_lb_0_io_rPort_19_backpressure),
    .io_rPort_19_output_0(x539_lb_0_io_rPort_19_output_0),
    .io_rPort_18_banks_0(x539_lb_0_io_rPort_18_banks_0),
    .io_rPort_18_ofs_0(x539_lb_0_io_rPort_18_ofs_0),
    .io_rPort_18_en_0(x539_lb_0_io_rPort_18_en_0),
    .io_rPort_18_backpressure(x539_lb_0_io_rPort_18_backpressure),
    .io_rPort_18_output_0(x539_lb_0_io_rPort_18_output_0),
    .io_rPort_17_banks_0(x539_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x539_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x539_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x539_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x539_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_0(x539_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x539_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x539_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x539_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x539_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_0(x539_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x539_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x539_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x539_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x539_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_0(x539_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x539_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x539_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x539_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x539_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_0(x539_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x539_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x539_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x539_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x539_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_0(x539_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x539_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x539_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x539_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x539_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_0(x539_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x539_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x539_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x539_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x539_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_0(x539_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x539_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x539_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x539_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x539_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_0(x539_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x539_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x539_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x539_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x539_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x539_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x539_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x539_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x539_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x539_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x539_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x539_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x539_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x539_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x539_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x539_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x539_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x539_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x539_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x539_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x539_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x539_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x539_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x539_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x539_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x539_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x539_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x539_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x539_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x539_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x539_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x539_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x539_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x539_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x539_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x539_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x539_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x539_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x539_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x539_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x539_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x539_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x539_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x539_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x539_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x539_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x539_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x539_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x539_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x539_lb_0_io_rPort_0_output_0),
    .io_wPort_7_banks_0(x539_lb_0_io_wPort_7_banks_0),
    .io_wPort_7_ofs_0(x539_lb_0_io_wPort_7_ofs_0),
    .io_wPort_7_data_0(x539_lb_0_io_wPort_7_data_0),
    .io_wPort_7_en_0(x539_lb_0_io_wPort_7_en_0),
    .io_wPort_6_banks_0(x539_lb_0_io_wPort_6_banks_0),
    .io_wPort_6_ofs_0(x539_lb_0_io_wPort_6_ofs_0),
    .io_wPort_6_data_0(x539_lb_0_io_wPort_6_data_0),
    .io_wPort_6_en_0(x539_lb_0_io_wPort_6_en_0),
    .io_wPort_5_banks_0(x539_lb_0_io_wPort_5_banks_0),
    .io_wPort_5_ofs_0(x539_lb_0_io_wPort_5_ofs_0),
    .io_wPort_5_data_0(x539_lb_0_io_wPort_5_data_0),
    .io_wPort_5_en_0(x539_lb_0_io_wPort_5_en_0),
    .io_wPort_4_banks_0(x539_lb_0_io_wPort_4_banks_0),
    .io_wPort_4_ofs_0(x539_lb_0_io_wPort_4_ofs_0),
    .io_wPort_4_data_0(x539_lb_0_io_wPort_4_data_0),
    .io_wPort_4_en_0(x539_lb_0_io_wPort_4_en_0),
    .io_wPort_3_banks_0(x539_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x539_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x539_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x539_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x539_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x539_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x539_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x539_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x539_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x539_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x539_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x539_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x539_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x539_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x539_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x539_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_148 RetimeWrapper ( // @[package.scala 93:22:@36936.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x553_sum x553_sum_1 ( // @[Math.scala 150:24:@37044.4]
    .clock(x553_sum_1_clock),
    .reset(x553_sum_1_reset),
    .io_a(x553_sum_1_io_a),
    .io_b(x553_sum_1_io_b),
    .io_flow(x553_sum_1_io_flow),
    .io_result(x553_sum_1_io_result)
  );
  RetimeWrapper_150 RetimeWrapper_1 ( // @[package.scala 93:22:@37054.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_2 ( // @[package.scala 93:22:@37063.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_152 RetimeWrapper_3 ( // @[package.scala 93:22:@37072.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_4 ( // @[package.scala 93:22:@37081.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_154 RetimeWrapper_5 ( // @[package.scala 93:22:@37090.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_6 ( // @[package.scala 93:22:@37103.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x553_sum x559_rdcol_1 ( // @[Math.scala 150:24:@37126.4]
    .clock(x559_rdcol_1_clock),
    .reset(x559_rdcol_1_reset),
    .io_a(x559_rdcol_1_io_a),
    .io_b(x559_rdcol_1_io_b),
    .io_flow(x559_rdcol_1_io_flow),
    .io_result(x559_rdcol_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_7 ( // @[package.scala 93:22:@37147.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x553_sum x563_sum_1 ( // @[Math.scala 150:24:@37156.4]
    .clock(x563_sum_1_clock),
    .reset(x563_sum_1_reset),
    .io_a(x563_sum_1_io_a),
    .io_b(x563_sum_1_io_b),
    .io_flow(x563_sum_1_io_flow),
    .io_result(x563_sum_1_io_result)
  );
  RetimeWrapper_159 RetimeWrapper_8 ( // @[package.scala 93:22:@37166.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_9 ( // @[package.scala 93:22:@37175.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_10 ( // @[package.scala 93:22:@37188.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x553_sum x568_rdcol_1 ( // @[Math.scala 150:24:@37211.4]
    .clock(x568_rdcol_1_clock),
    .reset(x568_rdcol_1_reset),
    .io_a(x568_rdcol_1_io_a),
    .io_b(x568_rdcol_1_io_b),
    .io_flow(x568_rdcol_1_io_flow),
    .io_result(x568_rdcol_1_io_result)
  );
  x553_sum x572_sum_1 ( // @[Math.scala 150:24:@37232.4]
    .clock(x572_sum_1_clock),
    .reset(x572_sum_1_reset),
    .io_a(x572_sum_1_io_a),
    .io_b(x572_sum_1_io_b),
    .io_flow(x572_sum_1_io_flow),
    .io_result(x572_sum_1_io_result)
  );
  RetimeWrapper_153 RetimeWrapper_11 ( // @[package.scala 93:22:@37242.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_12 ( // @[package.scala 93:22:@37251.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_13 ( // @[package.scala 93:22:@37264.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x553_sum x577_rdcol_1 ( // @[Math.scala 150:24:@37287.4]
    .clock(x577_rdcol_1_clock),
    .reset(x577_rdcol_1_reset),
    .io_a(x577_rdcol_1_io_a),
    .io_b(x577_rdcol_1_io_b),
    .io_flow(x577_rdcol_1_io_flow),
    .io_result(x577_rdcol_1_io_result)
  );
  x553_sum x581_sum_1 ( // @[Math.scala 150:24:@37308.4]
    .clock(x581_sum_1_clock),
    .reset(x581_sum_1_reset),
    .io_a(x581_sum_1_io_a),
    .io_b(x581_sum_1_io_b),
    .io_flow(x581_sum_1_io_flow),
    .io_result(x581_sum_1_io_result)
  );
  RetimeWrapper_153 RetimeWrapper_14 ( // @[package.scala 93:22:@37318.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_15 ( // @[package.scala 93:22:@37327.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_16 ( // @[package.scala 93:22:@37340.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  x553_sum x586_rdrow_1 ( // @[Math.scala 150:24:@37363.4]
    .clock(x586_rdrow_1_clock),
    .reset(x586_rdrow_1_reset),
    .io_a(x586_rdrow_1_io_a),
    .io_b(x586_rdrow_1_io_b),
    .io_flow(x586_rdrow_1_io_flow),
    .io_result(x586_rdrow_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_17 ( // @[package.scala 93:22:@37444.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x553_sum x595_sum_1 ( // @[Math.scala 150:24:@37453.4]
    .clock(x595_sum_1_clock),
    .reset(x595_sum_1_reset),
    .io_a(x595_sum_1_io_a),
    .io_b(x595_sum_1_io_b),
    .io_flow(x595_sum_1_io_flow),
    .io_result(x595_sum_1_io_result)
  );
  RetimeWrapper_154 RetimeWrapper_18 ( // @[package.scala 93:22:@37463.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_19 ( // @[package.scala 93:22:@37472.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_20 ( // @[package.scala 93:22:@37481.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_21 ( // @[package.scala 93:22:@37494.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  x553_sum x601_sum_1 ( // @[Math.scala 150:24:@37517.4]
    .clock(x601_sum_1_clock),
    .reset(x601_sum_1_reset),
    .io_a(x601_sum_1_io_a),
    .io_b(x601_sum_1_io_b),
    .io_flow(x601_sum_1_io_flow),
    .io_result(x601_sum_1_io_result)
  );
  RetimeWrapper_159 RetimeWrapper_22 ( // @[package.scala 93:22:@37527.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_23 ( // @[package.scala 93:22:@37536.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_24 ( // @[package.scala 93:22:@37549.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  x553_sum x606_sum_1 ( // @[Math.scala 150:24:@37572.4]
    .clock(x606_sum_1_clock),
    .reset(x606_sum_1_reset),
    .io_a(x606_sum_1_io_a),
    .io_b(x606_sum_1_io_b),
    .io_flow(x606_sum_1_io_flow),
    .io_result(x606_sum_1_io_result)
  );
  RetimeWrapper_159 RetimeWrapper_25 ( // @[package.scala 93:22:@37582.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_153 RetimeWrapper_26 ( // @[package.scala 93:22:@37591.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_27 ( // @[package.scala 93:22:@37604.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x553_sum x611_sum_1 ( // @[Math.scala 150:24:@37627.4]
    .clock(x611_sum_1_clock),
    .reset(x611_sum_1_reset),
    .io_a(x611_sum_1_io_a),
    .io_b(x611_sum_1_io_b),
    .io_flow(x611_sum_1_io_flow),
    .io_result(x611_sum_1_io_result)
  );
  RetimeWrapper_153 RetimeWrapper_28 ( // @[package.scala 93:22:@37637.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_159 RetimeWrapper_29 ( // @[package.scala 93:22:@37646.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_150 RetimeWrapper_30 ( // @[package.scala 93:22:@37659.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_31 ( // @[package.scala 93:22:@37680.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_32 ( // @[package.scala 93:22:@37707.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_33 ( // @[package.scala 93:22:@37749.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  x553_sum x623_sum_1 ( // @[Math.scala 150:24:@37758.4]
    .clock(x623_sum_1_clock),
    .reset(x623_sum_1_reset),
    .io_a(x623_sum_1_io_a),
    .io_b(x623_sum_1_io_b),
    .io_flow(x623_sum_1_io_flow),
    .io_result(x623_sum_1_io_result)
  );
  RetimeWrapper_195 RetimeWrapper_34 ( // @[package.scala 93:22:@37768.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_35 ( // @[package.scala 93:22:@37777.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_36 ( // @[package.scala 93:22:@37786.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper RetimeWrapper_37 ( // @[package.scala 93:22:@37795.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_38 ( // @[package.scala 93:22:@37809.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_39 ( // @[package.scala 93:22:@37830.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_40 ( // @[package.scala 93:22:@37852.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x553_sum x632_sum_1 ( // @[Math.scala 150:24:@37861.4]
    .clock(x632_sum_1_clock),
    .reset(x632_sum_1_reset),
    .io_a(x632_sum_1_io_a),
    .io_b(x632_sum_1_io_b),
    .io_flow(x632_sum_1_io_flow),
    .io_result(x632_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@37871.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_42 ( // @[package.scala 93:22:@37885.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_43 ( // @[package.scala 93:22:@37906.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_44 ( // @[package.scala 93:22:@37930.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  x553_sum x640_sum_1 ( // @[Math.scala 150:24:@37939.4]
    .clock(x640_sum_1_clock),
    .reset(x640_sum_1_reset),
    .io_a(x640_sum_1_io_a),
    .io_b(x640_sum_1_io_b),
    .io_flow(x640_sum_1_io_flow),
    .io_result(x640_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@37949.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_46 ( // @[package.scala 93:22:@37963.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_47 ( // @[package.scala 93:22:@37984.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper RetimeWrapper_48 ( // @[package.scala 93:22:@38000.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_212 RetimeWrapper_49 ( // @[package.scala 93:22:@38015.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x553_sum x648_sum_1 ( // @[Math.scala 150:24:@38024.4]
    .clock(x648_sum_1_clock),
    .reset(x648_sum_1_reset),
    .io_a(x648_sum_1_io_a),
    .io_b(x648_sum_1_io_b),
    .io_flow(x648_sum_1_io_flow),
    .io_result(x648_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_50 ( // @[package.scala 93:22:@38034.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_51 ( // @[package.scala 93:22:@38048.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x553_sum x653_rdcol_1 ( // @[Math.scala 150:24:@38071.4]
    .clock(x653_rdcol_1_clock),
    .reset(x653_rdcol_1_reset),
    .io_a(x653_rdcol_1_io_a),
    .io_b(x653_rdcol_1_io_b),
    .io_flow(x653_rdcol_1_io_flow),
    .io_result(x653_rdcol_1_io_result)
  );
  x553_sum x659_sum_1 ( // @[Math.scala 150:24:@38103.4]
    .clock(x659_sum_1_clock),
    .reset(x659_sum_1_reset),
    .io_a(x659_sum_1_io_a),
    .io_b(x659_sum_1_io_b),
    .io_flow(x659_sum_1_io_flow),
    .io_result(x659_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_52 ( // @[package.scala 93:22:@38113.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_53 ( // @[package.scala 93:22:@38127.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x553_sum x665_rdcol_1 ( // @[Math.scala 150:24:@38150.4]
    .clock(x665_rdcol_1_clock),
    .reset(x665_rdcol_1_reset),
    .io_a(x665_rdcol_1_io_a),
    .io_b(x665_rdcol_1_io_b),
    .io_flow(x665_rdcol_1_io_flow),
    .io_result(x665_rdcol_1_io_result)
  );
  x553_sum x671_sum_1 ( // @[Math.scala 150:24:@38182.4]
    .clock(x671_sum_1_clock),
    .reset(x671_sum_1_reset),
    .io_a(x671_sum_1_io_a),
    .io_b(x671_sum_1_io_b),
    .io_flow(x671_sum_1_io_flow),
    .io_result(x671_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_54 ( // @[package.scala 93:22:@38192.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_55 ( // @[package.scala 93:22:@38206.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_56 ( // @[package.scala 93:22:@38227.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@38254.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_58 ( // @[package.scala 93:22:@38289.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x553_sum x683_sum_1 ( // @[Math.scala 150:24:@38298.4]
    .clock(x683_sum_1_clock),
    .reset(x683_sum_1_reset),
    .io_a(x683_sum_1_io_a),
    .io_b(x683_sum_1_io_b),
    .io_flow(x683_sum_1_io_flow),
    .io_result(x683_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@38308.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_229 RetimeWrapper_60 ( // @[package.scala 93:22:@38317.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_61 ( // @[package.scala 93:22:@38331.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x553_sum x691_sum_1 ( // @[Math.scala 150:24:@38360.4]
    .clock(x691_sum_1_clock),
    .reset(x691_sum_1_reset),
    .io_a(x691_sum_1_io_a),
    .io_b(x691_sum_1_io_b),
    .io_flow(x691_sum_1_io_flow),
    .io_result(x691_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@38370.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_63 ( // @[package.scala 93:22:@38384.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x553_sum x698_sum_1 ( // @[Math.scala 150:24:@38411.4]
    .clock(x698_sum_1_clock),
    .reset(x698_sum_1_reset),
    .io_a(x698_sum_1_io_a),
    .io_b(x698_sum_1_io_b),
    .io_flow(x698_sum_1_io_flow),
    .io_result(x698_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_64 ( // @[package.scala 93:22:@38421.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_65 ( // @[package.scala 93:22:@38435.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_66 ( // @[package.scala 93:22:@38462.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x553_sum x705_sum_1 ( // @[Math.scala 150:24:@38471.4]
    .clock(x705_sum_1_clock),
    .reset(x705_sum_1_reset),
    .io_a(x705_sum_1_io_a),
    .io_b(x705_sum_1_io_b),
    .io_flow(x705_sum_1_io_flow),
    .io_result(x705_sum_1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@38481.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_149 RetimeWrapper_68 ( // @[package.scala 93:22:@38490.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_69 ( // @[package.scala 93:22:@38504.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x553_sum x712_sum_1 ( // @[Math.scala 150:24:@38531.4]
    .clock(x712_sum_1_clock),
    .reset(x712_sum_1_reset),
    .io_a(x712_sum_1_io_a),
    .io_b(x712_sum_1_io_b),
    .io_flow(x712_sum_1_io_flow),
    .io_result(x712_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_70 ( // @[package.scala 93:22:@38541.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_71 ( // @[package.scala 93:22:@38555.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x553_sum x719_sum_1 ( // @[Math.scala 150:24:@38582.4]
    .clock(x719_sum_1_clock),
    .reset(x719_sum_1_reset),
    .io_a(x719_sum_1_io_a),
    .io_b(x719_sum_1_io_b),
    .io_flow(x719_sum_1_io_flow),
    .io_result(x719_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_72 ( // @[package.scala 93:22:@38592.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_73 ( // @[package.scala 93:22:@38606.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x553_sum x724_rdrow_1 ( // @[Math.scala 150:24:@38629.4]
    .clock(x724_rdrow_1_clock),
    .reset(x724_rdrow_1_reset),
    .io_a(x724_rdrow_1_io_a),
    .io_b(x724_rdrow_1_io_b),
    .io_flow(x724_rdrow_1_io_flow),
    .io_result(x724_rdrow_1_io_result)
  );
  x553_sum x731_sum_1 ( // @[Math.scala 150:24:@38683.4]
    .clock(x731_sum_1_clock),
    .reset(x731_sum_1_reset),
    .io_a(x731_sum_1_io_a),
    .io_b(x731_sum_1_io_b),
    .io_flow(x731_sum_1_io_flow),
    .io_result(x731_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_74 ( // @[package.scala 93:22:@38693.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper RetimeWrapper_75 ( // @[package.scala 93:22:@38702.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_76 ( // @[package.scala 93:22:@38716.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x553_sum x739_sum_1 ( // @[Math.scala 150:24:@38745.4]
    .clock(x739_sum_1_clock),
    .reset(x739_sum_1_reset),
    .io_a(x739_sum_1_io_a),
    .io_b(x739_sum_1_io_b),
    .io_flow(x739_sum_1_io_flow),
    .io_result(x739_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_77 ( // @[package.scala 93:22:@38755.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_78 ( // @[package.scala 93:22:@38769.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x553_sum x746_sum_1 ( // @[Math.scala 150:24:@38796.4]
    .clock(x746_sum_1_clock),
    .reset(x746_sum_1_reset),
    .io_a(x746_sum_1_io_a),
    .io_b(x746_sum_1_io_b),
    .io_flow(x746_sum_1_io_flow),
    .io_result(x746_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_79 ( // @[package.scala 93:22:@38806.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_80 ( // @[package.scala 93:22:@38820.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x553_sum x753_sum_1 ( // @[Math.scala 150:24:@38847.4]
    .clock(x753_sum_1_clock),
    .reset(x753_sum_1_reset),
    .io_a(x753_sum_1_io_a),
    .io_b(x753_sum_1_io_b),
    .io_flow(x753_sum_1_io_flow),
    .io_result(x753_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_81 ( // @[package.scala 93:22:@38857.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_82 ( // @[package.scala 93:22:@38871.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x553_sum x760_sum_1 ( // @[Math.scala 150:24:@38898.4]
    .clock(x760_sum_1_clock),
    .reset(x760_sum_1_reset),
    .io_a(x760_sum_1_io_a),
    .io_b(x760_sum_1_io_b),
    .io_flow(x760_sum_1_io_flow),
    .io_result(x760_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_83 ( // @[package.scala 93:22:@38908.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_84 ( // @[package.scala 93:22:@38922.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x553_sum x767_sum_1 ( // @[Math.scala 150:24:@38949.4]
    .clock(x767_sum_1_clock),
    .reset(x767_sum_1_reset),
    .io_a(x767_sum_1_io_a),
    .io_b(x767_sum_1_io_b),
    .io_flow(x767_sum_1_io_flow),
    .io_result(x767_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@38959.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_86 ( // @[package.scala 93:22:@38973.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  x553_sum x772_rdrow_1 ( // @[Math.scala 150:24:@38996.4]
    .clock(x772_rdrow_1_clock),
    .reset(x772_rdrow_1_reset),
    .io_a(x772_rdrow_1_io_a),
    .io_b(x772_rdrow_1_io_b),
    .io_flow(x772_rdrow_1_io_flow),
    .io_result(x772_rdrow_1_io_result)
  );
  x553_sum x779_sum_1 ( // @[Math.scala 150:24:@39050.4]
    .clock(x779_sum_1_clock),
    .reset(x779_sum_1_reset),
    .io_a(x779_sum_1_io_a),
    .io_b(x779_sum_1_io_b),
    .io_flow(x779_sum_1_io_flow),
    .io_result(x779_sum_1_io_result)
  );
  RetimeWrapper_149 RetimeWrapper_87 ( // @[package.scala 93:22:@39060.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper RetimeWrapper_88 ( // @[package.scala 93:22:@39069.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_89 ( // @[package.scala 93:22:@39083.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  x553_sum x787_sum_1 ( // @[Math.scala 150:24:@39110.4]
    .clock(x787_sum_1_clock),
    .reset(x787_sum_1_reset),
    .io_a(x787_sum_1_io_a),
    .io_b(x787_sum_1_io_b),
    .io_flow(x787_sum_1_io_flow),
    .io_result(x787_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_90 ( // @[package.scala 93:22:@39120.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_91 ( // @[package.scala 93:22:@39134.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x553_sum x794_sum_1 ( // @[Math.scala 150:24:@39163.4]
    .clock(x794_sum_1_clock),
    .reset(x794_sum_1_reset),
    .io_a(x794_sum_1_io_a),
    .io_b(x794_sum_1_io_b),
    .io_flow(x794_sum_1_io_flow),
    .io_result(x794_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_92 ( // @[package.scala 93:22:@39173.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_93 ( // @[package.scala 93:22:@39187.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  x553_sum x801_sum_1 ( // @[Math.scala 150:24:@39214.4]
    .clock(x801_sum_1_clock),
    .reset(x801_sum_1_reset),
    .io_a(x801_sum_1_io_a),
    .io_b(x801_sum_1_io_b),
    .io_flow(x801_sum_1_io_flow),
    .io_result(x801_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_94 ( // @[package.scala 93:22:@39224.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_95 ( // @[package.scala 93:22:@39238.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  x553_sum x808_sum_1 ( // @[Math.scala 150:24:@39265.4]
    .clock(x808_sum_1_clock),
    .reset(x808_sum_1_reset),
    .io_a(x808_sum_1_io_a),
    .io_b(x808_sum_1_io_b),
    .io_flow(x808_sum_1_io_flow),
    .io_result(x808_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_96 ( // @[package.scala 93:22:@39275.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_97 ( // @[package.scala 93:22:@39289.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x553_sum x815_sum_1 ( // @[Math.scala 150:24:@39316.4]
    .clock(x815_sum_1_clock),
    .reset(x815_sum_1_reset),
    .io_a(x815_sum_1_io_a),
    .io_b(x815_sum_1_io_b),
    .io_flow(x815_sum_1_io_flow),
    .io_result(x815_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_98 ( // @[package.scala 93:22:@39326.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_195 RetimeWrapper_99 ( // @[package.scala 93:22:@39340.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x825_x17 x825_x17_1 ( // @[Math.scala 150:24:@39386.4]
    .clock(x825_x17_1_clock),
    .reset(x825_x17_1_reset),
    .io_a(x825_x17_1_io_a),
    .io_b(x825_x17_1_io_b),
    .io_flow(x825_x17_1_io_flow),
    .io_result(x825_x17_1_io_result)
  );
  x825_x17 x826_x18_1 ( // @[Math.scala 150:24:@39396.4]
    .clock(x826_x18_1_clock),
    .reset(x826_x18_1_reset),
    .io_a(x826_x18_1_io_a),
    .io_b(x826_x18_1_io_b),
    .io_flow(x826_x18_1_io_flow),
    .io_result(x826_x18_1_io_result)
  );
  x825_x17 x827_x17_1 ( // @[Math.scala 150:24:@39406.4]
    .clock(x827_x17_1_clock),
    .reset(x827_x17_1_reset),
    .io_a(x827_x17_1_io_a),
    .io_b(x827_x17_1_io_b),
    .io_flow(x827_x17_1_io_flow),
    .io_result(x827_x17_1_io_result)
  );
  x825_x17 x828_x18_1 ( // @[Math.scala 150:24:@39416.4]
    .clock(x828_x18_1_clock),
    .reset(x828_x18_1_reset),
    .io_a(x828_x18_1_io_a),
    .io_b(x828_x18_1_io_b),
    .io_flow(x828_x18_1_io_flow),
    .io_result(x828_x18_1_io_result)
  );
  x829_x17 x829_x17_1 ( // @[Math.scala 150:24:@39426.4]
    .io_a(x829_x17_1_io_a),
    .io_b(x829_x17_1_io_b),
    .io_result(x829_x17_1_io_result)
  );
  x829_x17 x830_x18_1 ( // @[Math.scala 150:24:@39436.4]
    .io_a(x830_x18_1_io_a),
    .io_b(x830_x18_1_io_b),
    .io_result(x830_x18_1_io_result)
  );
  x829_x17 x831_x17_1 ( // @[Math.scala 150:24:@39446.4]
    .io_a(x831_x17_1_io_a),
    .io_b(x831_x17_1_io_b),
    .io_result(x831_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_100 ( // @[package.scala 93:22:@39456.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  x829_x17 x832_sum_1 ( // @[Math.scala 150:24:@39465.4]
    .io_a(x832_sum_1_io_a),
    .io_b(x832_sum_1_io_b),
    .io_result(x832_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_101 ( // @[package.scala 93:22:@39479.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_102 ( // @[package.scala 93:22:@39489.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  x834_sub x834_sub_1 ( // @[Math.scala 191:24:@39498.4]
    .io_a(x834_sub_1_io_a),
    .io_b(x834_sub_1_io_b),
    .io_result(x834_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_103 ( // @[package.scala 93:22:@39523.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  x838_div x838_div_1 ( // @[Math.scala 327:24:@39534.4]
    .clock(x838_div_1_clock),
    .reset(x838_div_1_reset),
    .io_a(x838_div_1_io_a),
    .io_flow(x838_div_1_io_flow),
    .io_result(x838_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_104 ( // @[package.scala 93:22:@39544.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x829_x17 x839_sum_1 ( // @[Math.scala 150:24:@39553.4]
    .io_a(x839_sum_1_io_a),
    .io_b(x839_sum_1_io_b),
    .io_result(x839_sum_1_io_result)
  );
  RetimeWrapper_298 RetimeWrapper_105 ( // @[package.scala 93:22:@39563.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_299 RetimeWrapper_106 ( // @[package.scala 93:22:@39572.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x825_x17 x846_x17_1 ( // @[Math.scala 150:24:@39611.4]
    .clock(x846_x17_1_clock),
    .reset(x846_x17_1_reset),
    .io_a(x846_x17_1_io_a),
    .io_b(x846_x17_1_io_b),
    .io_flow(x846_x17_1_io_flow),
    .io_result(x846_x17_1_io_result)
  );
  x825_x17 x847_x18_1 ( // @[Math.scala 150:24:@39621.4]
    .clock(x847_x18_1_clock),
    .reset(x847_x18_1_reset),
    .io_a(x847_x18_1_io_a),
    .io_b(x847_x18_1_io_b),
    .io_flow(x847_x18_1_io_flow),
    .io_result(x847_x18_1_io_result)
  );
  x825_x17 x848_x17_1 ( // @[Math.scala 150:24:@39631.4]
    .clock(x848_x17_1_clock),
    .reset(x848_x17_1_reset),
    .io_a(x848_x17_1_io_a),
    .io_b(x848_x17_1_io_b),
    .io_flow(x848_x17_1_io_flow),
    .io_result(x848_x17_1_io_result)
  );
  x825_x17 x849_x18_1 ( // @[Math.scala 150:24:@39641.4]
    .clock(x849_x18_1_clock),
    .reset(x849_x18_1_reset),
    .io_a(x849_x18_1_io_a),
    .io_b(x849_x18_1_io_b),
    .io_flow(x849_x18_1_io_flow),
    .io_result(x849_x18_1_io_result)
  );
  x829_x17 x850_x17_1 ( // @[Math.scala 150:24:@39651.4]
    .io_a(x850_x17_1_io_a),
    .io_b(x850_x17_1_io_b),
    .io_result(x850_x17_1_io_result)
  );
  x829_x17 x851_x18_1 ( // @[Math.scala 150:24:@39661.4]
    .io_a(x851_x18_1_io_a),
    .io_b(x851_x18_1_io_b),
    .io_result(x851_x18_1_io_result)
  );
  x829_x17 x852_x17_1 ( // @[Math.scala 150:24:@39671.4]
    .io_a(x852_x17_1_io_a),
    .io_b(x852_x17_1_io_b),
    .io_result(x852_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_107 ( // @[package.scala 93:22:@39681.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x829_x17 x853_sum_1 ( // @[Math.scala 150:24:@39690.4]
    .io_a(x853_sum_1_io_a),
    .io_b(x853_sum_1_io_b),
    .io_result(x853_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_108 ( // @[package.scala 93:22:@39704.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_109 ( // @[package.scala 93:22:@39714.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  x834_sub x855_sub_1 ( // @[Math.scala 191:24:@39723.4]
    .io_a(x855_sub_1_io_a),
    .io_b(x855_sub_1_io_b),
    .io_result(x855_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_110 ( // @[package.scala 93:22:@39748.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  x838_div x859_div_1 ( // @[Math.scala 327:24:@39759.4]
    .clock(x859_div_1_clock),
    .reset(x859_div_1_reset),
    .io_a(x859_div_1_io_a),
    .io_flow(x859_div_1_io_flow),
    .io_result(x859_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_111 ( // @[package.scala 93:22:@39769.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  x829_x17 x860_sum_1 ( // @[Math.scala 150:24:@39778.4]
    .io_a(x860_sum_1_io_a),
    .io_b(x860_sum_1_io_b),
    .io_result(x860_sum_1_io_result)
  );
  RetimeWrapper_298 RetimeWrapper_112 ( // @[package.scala 93:22:@39788.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_299 RetimeWrapper_113 ( // @[package.scala 93:22:@39797.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  x825_x17 x866_x17_1 ( // @[Math.scala 150:24:@39829.4]
    .clock(x866_x17_1_clock),
    .reset(x866_x17_1_reset),
    .io_a(x866_x17_1_io_a),
    .io_b(x866_x17_1_io_b),
    .io_flow(x866_x17_1_io_flow),
    .io_result(x866_x17_1_io_result)
  );
  x825_x17 x867_x18_1 ( // @[Math.scala 150:24:@39839.4]
    .clock(x867_x18_1_clock),
    .reset(x867_x18_1_reset),
    .io_a(x867_x18_1_io_a),
    .io_b(x867_x18_1_io_b),
    .io_flow(x867_x18_1_io_flow),
    .io_result(x867_x18_1_io_result)
  );
  x825_x17 x868_x17_1 ( // @[Math.scala 150:24:@39849.4]
    .clock(x868_x17_1_clock),
    .reset(x868_x17_1_reset),
    .io_a(x868_x17_1_io_a),
    .io_b(x868_x17_1_io_b),
    .io_flow(x868_x17_1_io_flow),
    .io_result(x868_x17_1_io_result)
  );
  x825_x17 x869_x18_1 ( // @[Math.scala 150:24:@39859.4]
    .clock(x869_x18_1_clock),
    .reset(x869_x18_1_reset),
    .io_a(x869_x18_1_io_a),
    .io_b(x869_x18_1_io_b),
    .io_flow(x869_x18_1_io_flow),
    .io_result(x869_x18_1_io_result)
  );
  x829_x17 x870_x17_1 ( // @[Math.scala 150:24:@39869.4]
    .io_a(x870_x17_1_io_a),
    .io_b(x870_x17_1_io_b),
    .io_result(x870_x17_1_io_result)
  );
  x829_x17 x871_x18_1 ( // @[Math.scala 150:24:@39879.4]
    .io_a(x871_x18_1_io_a),
    .io_b(x871_x18_1_io_b),
    .io_result(x871_x18_1_io_result)
  );
  x829_x17 x872_x17_1 ( // @[Math.scala 150:24:@39889.4]
    .io_a(x872_x17_1_io_a),
    .io_b(x872_x17_1_io_b),
    .io_result(x872_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_114 ( // @[package.scala 93:22:@39899.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  x829_x17 x873_sum_1 ( // @[Math.scala 150:24:@39908.4]
    .io_a(x873_sum_1_io_a),
    .io_b(x873_sum_1_io_b),
    .io_result(x873_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_115 ( // @[package.scala 93:22:@39922.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_116 ( // @[package.scala 93:22:@39932.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  x834_sub x875_sub_1 ( // @[Math.scala 191:24:@39941.4]
    .io_a(x875_sub_1_io_a),
    .io_b(x875_sub_1_io_b),
    .io_result(x875_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_117 ( // @[package.scala 93:22:@39966.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  x838_div x879_div_1 ( // @[Math.scala 327:24:@39977.4]
    .clock(x879_div_1_clock),
    .reset(x879_div_1_reset),
    .io_a(x879_div_1_io_a),
    .io_flow(x879_div_1_io_flow),
    .io_result(x879_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_118 ( // @[package.scala 93:22:@39987.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  x829_x17 x880_sum_1 ( // @[Math.scala 150:24:@39998.4]
    .io_a(x880_sum_1_io_a),
    .io_b(x880_sum_1_io_b),
    .io_result(x880_sum_1_io_result)
  );
  RetimeWrapper_298 RetimeWrapper_119 ( // @[package.scala 93:22:@40008.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_299 RetimeWrapper_120 ( // @[package.scala 93:22:@40017.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  x825_x17 x886_x17_1 ( // @[Math.scala 150:24:@40049.4]
    .clock(x886_x17_1_clock),
    .reset(x886_x17_1_reset),
    .io_a(x886_x17_1_io_a),
    .io_b(x886_x17_1_io_b),
    .io_flow(x886_x17_1_io_flow),
    .io_result(x886_x17_1_io_result)
  );
  x825_x17 x887_x18_1 ( // @[Math.scala 150:24:@40059.4]
    .clock(x887_x18_1_clock),
    .reset(x887_x18_1_reset),
    .io_a(x887_x18_1_io_a),
    .io_b(x887_x18_1_io_b),
    .io_flow(x887_x18_1_io_flow),
    .io_result(x887_x18_1_io_result)
  );
  x825_x17 x888_x17_1 ( // @[Math.scala 150:24:@40069.4]
    .clock(x888_x17_1_clock),
    .reset(x888_x17_1_reset),
    .io_a(x888_x17_1_io_a),
    .io_b(x888_x17_1_io_b),
    .io_flow(x888_x17_1_io_flow),
    .io_result(x888_x17_1_io_result)
  );
  x825_x17 x889_x18_1 ( // @[Math.scala 150:24:@40079.4]
    .clock(x889_x18_1_clock),
    .reset(x889_x18_1_reset),
    .io_a(x889_x18_1_io_a),
    .io_b(x889_x18_1_io_b),
    .io_flow(x889_x18_1_io_flow),
    .io_result(x889_x18_1_io_result)
  );
  x829_x17 x890_x17_1 ( // @[Math.scala 150:24:@40089.4]
    .io_a(x890_x17_1_io_a),
    .io_b(x890_x17_1_io_b),
    .io_result(x890_x17_1_io_result)
  );
  x829_x17 x891_x18_1 ( // @[Math.scala 150:24:@40099.4]
    .io_a(x891_x18_1_io_a),
    .io_b(x891_x18_1_io_b),
    .io_result(x891_x18_1_io_result)
  );
  x829_x17 x892_x17_1 ( // @[Math.scala 150:24:@40109.4]
    .io_a(x892_x17_1_io_a),
    .io_b(x892_x17_1_io_b),
    .io_result(x892_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_121 ( // @[package.scala 93:22:@40119.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  x829_x17 x893_sum_1 ( // @[Math.scala 150:24:@40128.4]
    .io_a(x893_sum_1_io_a),
    .io_b(x893_sum_1_io_b),
    .io_result(x893_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_122 ( // @[package.scala 93:22:@40142.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_123 ( // @[package.scala 93:22:@40152.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  x834_sub x895_sub_1 ( // @[Math.scala 191:24:@40161.4]
    .io_a(x895_sub_1_io_a),
    .io_b(x895_sub_1_io_b),
    .io_result(x895_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_124 ( // @[package.scala 93:22:@40186.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  x838_div x899_div_1 ( // @[Math.scala 327:24:@40197.4]
    .clock(x899_div_1_clock),
    .reset(x899_div_1_reset),
    .io_a(x899_div_1_io_a),
    .io_flow(x899_div_1_io_flow),
    .io_result(x899_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_125 ( // @[package.scala 93:22:@40207.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  x829_x17 x900_sum_1 ( // @[Math.scala 150:24:@40216.4]
    .io_a(x900_sum_1_io_a),
    .io_b(x900_sum_1_io_b),
    .io_result(x900_sum_1_io_result)
  );
  RetimeWrapper_298 RetimeWrapper_126 ( // @[package.scala 93:22:@40226.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_299 RetimeWrapper_127 ( // @[package.scala 93:22:@40235.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  x825_x17 x905_x17_1 ( // @[Math.scala 150:24:@40262.4]
    .clock(x905_x17_1_clock),
    .reset(x905_x17_1_reset),
    .io_a(x905_x17_1_io_a),
    .io_b(x905_x17_1_io_b),
    .io_flow(x905_x17_1_io_flow),
    .io_result(x905_x17_1_io_result)
  );
  x825_x17 x906_x18_1 ( // @[Math.scala 150:24:@40272.4]
    .clock(x906_x18_1_clock),
    .reset(x906_x18_1_reset),
    .io_a(x906_x18_1_io_a),
    .io_b(x906_x18_1_io_b),
    .io_flow(x906_x18_1_io_flow),
    .io_result(x906_x18_1_io_result)
  );
  x825_x17 x907_x17_1 ( // @[Math.scala 150:24:@40282.4]
    .clock(x907_x17_1_clock),
    .reset(x907_x17_1_reset),
    .io_a(x907_x17_1_io_a),
    .io_b(x907_x17_1_io_b),
    .io_flow(x907_x17_1_io_flow),
    .io_result(x907_x17_1_io_result)
  );
  x825_x17 x908_x18_1 ( // @[Math.scala 150:24:@40292.4]
    .clock(x908_x18_1_clock),
    .reset(x908_x18_1_reset),
    .io_a(x908_x18_1_io_a),
    .io_b(x908_x18_1_io_b),
    .io_flow(x908_x18_1_io_flow),
    .io_result(x908_x18_1_io_result)
  );
  x829_x17 x909_x17_1 ( // @[Math.scala 150:24:@40302.4]
    .io_a(x909_x17_1_io_a),
    .io_b(x909_x17_1_io_b),
    .io_result(x909_x17_1_io_result)
  );
  x829_x17 x910_x18_1 ( // @[Math.scala 150:24:@40312.4]
    .io_a(x910_x18_1_io_a),
    .io_b(x910_x18_1_io_b),
    .io_result(x910_x18_1_io_result)
  );
  x829_x17 x911_x17_1 ( // @[Math.scala 150:24:@40322.4]
    .io_a(x911_x17_1_io_a),
    .io_b(x911_x17_1_io_b),
    .io_result(x911_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_128 ( // @[package.scala 93:22:@40332.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  x829_x17 x912_sum_1 ( // @[Math.scala 150:24:@40341.4]
    .io_a(x912_sum_1_io_a),
    .io_b(x912_sum_1_io_b),
    .io_result(x912_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_129 ( // @[package.scala 93:22:@40355.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_130 ( // @[package.scala 93:22:@40365.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  x834_sub x914_sub_1 ( // @[Math.scala 191:24:@40374.4]
    .io_a(x914_sub_1_io_a),
    .io_b(x914_sub_1_io_b),
    .io_result(x914_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_131 ( // @[package.scala 93:22:@40399.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  x838_div x918_div_1 ( // @[Math.scala 327:24:@40412.4]
    .clock(x918_div_1_clock),
    .reset(x918_div_1_reset),
    .io_a(x918_div_1_io_a),
    .io_flow(x918_div_1_io_flow),
    .io_result(x918_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_132 ( // @[package.scala 93:22:@40422.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  x829_x17 x919_sum_1 ( // @[Math.scala 150:24:@40431.4]
    .io_a(x919_sum_1_io_a),
    .io_b(x919_sum_1_io_b),
    .io_result(x919_sum_1_io_result)
  );
  RetimeWrapper_299 RetimeWrapper_133 ( // @[package.scala 93:22:@40441.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_298 RetimeWrapper_134 ( // @[package.scala 93:22:@40450.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  x825_x17 x923_x17_1 ( // @[Math.scala 150:24:@40472.4]
    .clock(x923_x17_1_clock),
    .reset(x923_x17_1_reset),
    .io_a(x923_x17_1_io_a),
    .io_b(x923_x17_1_io_b),
    .io_flow(x923_x17_1_io_flow),
    .io_result(x923_x17_1_io_result)
  );
  x825_x17 x924_x18_1 ( // @[Math.scala 150:24:@40482.4]
    .clock(x924_x18_1_clock),
    .reset(x924_x18_1_reset),
    .io_a(x924_x18_1_io_a),
    .io_b(x924_x18_1_io_b),
    .io_flow(x924_x18_1_io_flow),
    .io_result(x924_x18_1_io_result)
  );
  x825_x17 x925_x17_1 ( // @[Math.scala 150:24:@40492.4]
    .clock(x925_x17_1_clock),
    .reset(x925_x17_1_reset),
    .io_a(x925_x17_1_io_a),
    .io_b(x925_x17_1_io_b),
    .io_flow(x925_x17_1_io_flow),
    .io_result(x925_x17_1_io_result)
  );
  x825_x17 x926_x18_1 ( // @[Math.scala 150:24:@40502.4]
    .clock(x926_x18_1_clock),
    .reset(x926_x18_1_reset),
    .io_a(x926_x18_1_io_a),
    .io_b(x926_x18_1_io_b),
    .io_flow(x926_x18_1_io_flow),
    .io_result(x926_x18_1_io_result)
  );
  x829_x17 x927_x17_1 ( // @[Math.scala 150:24:@40512.4]
    .io_a(x927_x17_1_io_a),
    .io_b(x927_x17_1_io_b),
    .io_result(x927_x17_1_io_result)
  );
  x829_x17 x928_x18_1 ( // @[Math.scala 150:24:@40522.4]
    .io_a(x928_x18_1_io_a),
    .io_b(x928_x18_1_io_b),
    .io_result(x928_x18_1_io_result)
  );
  x829_x17 x929_x17_1 ( // @[Math.scala 150:24:@40532.4]
    .io_a(x929_x17_1_io_a),
    .io_b(x929_x17_1_io_b),
    .io_result(x929_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_135 ( // @[package.scala 93:22:@40542.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  x829_x17 x930_sum_1 ( // @[Math.scala 150:24:@40551.4]
    .io_a(x930_sum_1_io_a),
    .io_b(x930_sum_1_io_b),
    .io_result(x930_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_136 ( // @[package.scala 93:22:@40565.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_137 ( // @[package.scala 93:22:@40575.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  x834_sub x932_sub_1 ( // @[Math.scala 191:24:@40584.4]
    .io_a(x932_sub_1_io_a),
    .io_b(x932_sub_1_io_b),
    .io_result(x932_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_138 ( // @[package.scala 93:22:@40609.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  x838_div x936_div_1 ( // @[Math.scala 327:24:@40620.4]
    .clock(x936_div_1_clock),
    .reset(x936_div_1_reset),
    .io_a(x936_div_1_io_a),
    .io_flow(x936_div_1_io_flow),
    .io_result(x936_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_139 ( // @[package.scala 93:22:@40630.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  x829_x17 x937_sum_1 ( // @[Math.scala 150:24:@40639.4]
    .io_a(x937_sum_1_io_a),
    .io_b(x937_sum_1_io_b),
    .io_result(x937_sum_1_io_result)
  );
  RetimeWrapper_299 RetimeWrapper_140 ( // @[package.scala 93:22:@40649.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_298 RetimeWrapper_141 ( // @[package.scala 93:22:@40658.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  x825_x17 x941_x17_1 ( // @[Math.scala 150:24:@40680.4]
    .clock(x941_x17_1_clock),
    .reset(x941_x17_1_reset),
    .io_a(x941_x17_1_io_a),
    .io_b(x941_x17_1_io_b),
    .io_flow(x941_x17_1_io_flow),
    .io_result(x941_x17_1_io_result)
  );
  x825_x17 x942_x18_1 ( // @[Math.scala 150:24:@40690.4]
    .clock(x942_x18_1_clock),
    .reset(x942_x18_1_reset),
    .io_a(x942_x18_1_io_a),
    .io_b(x942_x18_1_io_b),
    .io_flow(x942_x18_1_io_flow),
    .io_result(x942_x18_1_io_result)
  );
  x825_x17 x943_x17_1 ( // @[Math.scala 150:24:@40700.4]
    .clock(x943_x17_1_clock),
    .reset(x943_x17_1_reset),
    .io_a(x943_x17_1_io_a),
    .io_b(x943_x17_1_io_b),
    .io_flow(x943_x17_1_io_flow),
    .io_result(x943_x17_1_io_result)
  );
  x825_x17 x944_x18_1 ( // @[Math.scala 150:24:@40710.4]
    .clock(x944_x18_1_clock),
    .reset(x944_x18_1_reset),
    .io_a(x944_x18_1_io_a),
    .io_b(x944_x18_1_io_b),
    .io_flow(x944_x18_1_io_flow),
    .io_result(x944_x18_1_io_result)
  );
  x829_x17 x945_x17_1 ( // @[Math.scala 150:24:@40720.4]
    .io_a(x945_x17_1_io_a),
    .io_b(x945_x17_1_io_b),
    .io_result(x945_x17_1_io_result)
  );
  x829_x17 x946_x18_1 ( // @[Math.scala 150:24:@40730.4]
    .io_a(x946_x18_1_io_a),
    .io_b(x946_x18_1_io_b),
    .io_result(x946_x18_1_io_result)
  );
  x829_x17 x947_x17_1 ( // @[Math.scala 150:24:@40740.4]
    .io_a(x947_x17_1_io_a),
    .io_b(x947_x17_1_io_b),
    .io_result(x947_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_142 ( // @[package.scala 93:22:@40750.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  x829_x17 x948_sum_1 ( // @[Math.scala 150:24:@40759.4]
    .io_a(x948_sum_1_io_a),
    .io_b(x948_sum_1_io_b),
    .io_result(x948_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_143 ( // @[package.scala 93:22:@40773.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_144 ( // @[package.scala 93:22:@40783.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  x834_sub x950_sub_1 ( // @[Math.scala 191:24:@40792.4]
    .io_a(x950_sub_1_io_a),
    .io_b(x950_sub_1_io_b),
    .io_result(x950_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_145 ( // @[package.scala 93:22:@40817.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  x838_div x954_div_1 ( // @[Math.scala 327:24:@40828.4]
    .clock(x954_div_1_clock),
    .reset(x954_div_1_reset),
    .io_a(x954_div_1_io_a),
    .io_flow(x954_div_1_io_flow),
    .io_result(x954_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_146 ( // @[package.scala 93:22:@40838.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  x829_x17 x955_sum_1 ( // @[Math.scala 150:24:@40849.4]
    .io_a(x955_sum_1_io_a),
    .io_b(x955_sum_1_io_b),
    .io_result(x955_sum_1_io_result)
  );
  RetimeWrapper_299 RetimeWrapper_147 ( // @[package.scala 93:22:@40859.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_298 RetimeWrapper_148 ( // @[package.scala 93:22:@40868.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  x825_x17 x960_x17_1 ( // @[Math.scala 150:24:@40895.4]
    .clock(x960_x17_1_clock),
    .reset(x960_x17_1_reset),
    .io_a(x960_x17_1_io_a),
    .io_b(x960_x17_1_io_b),
    .io_flow(x960_x17_1_io_flow),
    .io_result(x960_x17_1_io_result)
  );
  x825_x17 x961_x18_1 ( // @[Math.scala 150:24:@40905.4]
    .clock(x961_x18_1_clock),
    .reset(x961_x18_1_reset),
    .io_a(x961_x18_1_io_a),
    .io_b(x961_x18_1_io_b),
    .io_flow(x961_x18_1_io_flow),
    .io_result(x961_x18_1_io_result)
  );
  x825_x17 x962_x17_1 ( // @[Math.scala 150:24:@40915.4]
    .clock(x962_x17_1_clock),
    .reset(x962_x17_1_reset),
    .io_a(x962_x17_1_io_a),
    .io_b(x962_x17_1_io_b),
    .io_flow(x962_x17_1_io_flow),
    .io_result(x962_x17_1_io_result)
  );
  x825_x17 x963_x18_1 ( // @[Math.scala 150:24:@40925.4]
    .clock(x963_x18_1_clock),
    .reset(x963_x18_1_reset),
    .io_a(x963_x18_1_io_a),
    .io_b(x963_x18_1_io_b),
    .io_flow(x963_x18_1_io_flow),
    .io_result(x963_x18_1_io_result)
  );
  x829_x17 x964_x17_1 ( // @[Math.scala 150:24:@40935.4]
    .io_a(x964_x17_1_io_a),
    .io_b(x964_x17_1_io_b),
    .io_result(x964_x17_1_io_result)
  );
  x829_x17 x965_x18_1 ( // @[Math.scala 150:24:@40945.4]
    .io_a(x965_x18_1_io_a),
    .io_b(x965_x18_1_io_b),
    .io_result(x965_x18_1_io_result)
  );
  x829_x17 x966_x17_1 ( // @[Math.scala 150:24:@40955.4]
    .io_a(x966_x17_1_io_a),
    .io_b(x966_x17_1_io_b),
    .io_result(x966_x17_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_149 ( // @[package.scala 93:22:@40965.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  x829_x17 x967_sum_1 ( // @[Math.scala 150:24:@40974.4]
    .io_a(x967_sum_1_io_a),
    .io_b(x967_sum_1_io_b),
    .io_result(x967_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_150 ( // @[package.scala 93:22:@40988.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_294 RetimeWrapper_151 ( // @[package.scala 93:22:@40998.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  x834_sub x969_sub_1 ( // @[Math.scala 191:24:@41007.4]
    .io_a(x969_sub_1_io_a),
    .io_b(x969_sub_1_io_b),
    .io_result(x969_sub_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_152 ( // @[package.scala 93:22:@41032.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  x838_div x973_div_1 ( // @[Math.scala 327:24:@41043.4]
    .clock(x973_div_1_clock),
    .reset(x973_div_1_reset),
    .io_a(x973_div_1_io_a),
    .io_flow(x973_div_1_io_flow),
    .io_result(x973_div_1_io_result)
  );
  RetimeWrapper_297 RetimeWrapper_153 ( // @[package.scala 93:22:@41053.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  x829_x17 x974_sum_1 ( // @[Math.scala 150:24:@41062.4]
    .io_a(x974_sum_1_io_a),
    .io_b(x974_sum_1_io_b),
    .io_result(x974_sum_1_io_result)
  );
  RetimeWrapper_299 RetimeWrapper_154 ( // @[package.scala 93:22:@41072.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_298 RetimeWrapper_155 ( // @[package.scala 93:22:@41081.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_384 RetimeWrapper_156 ( // @[package.scala 93:22:@41111.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_157 ( // @[package.scala 93:22:@41120.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_158 ( // @[package.scala 93:22:@41129.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_159 ( // @[package.scala 93:22:@41138.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  assign b537 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 62:18:@36708.4]
  assign b538 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 63:18:@36709.4]
  assign _T_206 = b537 & b538; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 68:30:@36924.4]
  assign _T_207 = _T_206 & io_sigsIn_datapathEn; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 68:37:@36925.4]
  assign _T_211 = io_in_x526_TID == 8'h0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:76:@36930.4]
  assign _T_212 = _T_207 & _T_211; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:62:@36931.4]
  assign _T_214 = io_in_x526_TDEST == 8'h0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:101:@36932.4]
  assign x1058_x540_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@36941.4 package.scala 96:25:@36942.4]
  assign b535_number = __io_result; // @[Math.scala 712:22:@36693.4 Math.scala 713:14:@36694.4]
  assign _T_254 = $signed(b535_number); // @[Math.scala 499:52:@36969.4]
  assign x544 = $signed(32'sh1) == $signed(_T_254); // @[Math.scala 499:44:@36977.4]
  assign x545 = $signed(32'sh2) == $signed(_T_254); // @[Math.scala 499:44:@36984.4]
  assign x546 = $signed(32'sh3) == $signed(_T_254); // @[Math.scala 499:44:@36991.4]
  assign _T_301 = x544 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@37003.4]
  assign _T_303 = x545 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@37004.4]
  assign _T_305 = x546 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@37005.4]
  assign _T_307 = _T_301 | _T_303; // @[Mux.scala 19:72:@37007.4]
  assign x547_number = _T_307 | _T_305; // @[Mux.scala 19:72:@37008.4]
  assign _T_319 = $signed(x547_number); // @[Math.scala 406:49:@37018.4]
  assign _T_321 = $signed(_T_319) & $signed(32'sh3); // @[Math.scala 406:56:@37020.4]
  assign _T_322 = $signed(_T_321); // @[Math.scala 406:56:@37021.4]
  assign _T_327 = x547_number[31]; // @[FixedPoint.scala 50:25:@37027.4]
  assign _T_331 = _T_327 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37029.4]
  assign _T_332 = x547_number[31:2]; // @[FixedPoint.scala 18:52:@37030.4]
  assign b536_number = __1_io_result; // @[Math.scala 712:22:@36705.4 Math.scala 713:14:@36706.4]
  assign _T_337 = b536_number[31]; // @[FixedPoint.scala 50:25:@37036.4]
  assign _T_341 = _T_337 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37038.4]
  assign _T_342 = b536_number[31:2]; // @[FixedPoint.scala 18:52:@37039.4]
  assign _T_367 = ~ io_sigsIn_break; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:101:@37100.4]
  assign _T_371 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@37108.4 package.scala 96:25:@37109.4]
  assign _T_373 = io_rr ? _T_371 : 1'h0; // @[implicits.scala 55:10:@37110.4]
  assign _T_374 = _T_367 & _T_373; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:118:@37111.4]
  assign _T_376 = _T_374 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:205:@37113.4]
  assign _T_377 = _T_376 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:224:@37114.4]
  assign x1060_b537_D8 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@37068.4 package.scala 96:25:@37069.4]
  assign _T_378 = _T_377 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 113:250:@37115.4]
  assign x1059_b538_D8 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37059.4 package.scala 96:25:@37060.4]
  assign x559_rdcol_number = x559_rdcol_1_io_result; // @[Math.scala 154:22:@37132.4 Math.scala 155:14:@37133.4]
  assign _T_391 = x559_rdcol_number[31]; // @[FixedPoint.scala 50:25:@37139.4]
  assign _T_395 = _T_391 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37141.4]
  assign _T_396 = x559_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@37142.4]
  assign _T_419 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@37193.4 package.scala 96:25:@37194.4]
  assign _T_421 = io_rr ? _T_419 : 1'h0; // @[implicits.scala 55:10:@37195.4]
  assign _T_422 = _T_367 & _T_421; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:118:@37196.4]
  assign _T_424 = _T_422 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:205:@37198.4]
  assign _T_425 = _T_424 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:224:@37199.4]
  assign _T_426 = _T_425 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 132:250:@37200.4]
  assign x568_rdcol_number = x568_rdcol_1_io_result; // @[Math.scala 154:22:@37217.4 Math.scala 155:14:@37218.4]
  assign _T_439 = x568_rdcol_number[31]; // @[FixedPoint.scala 50:25:@37224.4]
  assign _T_443 = _T_439 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37226.4]
  assign _T_444 = x568_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@37227.4]
  assign _T_464 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@37269.4 package.scala 96:25:@37270.4]
  assign _T_466 = io_rr ? _T_464 : 1'h0; // @[implicits.scala 55:10:@37271.4]
  assign _T_467 = _T_367 & _T_466; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:118:@37272.4]
  assign _T_469 = _T_467 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:205:@37274.4]
  assign _T_470 = _T_469 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:224:@37275.4]
  assign _T_471 = _T_470 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 149:250:@37276.4]
  assign x577_rdcol_number = x577_rdcol_1_io_result; // @[Math.scala 154:22:@37293.4 Math.scala 155:14:@37294.4]
  assign _T_484 = x577_rdcol_number[31]; // @[FixedPoint.scala 50:25:@37300.4]
  assign _T_488 = _T_484 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37302.4]
  assign _T_489 = x577_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@37303.4]
  assign _T_509 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@37345.4 package.scala 96:25:@37346.4]
  assign _T_511 = io_rr ? _T_509 : 1'h0; // @[implicits.scala 55:10:@37347.4]
  assign _T_512 = _T_367 & _T_511; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:118:@37348.4]
  assign _T_514 = _T_512 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:205:@37350.4]
  assign _T_515 = _T_514 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:224:@37351.4]
  assign _T_516 = _T_515 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 166:250:@37352.4]
  assign x586_rdrow_number = x586_rdrow_1_io_result; // @[Math.scala 154:22:@37369.4 Math.scala 155:14:@37370.4]
  assign _T_531 = $signed(x586_rdrow_number); // @[Math.scala 499:52:@37376.4]
  assign x588 = $signed(32'sh1) == $signed(_T_531); // @[Math.scala 499:44:@37384.4]
  assign x589 = $signed(32'sh2) == $signed(_T_531); // @[Math.scala 499:44:@37391.4]
  assign x590 = $signed(32'sh3) == $signed(_T_531); // @[Math.scala 499:44:@37398.4]
  assign _T_578 = x588 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@37410.4]
  assign _T_580 = x589 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@37411.4]
  assign _T_582 = x590 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@37412.4]
  assign _T_584 = _T_578 | _T_580; // @[Mux.scala 19:72:@37414.4]
  assign x591_number = _T_584 | _T_582; // @[Mux.scala 19:72:@37415.4]
  assign _T_598 = $signed(x591_number); // @[Math.scala 406:49:@37427.4]
  assign _T_600 = $signed(_T_598) & $signed(32'sh3); // @[Math.scala 406:56:@37429.4]
  assign _T_601 = $signed(_T_600); // @[Math.scala 406:56:@37430.4]
  assign _T_606 = x591_number[31]; // @[FixedPoint.scala 50:25:@37436.4]
  assign _T_610 = _T_606 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37438.4]
  assign _T_611 = x591_number[31:2]; // @[FixedPoint.scala 18:52:@37439.4]
  assign _T_637 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@37499.4 package.scala 96:25:@37500.4]
  assign _T_639 = io_rr ? _T_637 : 1'h0; // @[implicits.scala 55:10:@37501.4]
  assign _T_640 = _T_367 & _T_639; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:166:@37502.4]
  assign _T_642 = _T_640 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:253:@37504.4]
  assign _T_643 = _T_642 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:272:@37505.4]
  assign _T_644 = _T_643 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 207:298:@37506.4]
  assign _T_665 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@37554.4 package.scala 96:25:@37555.4]
  assign _T_667 = io_rr ? _T_665 : 1'h0; // @[implicits.scala 55:10:@37556.4]
  assign _T_668 = _T_367 & _T_667; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:166:@37557.4]
  assign _T_670 = _T_668 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:253:@37559.4]
  assign _T_671 = _T_670 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:272:@37560.4]
  assign _T_672 = _T_671 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 220:298:@37561.4]
  assign _T_693 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@37609.4 package.scala 96:25:@37610.4]
  assign _T_695 = io_rr ? _T_693 : 1'h0; // @[implicits.scala 55:10:@37611.4]
  assign _T_696 = _T_367 & _T_695; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:166:@37612.4]
  assign _T_698 = _T_696 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:253:@37614.4]
  assign _T_699 = _T_698 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:272:@37615.4]
  assign _T_700 = _T_699 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 233:298:@37616.4]
  assign _T_721 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@37664.4 package.scala 96:25:@37665.4]
  assign _T_723 = io_rr ? _T_721 : 1'h0; // @[implicits.scala 55:10:@37666.4]
  assign _T_724 = _T_367 & _T_723; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:166:@37667.4]
  assign _T_726 = _T_724 & _T_367; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:253:@37669.4]
  assign _T_727 = _T_726 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:272:@37670.4]
  assign _T_728 = _T_727 & x1060_b537_D8; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 246:298:@37671.4]
  assign x1081_x586_rdrow_D11_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@37685.4 package.scala 96:25:@37686.4]
  assign _T_740 = $signed(x1081_x586_rdrow_D11_number); // @[Math.scala 406:49:@37692.4]
  assign _T_742 = $signed(_T_740) & $signed(32'sh3); // @[Math.scala 406:56:@37694.4]
  assign _T_743 = $signed(_T_742); // @[Math.scala 406:56:@37695.4]
  assign x1050_number = $unsigned(_T_743); // @[implicits.scala 133:21:@37696.4]
  assign x617 = $signed(_T_740) < $signed(32'sh0); // @[Math.scala 465:44:@37704.4]
  assign x1082_x577_rdcol_D11_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@37712.4 package.scala 96:25:@37713.4]
  assign _T_761 = $signed(x1082_x577_rdcol_D11_number); // @[Math.scala 465:37:@37718.4]
  assign x618 = $signed(_T_761) < $signed(32'sh0); // @[Math.scala 465:44:@37720.4]
  assign x619 = x617 | x618; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 259:24:@37723.4]
  assign _T_775 = $signed(x1050_number); // @[Math.scala 406:49:@37732.4]
  assign _T_777 = $signed(_T_775) & $signed(32'sh3); // @[Math.scala 406:56:@37734.4]
  assign _T_778 = $signed(_T_777); // @[Math.scala 406:56:@37735.4]
  assign _T_783 = x1050_number[31]; // @[FixedPoint.scala 50:25:@37741.4]
  assign _T_787 = _T_783 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@37743.4]
  assign _T_788 = x1050_number[31:2]; // @[FixedPoint.scala 18:52:@37744.4]
  assign _T_823 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@37814.4 package.scala 96:25:@37815.4]
  assign _T_825 = io_rr ? _T_823 : 1'h0; // @[implicits.scala 55:10:@37816.4]
  assign _T_826 = _T_367 & _T_825; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 282:194:@37817.4]
  assign x1087_x620_D1 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@37800.4 package.scala 96:25:@37801.4]
  assign _T_827 = _T_826 & x1087_x620_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 282:282:@37818.4]
  assign x1086_b537_D13 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@37791.4 package.scala 96:25:@37792.4]
  assign _T_828 = _T_827 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 282:291:@37819.4]
  assign x1084_b538_D13 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@37773.4 package.scala 96:25:@37774.4]
  assign x1088_x568_rdcol_D11_number = RetimeWrapper_39_io_out; // @[package.scala 96:25:@37835.4 package.scala 96:25:@37836.4]
  assign _T_839 = $signed(x1088_x568_rdcol_D11_number); // @[Math.scala 465:37:@37841.4]
  assign x629 = $signed(_T_839) < $signed(32'sh0); // @[Math.scala 465:44:@37843.4]
  assign x630 = x617 | x629; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 290:24:@37846.4]
  assign _T_870 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@37890.4 package.scala 96:25:@37891.4]
  assign _T_872 = io_rr ? _T_870 : 1'h0; // @[implicits.scala 55:10:@37892.4]
  assign _T_873 = _T_367 & _T_872; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:194:@37893.4]
  assign x1090_x631_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@37876.4 package.scala 96:25:@37877.4]
  assign _T_874 = _T_873 & x1090_x631_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:282:@37894.4]
  assign _T_875 = _T_874 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:326:@37895.4]
  assign x1091_x559_rdcol_D11_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@37911.4 package.scala 96:25:@37912.4]
  assign _T_888 = $signed(x1091_x559_rdcol_D11_number); // @[Math.scala 465:37:@37919.4]
  assign x637 = $signed(_T_888) < $signed(32'sh0); // @[Math.scala 465:44:@37921.4]
  assign x638 = x617 | x637; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 319:59:@37924.4]
  assign _T_919 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@37968.4 package.scala 96:25:@37969.4]
  assign _T_921 = io_rr ? _T_919 : 1'h0; // @[implicits.scala 55:10:@37970.4]
  assign _T_922 = _T_367 & _T_921; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:194:@37971.4]
  assign x1093_x639_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@37954.4 package.scala 96:25:@37955.4]
  assign _T_923 = _T_922 & x1093_x639_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:282:@37972.4]
  assign _T_924 = _T_923 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:291:@37973.4]
  assign x1094_b536_D11_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@37989.4 package.scala 96:25:@37990.4]
  assign _T_935 = $signed(x1094_b536_D11_number); // @[Math.scala 465:37:@37995.4]
  assign x645 = $signed(_T_935) < $signed(32'sh0); // @[Math.scala 465:44:@37997.4]
  assign x1095_x645_D1 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@38005.4 package.scala 96:25:@38006.4]
  assign x646 = x617 | x1095_x645_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 342:59:@38009.4]
  assign _T_969 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@38053.4 package.scala 96:25:@38054.4]
  assign _T_971 = io_rr ? _T_969 : 1'h0; // @[implicits.scala 55:10:@38055.4]
  assign _T_972 = _T_367 & _T_971; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:194:@38056.4]
  assign x1097_x647_D1 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@38039.4 package.scala 96:25:@38040.4]
  assign _T_973 = _T_972 & x1097_x647_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:282:@38057.4]
  assign _T_974 = _T_973 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:291:@38058.4]
  assign x653_rdcol_number = x653_rdcol_1_io_result; // @[Math.scala 154:22:@38077.4 Math.scala 155:14:@38078.4]
  assign _T_989 = $signed(x653_rdcol_number); // @[Math.scala 465:37:@38083.4]
  assign x654 = $signed(_T_989) < $signed(32'sh0); // @[Math.scala 465:44:@38085.4]
  assign x655 = x617 | x654; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 363:59:@38088.4]
  assign _T_999 = x653_rdcol_number[31]; // @[FixedPoint.scala 50:25:@38095.4]
  assign _T_1003 = _T_999 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@38097.4]
  assign _T_1004 = x653_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@38098.4]
  assign _T_1027 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@38132.4 package.scala 96:25:@38133.4]
  assign _T_1029 = io_rr ? _T_1027 : 1'h0; // @[implicits.scala 55:10:@38134.4]
  assign _T_1030 = _T_367 & _T_1029; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:194:@38135.4]
  assign x1098_x656_D1 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@38118.4 package.scala 96:25:@38119.4]
  assign _T_1031 = _T_1030 & x1098_x656_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:282:@38136.4]
  assign _T_1032 = _T_1031 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:291:@38137.4]
  assign x665_rdcol_number = x665_rdcol_1_io_result; // @[Math.scala 154:22:@38156.4 Math.scala 155:14:@38157.4]
  assign _T_1047 = $signed(x665_rdcol_number); // @[Math.scala 465:37:@38162.4]
  assign x666 = $signed(_T_1047) < $signed(32'sh0); // @[Math.scala 465:44:@38164.4]
  assign x667 = x617 | x666; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 384:59:@38167.4]
  assign _T_1057 = x665_rdcol_number[31]; // @[FixedPoint.scala 50:25:@38174.4]
  assign _T_1061 = _T_1057 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@38176.4]
  assign _T_1062 = x665_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@38177.4]
  assign _T_1085 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@38211.4 package.scala 96:25:@38212.4]
  assign _T_1087 = io_rr ? _T_1085 : 1'h0; // @[implicits.scala 55:10:@38213.4]
  assign _T_1088 = _T_367 & _T_1087; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 397:194:@38214.4]
  assign x1099_x668_D1 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@38197.4 package.scala 96:25:@38198.4]
  assign _T_1089 = _T_1088 & x1099_x668_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 397:282:@38215.4]
  assign _T_1090 = _T_1089 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 397:291:@38216.4]
  assign x1100_b535_D11_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@38232.4 package.scala 96:25:@38233.4]
  assign _T_1103 = $signed(x1100_b535_D11_number); // @[Math.scala 406:49:@38239.4]
  assign _T_1105 = $signed(_T_1103) & $signed(32'sh3); // @[Math.scala 406:56:@38241.4]
  assign _T_1106 = $signed(_T_1105); // @[Math.scala 406:56:@38242.4]
  assign x1052_number = $unsigned(_T_1106); // @[implicits.scala 133:21:@38243.4]
  assign x678 = $signed(_T_1103) < $signed(32'sh0); // @[Math.scala 465:44:@38251.4]
  assign x1101_x678_D1 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@38259.4 package.scala 96:25:@38260.4]
  assign x679 = x1101_x678_D1 | x618; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 409:25:@38263.4]
  assign _T_1130 = $signed(x1052_number); // @[Math.scala 406:49:@38272.4]
  assign _T_1132 = $signed(_T_1130) & $signed(32'sh3); // @[Math.scala 406:56:@38274.4]
  assign _T_1133 = $signed(_T_1132); // @[Math.scala 406:56:@38275.4]
  assign _T_1138 = x1052_number[31]; // @[FixedPoint.scala 50:25:@38281.4]
  assign _T_1142 = _T_1138 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@38283.4]
  assign _T_1143 = x1052_number[31:2]; // @[FixedPoint.scala 18:52:@38284.4]
  assign _T_1172 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@38336.4 package.scala 96:25:@38337.4]
  assign _T_1174 = io_rr ? _T_1172 : 1'h0; // @[implicits.scala 55:10:@38338.4]
  assign _T_1175 = _T_367 & _T_1174; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:194:@38339.4]
  assign x1103_x680_D1 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@38313.4 package.scala 96:25:@38314.4]
  assign _T_1176 = _T_1175 & x1103_x680_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:282:@38340.4]
  assign _T_1177 = _T_1176 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:291:@38341.4]
  assign x689 = x1101_x678_D1 | x629; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 438:60:@38352.4]
  assign _T_1207 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@38389.4 package.scala 96:25:@38390.4]
  assign _T_1209 = io_rr ? _T_1207 : 1'h0; // @[implicits.scala 55:10:@38391.4]
  assign _T_1210 = _T_367 & _T_1209; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:194:@38392.4]
  assign x1105_x690_D1 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@38375.4 package.scala 96:25:@38376.4]
  assign _T_1211 = _T_1210 & x1105_x690_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:282:@38393.4]
  assign _T_1212 = _T_1211 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:291:@38394.4]
  assign x696 = x1101_x678_D1 | x637; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 455:60:@38405.4]
  assign _T_1240 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@38440.4 package.scala 96:25:@38441.4]
  assign _T_1242 = io_rr ? _T_1240 : 1'h0; // @[implicits.scala 55:10:@38442.4]
  assign _T_1243 = _T_367 & _T_1242; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:194:@38443.4]
  assign x1106_x697_D1 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@38426.4 package.scala 96:25:@38427.4]
  assign _T_1244 = _T_1243 & x1106_x697_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:282:@38444.4]
  assign _T_1245 = _T_1244 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:291:@38445.4]
  assign x703 = x678 | x645; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 470:59:@38456.4]
  assign _T_1279 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@38509.4 package.scala 96:25:@38510.4]
  assign _T_1281 = io_rr ? _T_1279 : 1'h0; // @[implicits.scala 55:10:@38511.4]
  assign _T_1282 = _T_367 & _T_1281; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:194:@38512.4]
  assign x1108_x704_D2 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@38486.4 package.scala 96:25:@38487.4]
  assign _T_1283 = _T_1282 & x1108_x704_D2; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:282:@38513.4]
  assign _T_1284 = _T_1283 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:291:@38514.4]
  assign x710 = x1101_x678_D1 | x654; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 489:60:@38525.4]
  assign _T_1312 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@38560.4 package.scala 96:25:@38561.4]
  assign _T_1314 = io_rr ? _T_1312 : 1'h0; // @[implicits.scala 55:10:@38562.4]
  assign _T_1315 = _T_367 & _T_1314; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:194:@38563.4]
  assign x1110_x711_D1 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@38546.4 package.scala 96:25:@38547.4]
  assign _T_1316 = _T_1315 & x1110_x711_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:282:@38564.4]
  assign _T_1317 = _T_1316 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:291:@38565.4]
  assign x717 = x1101_x678_D1 | x666; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 504:60:@38576.4]
  assign _T_1345 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@38611.4 package.scala 96:25:@38612.4]
  assign _T_1347 = io_rr ? _T_1345 : 1'h0; // @[implicits.scala 55:10:@38613.4]
  assign _T_1348 = _T_367 & _T_1347; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:194:@38614.4]
  assign x1111_x718_D1 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@38597.4 package.scala 96:25:@38598.4]
  assign _T_1349 = _T_1348 & x1111_x718_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:282:@38615.4]
  assign _T_1350 = _T_1349 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:291:@38616.4]
  assign x724_rdrow_number = x724_rdrow_1_io_result; // @[Math.scala 154:22:@38635.4 Math.scala 155:14:@38636.4]
  assign _T_1367 = $signed(x724_rdrow_number); // @[Math.scala 406:49:@38642.4]
  assign _T_1369 = $signed(_T_1367) & $signed(32'sh3); // @[Math.scala 406:56:@38644.4]
  assign _T_1370 = $signed(_T_1369); // @[Math.scala 406:56:@38645.4]
  assign x1054_number = $unsigned(_T_1370); // @[implicits.scala 133:21:@38646.4]
  assign x726 = $signed(_T_1367) < $signed(32'sh0); // @[Math.scala 465:44:@38654.4]
  assign x727 = x726 | x618; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 525:24:@38657.4]
  assign _T_1391 = $signed(x1054_number); // @[Math.scala 406:49:@38666.4]
  assign _T_1393 = $signed(_T_1391) & $signed(32'sh3); // @[Math.scala 406:56:@38668.4]
  assign _T_1394 = $signed(_T_1393); // @[Math.scala 406:56:@38669.4]
  assign _T_1399 = x1054_number[31]; // @[FixedPoint.scala 50:25:@38675.4]
  assign _T_1403 = _T_1399 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@38677.4]
  assign _T_1404 = x1054_number[31:2]; // @[FixedPoint.scala 18:52:@38678.4]
  assign _T_1430 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@38721.4 package.scala 96:25:@38722.4]
  assign _T_1432 = io_rr ? _T_1430 : 1'h0; // @[implicits.scala 55:10:@38723.4]
  assign _T_1433 = _T_367 & _T_1432; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:194:@38724.4]
  assign x1113_x728_D1 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@38707.4 package.scala 96:25:@38708.4]
  assign _T_1434 = _T_1433 & x1113_x728_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:282:@38725.4]
  assign _T_1435 = _T_1434 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:291:@38726.4]
  assign x737 = x726 | x629; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 546:24:@38737.4]
  assign _T_1465 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@38774.4 package.scala 96:25:@38775.4]
  assign _T_1467 = io_rr ? _T_1465 : 1'h0; // @[implicits.scala 55:10:@38776.4]
  assign _T_1468 = _T_367 & _T_1467; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:194:@38777.4]
  assign x1114_x738_D1 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@38760.4 package.scala 96:25:@38761.4]
  assign _T_1469 = _T_1468 & x1114_x738_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:282:@38778.4]
  assign _T_1470 = _T_1469 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:291:@38779.4]
  assign x744 = x726 | x637; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 569:59:@38790.4]
  assign _T_1498 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@38825.4 package.scala 96:25:@38826.4]
  assign _T_1500 = io_rr ? _T_1498 : 1'h0; // @[implicits.scala 55:10:@38827.4]
  assign _T_1501 = _T_367 & _T_1500; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:194:@38828.4]
  assign x1115_x745_D1 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@38811.4 package.scala 96:25:@38812.4]
  assign _T_1502 = _T_1501 & x1115_x745_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:282:@38829.4]
  assign _T_1503 = _T_1502 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:291:@38830.4]
  assign x751 = x726 | x1095_x645_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 584:59:@38841.4]
  assign _T_1531 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@38876.4 package.scala 96:25:@38877.4]
  assign _T_1533 = io_rr ? _T_1531 : 1'h0; // @[implicits.scala 55:10:@38878.4]
  assign _T_1534 = _T_367 & _T_1533; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:194:@38879.4]
  assign x1116_x752_D1 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@38862.4 package.scala 96:25:@38863.4]
  assign _T_1535 = _T_1534 & x1116_x752_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:282:@38880.4]
  assign _T_1536 = _T_1535 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:291:@38881.4]
  assign x758 = x726 | x654; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 599:59:@38892.4]
  assign _T_1564 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@38927.4 package.scala 96:25:@38928.4]
  assign _T_1566 = io_rr ? _T_1564 : 1'h0; // @[implicits.scala 55:10:@38929.4]
  assign _T_1567 = _T_367 & _T_1566; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:194:@38930.4]
  assign x1117_x759_D1 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@38913.4 package.scala 96:25:@38914.4]
  assign _T_1568 = _T_1567 & x1117_x759_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:282:@38931.4]
  assign _T_1569 = _T_1568 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:291:@38932.4]
  assign x765 = x726 | x666; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 614:59:@38943.4]
  assign _T_1597 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@38978.4 package.scala 96:25:@38979.4]
  assign _T_1599 = io_rr ? _T_1597 : 1'h0; // @[implicits.scala 55:10:@38980.4]
  assign _T_1600 = _T_367 & _T_1599; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:194:@38981.4]
  assign x1118_x766_D1 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@38964.4 package.scala 96:25:@38965.4]
  assign _T_1601 = _T_1600 & x1118_x766_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:282:@38982.4]
  assign _T_1602 = _T_1601 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:291:@38983.4]
  assign x772_rdrow_number = x772_rdrow_1_io_result; // @[Math.scala 154:22:@39002.4 Math.scala 155:14:@39003.4]
  assign _T_1619 = $signed(x772_rdrow_number); // @[Math.scala 406:49:@39009.4]
  assign _T_1621 = $signed(_T_1619) & $signed(32'sh3); // @[Math.scala 406:56:@39011.4]
  assign _T_1622 = $signed(_T_1621); // @[Math.scala 406:56:@39012.4]
  assign x1056_number = $unsigned(_T_1622); // @[implicits.scala 133:21:@39013.4]
  assign x774 = $signed(_T_1619) < $signed(32'sh0); // @[Math.scala 465:44:@39021.4]
  assign x775 = x774 | x618; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 635:24:@39024.4]
  assign _T_1643 = $signed(x1056_number); // @[Math.scala 406:49:@39033.4]
  assign _T_1645 = $signed(_T_1643) & $signed(32'sh3); // @[Math.scala 406:56:@39035.4]
  assign _T_1646 = $signed(_T_1645); // @[Math.scala 406:56:@39036.4]
  assign _T_1651 = x1056_number[31]; // @[FixedPoint.scala 50:25:@39042.4]
  assign _T_1655 = _T_1651 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@39044.4]
  assign _T_1656 = x1056_number[31:2]; // @[FixedPoint.scala 18:52:@39045.4]
  assign _T_1682 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@39088.4 package.scala 96:25:@39089.4]
  assign _T_1684 = io_rr ? _T_1682 : 1'h0; // @[implicits.scala 55:10:@39090.4]
  assign _T_1685 = _T_367 & _T_1684; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 652:194:@39091.4]
  assign x1120_x776_D1 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@39074.4 package.scala 96:25:@39075.4]
  assign _T_1686 = _T_1685 & x1120_x776_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 652:282:@39092.4]
  assign _T_1687 = _T_1686 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 652:291:@39093.4]
  assign x785 = x774 | x629; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 656:24:@39104.4]
  assign _T_1715 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@39139.4 package.scala 96:25:@39140.4]
  assign _T_1717 = io_rr ? _T_1715 : 1'h0; // @[implicits.scala 55:10:@39141.4]
  assign _T_1718 = _T_367 & _T_1717; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:194:@39142.4]
  assign x1121_x786_D1 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@39125.4 package.scala 96:25:@39126.4]
  assign _T_1719 = _T_1718 & x1121_x786_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:282:@39143.4]
  assign _T_1720 = _T_1719 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:291:@39144.4]
  assign x792 = x774 | x637; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 671:24:@39155.4]
  assign _T_1750 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@39192.4 package.scala 96:25:@39193.4]
  assign _T_1752 = io_rr ? _T_1750 : 1'h0; // @[implicits.scala 55:10:@39194.4]
  assign _T_1753 = _T_367 & _T_1752; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:194:@39195.4]
  assign x1122_x793_D1 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@39178.4 package.scala 96:25:@39179.4]
  assign _T_1754 = _T_1753 & x1122_x793_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:282:@39196.4]
  assign _T_1755 = _T_1754 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:291:@39197.4]
  assign x799 = x774 | x1095_x645_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 694:59:@39208.4]
  assign _T_1783 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@39243.4 package.scala 96:25:@39244.4]
  assign _T_1785 = io_rr ? _T_1783 : 1'h0; // @[implicits.scala 55:10:@39245.4]
  assign _T_1786 = _T_367 & _T_1785; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:194:@39246.4]
  assign x1123_x800_D1 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@39229.4 package.scala 96:25:@39230.4]
  assign _T_1787 = _T_1786 & x1123_x800_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:282:@39247.4]
  assign _T_1788 = _T_1787 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:291:@39248.4]
  assign x806 = x774 | x654; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 709:59:@39259.4]
  assign _T_1816 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@39294.4 package.scala 96:25:@39295.4]
  assign _T_1818 = io_rr ? _T_1816 : 1'h0; // @[implicits.scala 55:10:@39296.4]
  assign _T_1819 = _T_367 & _T_1818; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:194:@39297.4]
  assign x1124_x807_D1 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@39280.4 package.scala 96:25:@39281.4]
  assign _T_1820 = _T_1819 & x1124_x807_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:282:@39298.4]
  assign _T_1821 = _T_1820 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:291:@39299.4]
  assign x813 = x774 | x666; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 724:59:@39310.4]
  assign _T_1849 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@39345.4 package.scala 96:25:@39346.4]
  assign _T_1851 = io_rr ? _T_1849 : 1'h0; // @[implicits.scala 55:10:@39347.4]
  assign _T_1852 = _T_367 & _T_1851; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 735:194:@39348.4]
  assign x1125_x814_D1 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@39331.4 package.scala 96:25:@39332.4]
  assign _T_1853 = _T_1852 & x1125_x814_D1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 735:282:@39349.4]
  assign _T_1854 = _T_1853 & x1086_b537_D13; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 735:291:@39350.4]
  assign x635_rd_0_number = x539_lb_0_io_rPort_22_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 305:29:@37879.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 309:445:@37902.4]
  assign _GEN_0 = {{1'd0}, x635_rd_0_number}; // @[Math.scala 450:32:@39362.4]
  assign _T_1860 = _GEN_0 << 1; // @[Math.scala 450:32:@39362.4]
  assign x687_rd_0_number = x539_lb_0_io_rPort_5_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 430:29:@38325.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 434:410:@38348.4]
  assign _GEN_1 = {{1'd0}, x687_rd_0_number}; // @[Math.scala 450:32:@39367.4]
  assign _T_1864 = _GEN_1 << 1; // @[Math.scala 450:32:@39367.4]
  assign x694_rd_0_number = x539_lb_0_io_rPort_9_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 447:29:@38378.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 451:410:@38401.4]
  assign _GEN_2 = {{2'd0}, x694_rd_0_number}; // @[Math.scala 450:32:@39372.4]
  assign _T_1868 = _GEN_2 << 2; // @[Math.scala 450:32:@39372.4]
  assign x701_rd_0_number = x539_lb_0_io_rPort_8_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 462:29:@38429.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 466:410:@38452.4]
  assign _GEN_3 = {{1'd0}, x701_rd_0_number}; // @[Math.scala 450:32:@39377.4]
  assign _T_1872 = _GEN_3 << 1; // @[Math.scala 450:32:@39377.4]
  assign x742_rd_0_number = x539_lb_0_io_rPort_6_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 561:29:@38763.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 565:410:@38786.4]
  assign _GEN_4 = {{1'd0}, x742_rd_0_number}; // @[Math.scala 450:32:@39382.4]
  assign _T_1876 = _GEN_4 << 1; // @[Math.scala 450:32:@39382.4]
  assign x832_sum_number = x832_sum_1_io_result; // @[Math.scala 154:22:@39471.4 Math.scala 155:14:@39472.4]
  assign _T_1912 = x832_sum_number[7:4]; // @[FixedPoint.scala 18:52:@39477.4]
  assign x834_sub_number = x834_sub_1_io_result; // @[Math.scala 195:22:@39504.4 Math.scala 196:14:@39505.4]
  assign x835 = 8'hf < x834_sub_number; // @[Math.scala 466:37:@39510.4]
  assign x833_number = RetimeWrapper_101_io_out; // @[package.scala 96:25:@39484.4 package.scala 96:25:@39485.4]
  assign x1131_x837_D6 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@39577.4 package.scala 96:25:@39578.4]
  assign x1130_x833_D6_number = RetimeWrapper_105_io_out; // @[package.scala 96:25:@39568.4 package.scala 96:25:@39569.4]
  assign x839_sum_number = x839_sum_1_io_result; // @[Math.scala 154:22:@39559.4 Math.scala 155:14:@39560.4]
  assign x840_number = x1131_x837_D6 ? x1130_x833_D6_number : x839_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 791:24:@39581.4]
  assign x643_rd_0_number = x539_lb_0_io_rPort_16_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 328:29:@37957.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 332:410:@37980.4]
  assign _GEN_5 = {{1'd0}, x643_rd_0_number}; // @[Math.scala 450:32:@39587.4]
  assign _T_1969 = _GEN_5 << 1; // @[Math.scala 450:32:@39587.4]
  assign _GEN_6 = {{1'd0}, x694_rd_0_number}; // @[Math.scala 450:32:@39592.4]
  assign _T_1973 = _GEN_6 << 1; // @[Math.scala 450:32:@39592.4]
  assign _GEN_7 = {{2'd0}, x701_rd_0_number}; // @[Math.scala 450:32:@39597.4]
  assign _T_1977 = _GEN_7 << 2; // @[Math.scala 450:32:@39597.4]
  assign x708_rd_0_number = x539_lb_0_io_rPort_23_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 481:29:@38498.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 485:410:@38521.4]
  assign _GEN_8 = {{1'd0}, x708_rd_0_number}; // @[Math.scala 450:32:@39602.4]
  assign _T_1981 = _GEN_8 << 1; // @[Math.scala 450:32:@39602.4]
  assign x749_rd_0_number = x539_lb_0_io_rPort_15_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 576:29:@38814.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 580:410:@38837.4]
  assign _GEN_9 = {{1'd0}, x749_rd_0_number}; // @[Math.scala 450:32:@39607.4]
  assign _T_1985 = _GEN_9 << 1; // @[Math.scala 450:32:@39607.4]
  assign x853_sum_number = x853_sum_1_io_result; // @[Math.scala 154:22:@39696.4 Math.scala 155:14:@39697.4]
  assign _T_2021 = x853_sum_number[7:4]; // @[FixedPoint.scala 18:52:@39702.4]
  assign x855_sub_number = x855_sub_1_io_result; // @[Math.scala 195:22:@39729.4 Math.scala 196:14:@39730.4]
  assign x856 = 8'hf < x855_sub_number; // @[Math.scala 466:37:@39735.4]
  assign x854_number = RetimeWrapper_108_io_out; // @[package.scala 96:25:@39709.4 package.scala 96:25:@39710.4]
  assign x1137_x858_D6 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@39802.4 package.scala 96:25:@39803.4]
  assign x1136_x854_D6_number = RetimeWrapper_112_io_out; // @[package.scala 96:25:@39793.4 package.scala 96:25:@39794.4]
  assign x860_sum_number = x860_sum_1_io_result; // @[Math.scala 154:22:@39784.4 Math.scala 155:14:@39785.4]
  assign x861_number = x1137_x858_D6 ? x1136_x854_D6_number : x860_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 853:24:@39806.4]
  assign x651_rd_0_number = x539_lb_0_io_rPort_2_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 351:29:@38042.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 355:410:@38065.4]
  assign _GEN_10 = {{1'd0}, x651_rd_0_number}; // @[Math.scala 450:32:@39810.4]
  assign _T_2076 = _GEN_10 << 1; // @[Math.scala 450:32:@39810.4]
  assign _GEN_11 = {{2'd0}, x708_rd_0_number}; // @[Math.scala 450:32:@39815.4]
  assign _T_2080 = _GEN_11 << 2; // @[Math.scala 450:32:@39815.4]
  assign x715_rd_0_number = x539_lb_0_io_rPort_1_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 496:29:@38549.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 500:410:@38572.4]
  assign _GEN_12 = {{1'd0}, x715_rd_0_number}; // @[Math.scala 450:32:@39820.4]
  assign _T_2084 = _GEN_12 << 1; // @[Math.scala 450:32:@39820.4]
  assign x756_rd_0_number = x539_lb_0_io_rPort_4_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 591:29:@38865.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 595:410:@38888.4]
  assign _GEN_13 = {{1'd0}, x756_rd_0_number}; // @[Math.scala 450:32:@39825.4]
  assign _T_2088 = _GEN_13 << 1; // @[Math.scala 450:32:@39825.4]
  assign x873_sum_number = x873_sum_1_io_result; // @[Math.scala 154:22:@39914.4 Math.scala 155:14:@39915.4]
  assign _T_2124 = x873_sum_number[7:4]; // @[FixedPoint.scala 18:52:@39920.4]
  assign x875_sub_number = x875_sub_1_io_result; // @[Math.scala 195:22:@39947.4 Math.scala 196:14:@39948.4]
  assign x876 = 8'hf < x875_sub_number; // @[Math.scala 466:37:@39953.4]
  assign x874_number = RetimeWrapper_115_io_out; // @[package.scala 96:25:@39927.4 package.scala 96:25:@39928.4]
  assign x1143_x878_D6 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@40022.4 package.scala 96:25:@40023.4]
  assign x1142_x874_D6_number = RetimeWrapper_119_io_out; // @[package.scala 96:25:@40013.4 package.scala 96:25:@40014.4]
  assign x880_sum_number = x880_sum_1_io_result; // @[Math.scala 154:22:@40004.4 Math.scala 155:14:@40005.4]
  assign x881_number = x1143_x878_D6 ? x1142_x874_D6_number : x880_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 913:24:@40026.4]
  assign x663_rd_0_number = x539_lb_0_io_rPort_14_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 372:29:@38121.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 376:410:@38144.4]
  assign _GEN_14 = {{1'd0}, x663_rd_0_number}; // @[Math.scala 450:32:@40030.4]
  assign _T_2181 = _GEN_14 << 1; // @[Math.scala 450:32:@40030.4]
  assign _GEN_15 = {{2'd0}, x715_rd_0_number}; // @[Math.scala 450:32:@40035.4]
  assign _T_2185 = _GEN_15 << 2; // @[Math.scala 450:32:@40035.4]
  assign x722_rd_0_number = x539_lb_0_io_rPort_12_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 511:29:@38600.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 515:410:@38623.4]
  assign _GEN_16 = {{1'd0}, x722_rd_0_number}; // @[Math.scala 450:32:@40040.4]
  assign _T_2189 = _GEN_16 << 1; // @[Math.scala 450:32:@40040.4]
  assign x763_rd_0_number = x539_lb_0_io_rPort_18_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 606:29:@38916.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 610:410:@38939.4]
  assign _GEN_17 = {{1'd0}, x763_rd_0_number}; // @[Math.scala 450:32:@40045.4]
  assign _T_2193 = _GEN_17 << 1; // @[Math.scala 450:32:@40045.4]
  assign x893_sum_number = x893_sum_1_io_result; // @[Math.scala 154:22:@40134.4 Math.scala 155:14:@40135.4]
  assign _T_2229 = x893_sum_number[7:4]; // @[FixedPoint.scala 18:52:@40140.4]
  assign x895_sub_number = x895_sub_1_io_result; // @[Math.scala 195:22:@40167.4 Math.scala 196:14:@40168.4]
  assign x896 = 8'hf < x895_sub_number; // @[Math.scala 466:37:@40173.4]
  assign x894_number = RetimeWrapper_122_io_out; // @[package.scala 96:25:@40147.4 package.scala 96:25:@40148.4]
  assign x1149_x898_D6 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@40240.4 package.scala 96:25:@40241.4]
  assign x1148_x894_D6_number = RetimeWrapper_126_io_out; // @[package.scala 96:25:@40231.4 package.scala 96:25:@40232.4]
  assign x900_sum_number = x900_sum_1_io_result; // @[Math.scala 154:22:@40222.4 Math.scala 155:14:@40223.4]
  assign x901_number = x1149_x898_D6 ? x1148_x894_D6_number : x900_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 965:24:@40244.4]
  assign x735_rd_0_number = x539_lb_0_io_rPort_21_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 538:29:@38710.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 542:410:@38733.4]
  assign _GEN_18 = {{1'd0}, x735_rd_0_number}; // @[Math.scala 450:32:@40248.4]
  assign _T_2284 = _GEN_18 << 1; // @[Math.scala 450:32:@40248.4]
  assign _GEN_19 = {{2'd0}, x742_rd_0_number}; // @[Math.scala 450:32:@40253.4]
  assign _T_2288 = _GEN_19 << 2; // @[Math.scala 450:32:@40253.4]
  assign x790_rd_0_number = x539_lb_0_io_rPort_20_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 663:29:@39128.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 667:410:@39151.4]
  assign _GEN_20 = {{1'd0}, x790_rd_0_number}; // @[Math.scala 450:32:@40258.4]
  assign _T_2292 = _GEN_20 << 1; // @[Math.scala 450:32:@40258.4]
  assign x912_sum_number = x912_sum_1_io_result; // @[Math.scala 154:22:@40347.4 Math.scala 155:14:@40348.4]
  assign _T_2328 = x912_sum_number[7:4]; // @[FixedPoint.scala 18:52:@40353.4]
  assign x914_sub_number = x914_sub_1_io_result; // @[Math.scala 195:22:@40380.4 Math.scala 196:14:@40381.4]
  assign x915 = 8'hf < x914_sub_number; // @[Math.scala 466:37:@40386.4]
  assign x913_number = RetimeWrapper_129_io_out; // @[package.scala 96:25:@40360.4 package.scala 96:25:@40361.4]
  assign x1154_x917_D6 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@40446.4 package.scala 96:25:@40447.4]
  assign x1155_x913_D6_number = RetimeWrapper_134_io_out; // @[package.scala 96:25:@40455.4 package.scala 96:25:@40456.4]
  assign x919_sum_number = x919_sum_1_io_result; // @[Math.scala 154:22:@40437.4 Math.scala 155:14:@40438.4]
  assign x920_number = x1154_x917_D6 ? x1155_x913_D6_number : x919_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1023:24:@40459.4]
  assign _GEN_21 = {{2'd0}, x749_rd_0_number}; // @[Math.scala 450:32:@40463.4]
  assign _T_2385 = _GEN_21 << 2; // @[Math.scala 450:32:@40463.4]
  assign x797_rd_0_number = x539_lb_0_io_rPort_0_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 686:29:@39181.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 690:410:@39204.4]
  assign _GEN_22 = {{1'd0}, x797_rd_0_number}; // @[Math.scala 450:32:@40468.4]
  assign _T_2389 = _GEN_22 << 1; // @[Math.scala 450:32:@40468.4]
  assign x930_sum_number = x930_sum_1_io_result; // @[Math.scala 154:22:@40557.4 Math.scala 155:14:@40558.4]
  assign _T_2425 = x930_sum_number[7:4]; // @[FixedPoint.scala 18:52:@40563.4]
  assign x932_sub_number = x932_sub_1_io_result; // @[Math.scala 195:22:@40590.4 Math.scala 196:14:@40591.4]
  assign x933 = 8'hf < x932_sub_number; // @[Math.scala 466:37:@40596.4]
  assign x931_number = RetimeWrapper_136_io_out; // @[package.scala 96:25:@40570.4 package.scala 96:25:@40571.4]
  assign x1160_x935_D6 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@40654.4 package.scala 96:25:@40655.4]
  assign x1161_x931_D6_number = RetimeWrapper_141_io_out; // @[package.scala 96:25:@40663.4 package.scala 96:25:@40664.4]
  assign x937_sum_number = x937_sum_1_io_result; // @[Math.scala 154:22:@40645.4 Math.scala 155:14:@40646.4]
  assign x938_number = x1160_x935_D6 ? x1161_x931_D6_number : x937_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1071:24:@40667.4]
  assign _GEN_23 = {{2'd0}, x756_rd_0_number}; // @[Math.scala 450:32:@40671.4]
  assign _T_2480 = _GEN_23 << 2; // @[Math.scala 450:32:@40671.4]
  assign x804_rd_0_number = x539_lb_0_io_rPort_10_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 701:29:@39232.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 705:410:@39255.4]
  assign _GEN_24 = {{1'd0}, x804_rd_0_number}; // @[Math.scala 450:32:@40676.4]
  assign _T_2484 = _GEN_24 << 1; // @[Math.scala 450:32:@40676.4]
  assign x948_sum_number = x948_sum_1_io_result; // @[Math.scala 154:22:@40765.4 Math.scala 155:14:@40766.4]
  assign _T_2520 = x948_sum_number[7:4]; // @[FixedPoint.scala 18:52:@40771.4]
  assign x950_sub_number = x950_sub_1_io_result; // @[Math.scala 195:22:@40798.4 Math.scala 196:14:@40799.4]
  assign x951 = 8'hf < x950_sub_number; // @[Math.scala 466:37:@40804.4]
  assign x949_number = RetimeWrapper_143_io_out; // @[package.scala 96:25:@40778.4 package.scala 96:25:@40779.4]
  assign x1166_x953_D6 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@40864.4 package.scala 96:25:@40865.4]
  assign x1167_x949_D6_number = RetimeWrapper_148_io_out; // @[package.scala 96:25:@40873.4 package.scala 96:25:@40874.4]
  assign x955_sum_number = x955_sum_1_io_result; // @[Math.scala 154:22:@40855.4 Math.scala 155:14:@40856.4]
  assign x956_number = x1166_x953_D6 ? x1167_x949_D6_number : x955_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1127:24:@40877.4]
  assign _GEN_25 = {{2'd0}, x763_rd_0_number}; // @[Math.scala 450:32:@40881.4]
  assign _T_2577 = _GEN_25 << 2; // @[Math.scala 450:32:@40881.4]
  assign x770_rd_0_number = x539_lb_0_io_rPort_3_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 621:29:@38967.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 625:410:@38990.4]
  assign _GEN_26 = {{1'd0}, x770_rd_0_number}; // @[Math.scala 450:32:@40886.4]
  assign _T_2581 = _GEN_26 << 1; // @[Math.scala 450:32:@40886.4]
  assign x811_rd_0_number = x539_lb_0_io_rPort_11_output_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 716:29:@39283.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 720:410:@39306.4]
  assign _GEN_27 = {{1'd0}, x811_rd_0_number}; // @[Math.scala 450:32:@40891.4]
  assign _T_2585 = _GEN_27 << 1; // @[Math.scala 450:32:@40891.4]
  assign x967_sum_number = x967_sum_1_io_result; // @[Math.scala 154:22:@40980.4 Math.scala 155:14:@40981.4]
  assign _T_2621 = x967_sum_number[7:4]; // @[FixedPoint.scala 18:52:@40986.4]
  assign x969_sub_number = x969_sub_1_io_result; // @[Math.scala 195:22:@41013.4 Math.scala 196:14:@41014.4]
  assign x970 = 8'hf < x969_sub_number; // @[Math.scala 466:37:@41019.4]
  assign x968_number = RetimeWrapper_150_io_out; // @[package.scala 96:25:@40993.4 package.scala 96:25:@40994.4]
  assign x1172_x972_D6 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@41077.4 package.scala 96:25:@41078.4]
  assign x1173_x968_D6_number = RetimeWrapper_155_io_out; // @[package.scala 96:25:@41086.4 package.scala 96:25:@41087.4]
  assign x974_sum_number = x974_sum_1_io_result; // @[Math.scala 154:22:@41068.4 Math.scala 155:14:@41069.4]
  assign x975_number = x1172_x972_D6 ? x1173_x968_D6_number : x974_sum_number; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1177:24:@41090.4]
  assign _T_2690 = {x920_number,x938_number,x956_number,x975_number}; // @[Cat.scala 30:58:@41104.4]
  assign _T_2693 = {x840_number,x861_number,x881_number,x901_number}; // @[Cat.scala 30:58:@41107.4]
  assign _T_2706 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@41143.4 package.scala 96:25:@41144.4]
  assign _T_2708 = io_rr ? _T_2706 : 1'h0; // @[implicits.scala 55:10:@41145.4]
  assign x1174_b537_D26 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@41125.4 package.scala 96:25:@41126.4]
  assign _T_2709 = _T_2708 & x1174_b537_D26; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1187:116:@41146.4]
  assign x1175_b538_D26 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@41134.4 package.scala 96:25:@41135.4]
  assign _T_2710 = _T_2709 & x1175_b538_D26; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1187:123:@41147.4]
  assign x1061_x1048_D8_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@37077.4 package.scala 96:25:@37078.4]
  assign x1063_x553_sum_D7_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@37095.4 package.scala 96:25:@37096.4]
  assign x1065_x563_sum_D6_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@37171.4 package.scala 96:25:@37172.4]
  assign x1068_x572_sum_D6_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@37256.4 package.scala 96:25:@37257.4]
  assign x1070_x581_sum_D6_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@37332.4 package.scala 96:25:@37333.4]
  assign x1072_x1049_D7_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@37468.4 package.scala 96:25:@37469.4]
  assign x1073_x595_sum_D6_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@37477.4 package.scala 96:25:@37478.4]
  assign x1075_x601_sum_D6_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@37532.4 package.scala 96:25:@37533.4]
  assign x1077_x606_sum_D6_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@37587.4 package.scala 96:25:@37588.4]
  assign x1080_x611_sum_D6_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@37651.4 package.scala 96:25:@37652.4]
  assign x623_sum_number = x623_sum_1_io_result; // @[Math.scala 154:22:@37764.4 Math.scala 155:14:@37765.4]
  assign x1085_x1051_D1_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@37782.4 package.scala 96:25:@37783.4]
  assign x632_sum_number = x632_sum_1_io_result; // @[Math.scala 154:22:@37867.4 Math.scala 155:14:@37868.4]
  assign x640_sum_number = x640_sum_1_io_result; // @[Math.scala 154:22:@37945.4 Math.scala 155:14:@37946.4]
  assign x648_sum_number = x648_sum_1_io_result; // @[Math.scala 154:22:@38030.4 Math.scala 155:14:@38031.4]
  assign x659_sum_number = x659_sum_1_io_result; // @[Math.scala 154:22:@38109.4 Math.scala 155:14:@38110.4]
  assign x671_sum_number = x671_sum_1_io_result; // @[Math.scala 154:22:@38188.4 Math.scala 155:14:@38189.4]
  assign x683_sum_number = x683_sum_1_io_result; // @[Math.scala 154:22:@38304.4 Math.scala 155:14:@38305.4]
  assign x1104_x1053_D2_number = RetimeWrapper_60_io_out; // @[package.scala 96:25:@38322.4 package.scala 96:25:@38323.4]
  assign x691_sum_number = x691_sum_1_io_result; // @[Math.scala 154:22:@38366.4 Math.scala 155:14:@38367.4]
  assign x698_sum_number = x698_sum_1_io_result; // @[Math.scala 154:22:@38417.4 Math.scala 155:14:@38418.4]
  assign x1109_x705_sum_D1_number = RetimeWrapper_68_io_out; // @[package.scala 96:25:@38495.4 package.scala 96:25:@38496.4]
  assign x712_sum_number = x712_sum_1_io_result; // @[Math.scala 154:22:@38537.4 Math.scala 155:14:@38538.4]
  assign x719_sum_number = x719_sum_1_io_result; // @[Math.scala 154:22:@38588.4 Math.scala 155:14:@38589.4]
  assign x731_sum_number = x731_sum_1_io_result; // @[Math.scala 154:22:@38689.4 Math.scala 155:14:@38690.4]
  assign x1112_x1055_D1_number = RetimeWrapper_74_io_out; // @[package.scala 96:25:@38698.4 package.scala 96:25:@38699.4]
  assign x739_sum_number = x739_sum_1_io_result; // @[Math.scala 154:22:@38751.4 Math.scala 155:14:@38752.4]
  assign x746_sum_number = x746_sum_1_io_result; // @[Math.scala 154:22:@38802.4 Math.scala 155:14:@38803.4]
  assign x753_sum_number = x753_sum_1_io_result; // @[Math.scala 154:22:@38853.4 Math.scala 155:14:@38854.4]
  assign x760_sum_number = x760_sum_1_io_result; // @[Math.scala 154:22:@38904.4 Math.scala 155:14:@38905.4]
  assign x767_sum_number = x767_sum_1_io_result; // @[Math.scala 154:22:@38955.4 Math.scala 155:14:@38956.4]
  assign x779_sum_number = x779_sum_1_io_result; // @[Math.scala 154:22:@39056.4 Math.scala 155:14:@39057.4]
  assign x1119_x1057_D1_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@39065.4 package.scala 96:25:@39066.4]
  assign x787_sum_number = x787_sum_1_io_result; // @[Math.scala 154:22:@39116.4 Math.scala 155:14:@39117.4]
  assign x794_sum_number = x794_sum_1_io_result; // @[Math.scala 154:22:@39169.4 Math.scala 155:14:@39170.4]
  assign x801_sum_number = x801_sum_1_io_result; // @[Math.scala 154:22:@39220.4 Math.scala 155:14:@39221.4]
  assign x808_sum_number = x808_sum_1_io_result; // @[Math.scala 154:22:@39271.4 Math.scala 155:14:@39272.4]
  assign x815_sum_number = x815_sum_1_io_result; // @[Math.scala 154:22:@39322.4 Math.scala 155:14:@39323.4]
  assign io_in_x527_TVALID = _T_2710 & io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1187:22:@41149.4]
  assign io_in_x527_TDATA = {{192'd0}, RetimeWrapper_156_io_out}; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1188:24:@41150.4]
  assign io_in_x526_TREADY = _T_212 & _T_214; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 68:22:@36926.4 sm_x980_inr_Foreach_SAMPLER_BOX.scala 70:22:@36934.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@36691.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@36703.4]
  assign x539_lb_0_clock = clock; // @[:@36711.4]
  assign x539_lb_0_reset = reset; // @[:@36712.4]
  assign x539_lb_0_io_rPort_23_banks_0 = x1104_x1053_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@38516.4]
  assign x539_lb_0_io_rPort_23_ofs_0 = x1109_x705_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@38518.4]
  assign x539_lb_0_io_rPort_23_en_0 = _T_1284 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38520.4]
  assign x539_lb_0_io_rPort_23_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38519.4]
  assign x539_lb_0_io_rPort_22_banks_0 = x1085_x1051_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@37897.4]
  assign x539_lb_0_io_rPort_22_ofs_0 = x632_sum_number[0]; // @[MemInterfaceType.scala 107:54:@37899.4]
  assign x539_lb_0_io_rPort_22_en_0 = _T_875 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@37901.4]
  assign x539_lb_0_io_rPort_22_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@37900.4]
  assign x539_lb_0_io_rPort_21_banks_0 = x1112_x1055_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38728.4]
  assign x539_lb_0_io_rPort_21_ofs_0 = x731_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38730.4]
  assign x539_lb_0_io_rPort_21_en_0 = _T_1435 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38732.4]
  assign x539_lb_0_io_rPort_21_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38731.4]
  assign x539_lb_0_io_rPort_20_banks_0 = x1119_x1057_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@39146.4]
  assign x539_lb_0_io_rPort_20_ofs_0 = x787_sum_number[0]; // @[MemInterfaceType.scala 107:54:@39148.4]
  assign x539_lb_0_io_rPort_20_en_0 = _T_1720 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@39150.4]
  assign x539_lb_0_io_rPort_20_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39149.4]
  assign x539_lb_0_io_rPort_19_banks_0 = x1119_x1057_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@39352.4]
  assign x539_lb_0_io_rPort_19_ofs_0 = x815_sum_number[0]; // @[MemInterfaceType.scala 107:54:@39354.4]
  assign x539_lb_0_io_rPort_19_en_0 = _T_1854 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@39356.4]
  assign x539_lb_0_io_rPort_19_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39355.4]
  assign x539_lb_0_io_rPort_18_banks_0 = x1112_x1055_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38934.4]
  assign x539_lb_0_io_rPort_18_ofs_0 = x760_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38936.4]
  assign x539_lb_0_io_rPort_18_en_0 = _T_1569 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38938.4]
  assign x539_lb_0_io_rPort_18_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38937.4]
  assign x539_lb_0_io_rPort_17_banks_0 = x1085_x1051_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@37821.4]
  assign x539_lb_0_io_rPort_17_ofs_0 = x623_sum_number[0]; // @[MemInterfaceType.scala 107:54:@37823.4]
  assign x539_lb_0_io_rPort_17_en_0 = _T_828 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@37825.4]
  assign x539_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@37824.4]
  assign x539_lb_0_io_rPort_16_banks_0 = x1085_x1051_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@37975.4]
  assign x539_lb_0_io_rPort_16_ofs_0 = x640_sum_number[0]; // @[MemInterfaceType.scala 107:54:@37977.4]
  assign x539_lb_0_io_rPort_16_en_0 = _T_924 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@37979.4]
  assign x539_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@37978.4]
  assign x539_lb_0_io_rPort_15_banks_0 = x1112_x1055_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38832.4]
  assign x539_lb_0_io_rPort_15_ofs_0 = x746_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38834.4]
  assign x539_lb_0_io_rPort_15_en_0 = _T_1503 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38836.4]
  assign x539_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38835.4]
  assign x539_lb_0_io_rPort_14_banks_0 = x1085_x1051_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38139.4]
  assign x539_lb_0_io_rPort_14_ofs_0 = x659_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38141.4]
  assign x539_lb_0_io_rPort_14_en_0 = _T_1032 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38143.4]
  assign x539_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38142.4]
  assign x539_lb_0_io_rPort_13_banks_0 = x1085_x1051_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38218.4]
  assign x539_lb_0_io_rPort_13_ofs_0 = x671_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38220.4]
  assign x539_lb_0_io_rPort_13_en_0 = _T_1090 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38222.4]
  assign x539_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38221.4]
  assign x539_lb_0_io_rPort_12_banks_0 = x1104_x1053_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@38618.4]
  assign x539_lb_0_io_rPort_12_ofs_0 = x719_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38620.4]
  assign x539_lb_0_io_rPort_12_en_0 = _T_1350 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38622.4]
  assign x539_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38621.4]
  assign x539_lb_0_io_rPort_11_banks_0 = x1119_x1057_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@39301.4]
  assign x539_lb_0_io_rPort_11_ofs_0 = x808_sum_number[0]; // @[MemInterfaceType.scala 107:54:@39303.4]
  assign x539_lb_0_io_rPort_11_en_0 = _T_1821 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@39305.4]
  assign x539_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39304.4]
  assign x539_lb_0_io_rPort_10_banks_0 = x1119_x1057_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@39250.4]
  assign x539_lb_0_io_rPort_10_ofs_0 = x801_sum_number[0]; // @[MemInterfaceType.scala 107:54:@39252.4]
  assign x539_lb_0_io_rPort_10_en_0 = _T_1788 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@39254.4]
  assign x539_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39253.4]
  assign x539_lb_0_io_rPort_9_banks_0 = x1104_x1053_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@38396.4]
  assign x539_lb_0_io_rPort_9_ofs_0 = x691_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38398.4]
  assign x539_lb_0_io_rPort_9_en_0 = _T_1212 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38400.4]
  assign x539_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38399.4]
  assign x539_lb_0_io_rPort_8_banks_0 = x1104_x1053_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@38447.4]
  assign x539_lb_0_io_rPort_8_ofs_0 = x698_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38449.4]
  assign x539_lb_0_io_rPort_8_en_0 = _T_1245 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38451.4]
  assign x539_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38450.4]
  assign x539_lb_0_io_rPort_7_banks_0 = x1119_x1057_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@39095.4]
  assign x539_lb_0_io_rPort_7_ofs_0 = x779_sum_number[0]; // @[MemInterfaceType.scala 107:54:@39097.4]
  assign x539_lb_0_io_rPort_7_en_0 = _T_1687 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@39099.4]
  assign x539_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39098.4]
  assign x539_lb_0_io_rPort_6_banks_0 = x1112_x1055_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38781.4]
  assign x539_lb_0_io_rPort_6_ofs_0 = x739_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38783.4]
  assign x539_lb_0_io_rPort_6_en_0 = _T_1470 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38785.4]
  assign x539_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38784.4]
  assign x539_lb_0_io_rPort_5_banks_0 = x1104_x1053_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@38343.4]
  assign x539_lb_0_io_rPort_5_ofs_0 = x683_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38345.4]
  assign x539_lb_0_io_rPort_5_en_0 = _T_1177 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38347.4]
  assign x539_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38346.4]
  assign x539_lb_0_io_rPort_4_banks_0 = x1112_x1055_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38883.4]
  assign x539_lb_0_io_rPort_4_ofs_0 = x753_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38885.4]
  assign x539_lb_0_io_rPort_4_en_0 = _T_1536 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38887.4]
  assign x539_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38886.4]
  assign x539_lb_0_io_rPort_3_banks_0 = x1112_x1055_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38985.4]
  assign x539_lb_0_io_rPort_3_ofs_0 = x767_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38987.4]
  assign x539_lb_0_io_rPort_3_en_0 = _T_1602 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38989.4]
  assign x539_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38988.4]
  assign x539_lb_0_io_rPort_2_banks_0 = x1085_x1051_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@38060.4]
  assign x539_lb_0_io_rPort_2_ofs_0 = x648_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38062.4]
  assign x539_lb_0_io_rPort_2_en_0 = _T_974 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38064.4]
  assign x539_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38063.4]
  assign x539_lb_0_io_rPort_1_banks_0 = x1104_x1053_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@38567.4]
  assign x539_lb_0_io_rPort_1_ofs_0 = x712_sum_number[0]; // @[MemInterfaceType.scala 107:54:@38569.4]
  assign x539_lb_0_io_rPort_1_en_0 = _T_1317 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@38571.4]
  assign x539_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38570.4]
  assign x539_lb_0_io_rPort_0_banks_0 = x1119_x1057_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@39199.4]
  assign x539_lb_0_io_rPort_0_ofs_0 = x794_sum_number[0]; // @[MemInterfaceType.scala 107:54:@39201.4]
  assign x539_lb_0_io_rPort_0_en_0 = _T_1755 & x1084_b538_D13; // @[MemInterfaceType.scala 110:79:@39203.4]
  assign x539_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@39202.4]
  assign x539_lb_0_io_wPort_7_banks_0 = x1061_x1048_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@37278.4]
  assign x539_lb_0_io_wPort_7_ofs_0 = x1068_x572_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37280.4]
  assign x539_lb_0_io_wPort_7_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@37281.4]
  assign x539_lb_0_io_wPort_7_en_0 = _T_471 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37283.4]
  assign x539_lb_0_io_wPort_6_banks_0 = x1061_x1048_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@37354.4]
  assign x539_lb_0_io_wPort_6_ofs_0 = x1070_x581_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37356.4]
  assign x539_lb_0_io_wPort_6_data_0 = RetimeWrapper_14_io_out; // @[MemInterfaceType.scala 90:56:@37357.4]
  assign x539_lb_0_io_wPort_6_en_0 = _T_516 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37359.4]
  assign x539_lb_0_io_wPort_5_banks_0 = x1072_x1049_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@37618.4]
  assign x539_lb_0_io_wPort_5_ofs_0 = x1077_x606_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37620.4]
  assign x539_lb_0_io_wPort_5_data_0 = RetimeWrapper_26_io_out; // @[MemInterfaceType.scala 90:56:@37621.4]
  assign x539_lb_0_io_wPort_5_en_0 = _T_700 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37623.4]
  assign x539_lb_0_io_wPort_4_banks_0 = x1072_x1049_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@37508.4]
  assign x539_lb_0_io_wPort_4_ofs_0 = x1073_x595_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37510.4]
  assign x539_lb_0_io_wPort_4_data_0 = RetimeWrapper_20_io_out; // @[MemInterfaceType.scala 90:56:@37511.4]
  assign x539_lb_0_io_wPort_4_en_0 = _T_644 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37513.4]
  assign x539_lb_0_io_wPort_3_banks_0 = x1061_x1048_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@37202.4]
  assign x539_lb_0_io_wPort_3_ofs_0 = x1065_x563_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37204.4]
  assign x539_lb_0_io_wPort_3_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@37205.4]
  assign x539_lb_0_io_wPort_3_en_0 = _T_426 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37207.4]
  assign x539_lb_0_io_wPort_2_banks_0 = x1072_x1049_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@37563.4]
  assign x539_lb_0_io_wPort_2_ofs_0 = x1075_x601_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37565.4]
  assign x539_lb_0_io_wPort_2_data_0 = RetimeWrapper_23_io_out; // @[MemInterfaceType.scala 90:56:@37566.4]
  assign x539_lb_0_io_wPort_2_en_0 = _T_672 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37568.4]
  assign x539_lb_0_io_wPort_1_banks_0 = x1061_x1048_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@37117.4]
  assign x539_lb_0_io_wPort_1_ofs_0 = x1063_x553_sum_D7_number[0]; // @[MemInterfaceType.scala 89:54:@37119.4]
  assign x539_lb_0_io_wPort_1_data_0 = RetimeWrapper_4_io_out; // @[MemInterfaceType.scala 90:56:@37120.4]
  assign x539_lb_0_io_wPort_1_en_0 = _T_378 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37122.4]
  assign x539_lb_0_io_wPort_0_banks_0 = x1072_x1049_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@37673.4]
  assign x539_lb_0_io_wPort_0_ofs_0 = x1080_x611_sum_D6_number[0]; // @[MemInterfaceType.scala 89:54:@37675.4]
  assign x539_lb_0_io_wPort_0_data_0 = RetimeWrapper_28_io_out; // @[MemInterfaceType.scala 90:56:@37676.4]
  assign x539_lb_0_io_wPort_0_en_0 = _T_728 & x1059_b538_D8; // @[MemInterfaceType.scala 93:57:@37678.4]
  assign RetimeWrapper_clock = clock; // @[:@36937.4]
  assign RetimeWrapper_reset = reset; // @[:@36938.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36940.4]
  assign RetimeWrapper_io_in = io_in_x526_TDATA[63:0]; // @[package.scala 94:16:@36939.4]
  assign x553_sum_1_clock = clock; // @[:@37045.4]
  assign x553_sum_1_reset = reset; // @[:@37046.4]
  assign x553_sum_1_io_a = {_T_331,_T_332}; // @[Math.scala 151:17:@37047.4]
  assign x553_sum_1_io_b = {_T_341,_T_342}; // @[Math.scala 152:17:@37048.4]
  assign x553_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37049.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37055.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37056.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37058.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@37057.4]
  assign RetimeWrapper_2_clock = clock; // @[:@37064.4]
  assign RetimeWrapper_2_reset = reset; // @[:@37065.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37067.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@37066.4]
  assign RetimeWrapper_3_clock = clock; // @[:@37073.4]
  assign RetimeWrapper_3_reset = reset; // @[:@37074.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37076.4]
  assign RetimeWrapper_3_io_in = $unsigned(_T_322); // @[package.scala 94:16:@37075.4]
  assign RetimeWrapper_4_clock = clock; // @[:@37082.4]
  assign RetimeWrapper_4_reset = reset; // @[:@37083.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37085.4]
  assign RetimeWrapper_4_io_in = x1058_x540_D1_0_number[7:0]; // @[package.scala 94:16:@37084.4]
  assign RetimeWrapper_5_clock = clock; // @[:@37091.4]
  assign RetimeWrapper_5_reset = reset; // @[:@37092.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37094.4]
  assign RetimeWrapper_5_io_in = x553_sum_1_io_result; // @[package.scala 94:16:@37093.4]
  assign RetimeWrapper_6_clock = clock; // @[:@37104.4]
  assign RetimeWrapper_6_reset = reset; // @[:@37105.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37107.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37106.4]
  assign x559_rdcol_1_clock = clock; // @[:@37127.4]
  assign x559_rdcol_1_reset = reset; // @[:@37128.4]
  assign x559_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@37129.4]
  assign x559_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@37130.4]
  assign x559_rdcol_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37131.4]
  assign RetimeWrapper_7_clock = clock; // @[:@37148.4]
  assign RetimeWrapper_7_reset = reset; // @[:@37149.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37151.4]
  assign RetimeWrapper_7_io_in = {_T_331,_T_332}; // @[package.scala 94:16:@37150.4]
  assign x563_sum_1_clock = clock; // @[:@37157.4]
  assign x563_sum_1_reset = reset; // @[:@37158.4]
  assign x563_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@37159.4]
  assign x563_sum_1_io_b = {_T_395,_T_396}; // @[Math.scala 152:17:@37160.4]
  assign x563_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37161.4]
  assign RetimeWrapper_8_clock = clock; // @[:@37167.4]
  assign RetimeWrapper_8_reset = reset; // @[:@37168.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37170.4]
  assign RetimeWrapper_8_io_in = x563_sum_1_io_result; // @[package.scala 94:16:@37169.4]
  assign RetimeWrapper_9_clock = clock; // @[:@37176.4]
  assign RetimeWrapper_9_reset = reset; // @[:@37177.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37179.4]
  assign RetimeWrapper_9_io_in = x1058_x540_D1_0_number[15:8]; // @[package.scala 94:16:@37178.4]
  assign RetimeWrapper_10_clock = clock; // @[:@37189.4]
  assign RetimeWrapper_10_reset = reset; // @[:@37190.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37192.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37191.4]
  assign x568_rdcol_1_clock = clock; // @[:@37212.4]
  assign x568_rdcol_1_reset = reset; // @[:@37213.4]
  assign x568_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@37214.4]
  assign x568_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@37215.4]
  assign x568_rdcol_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37216.4]
  assign x572_sum_1_clock = clock; // @[:@37233.4]
  assign x572_sum_1_reset = reset; // @[:@37234.4]
  assign x572_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@37235.4]
  assign x572_sum_1_io_b = {_T_443,_T_444}; // @[Math.scala 152:17:@37236.4]
  assign x572_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37237.4]
  assign RetimeWrapper_11_clock = clock; // @[:@37243.4]
  assign RetimeWrapper_11_reset = reset; // @[:@37244.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37246.4]
  assign RetimeWrapper_11_io_in = x1058_x540_D1_0_number[23:16]; // @[package.scala 94:16:@37245.4]
  assign RetimeWrapper_12_clock = clock; // @[:@37252.4]
  assign RetimeWrapper_12_reset = reset; // @[:@37253.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37255.4]
  assign RetimeWrapper_12_io_in = x572_sum_1_io_result; // @[package.scala 94:16:@37254.4]
  assign RetimeWrapper_13_clock = clock; // @[:@37265.4]
  assign RetimeWrapper_13_reset = reset; // @[:@37266.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37268.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37267.4]
  assign x577_rdcol_1_clock = clock; // @[:@37288.4]
  assign x577_rdcol_1_reset = reset; // @[:@37289.4]
  assign x577_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@37290.4]
  assign x577_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@37291.4]
  assign x577_rdcol_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37292.4]
  assign x581_sum_1_clock = clock; // @[:@37309.4]
  assign x581_sum_1_reset = reset; // @[:@37310.4]
  assign x581_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@37311.4]
  assign x581_sum_1_io_b = {_T_488,_T_489}; // @[Math.scala 152:17:@37312.4]
  assign x581_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37313.4]
  assign RetimeWrapper_14_clock = clock; // @[:@37319.4]
  assign RetimeWrapper_14_reset = reset; // @[:@37320.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37322.4]
  assign RetimeWrapper_14_io_in = x1058_x540_D1_0_number[31:24]; // @[package.scala 94:16:@37321.4]
  assign RetimeWrapper_15_clock = clock; // @[:@37328.4]
  assign RetimeWrapper_15_reset = reset; // @[:@37329.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37331.4]
  assign RetimeWrapper_15_io_in = x581_sum_1_io_result; // @[package.scala 94:16:@37330.4]
  assign RetimeWrapper_16_clock = clock; // @[:@37341.4]
  assign RetimeWrapper_16_reset = reset; // @[:@37342.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37344.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37343.4]
  assign x586_rdrow_1_clock = clock; // @[:@37364.4]
  assign x586_rdrow_1_reset = reset; // @[:@37365.4]
  assign x586_rdrow_1_io_a = __io_result; // @[Math.scala 151:17:@37366.4]
  assign x586_rdrow_1_io_b = 32'h1; // @[Math.scala 152:17:@37367.4]
  assign x586_rdrow_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37368.4]
  assign RetimeWrapper_17_clock = clock; // @[:@37445.4]
  assign RetimeWrapper_17_reset = reset; // @[:@37446.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37448.4]
  assign RetimeWrapper_17_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@37447.4]
  assign x595_sum_1_clock = clock; // @[:@37454.4]
  assign x595_sum_1_reset = reset; // @[:@37455.4]
  assign x595_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@37456.4]
  assign x595_sum_1_io_b = RetimeWrapper_17_io_out; // @[Math.scala 152:17:@37457.4]
  assign x595_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37458.4]
  assign RetimeWrapper_18_clock = clock; // @[:@37464.4]
  assign RetimeWrapper_18_reset = reset; // @[:@37465.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37467.4]
  assign RetimeWrapper_18_io_in = $unsigned(_T_601); // @[package.scala 94:16:@37466.4]
  assign RetimeWrapper_19_clock = clock; // @[:@37473.4]
  assign RetimeWrapper_19_reset = reset; // @[:@37474.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37476.4]
  assign RetimeWrapper_19_io_in = x595_sum_1_io_result; // @[package.scala 94:16:@37475.4]
  assign RetimeWrapper_20_clock = clock; // @[:@37482.4]
  assign RetimeWrapper_20_reset = reset; // @[:@37483.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37485.4]
  assign RetimeWrapper_20_io_in = x1058_x540_D1_0_number[39:32]; // @[package.scala 94:16:@37484.4]
  assign RetimeWrapper_21_clock = clock; // @[:@37495.4]
  assign RetimeWrapper_21_reset = reset; // @[:@37496.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37498.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37497.4]
  assign x601_sum_1_clock = clock; // @[:@37518.4]
  assign x601_sum_1_reset = reset; // @[:@37519.4]
  assign x601_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@37520.4]
  assign x601_sum_1_io_b = {_T_395,_T_396}; // @[Math.scala 152:17:@37521.4]
  assign x601_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37522.4]
  assign RetimeWrapper_22_clock = clock; // @[:@37528.4]
  assign RetimeWrapper_22_reset = reset; // @[:@37529.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37531.4]
  assign RetimeWrapper_22_io_in = x601_sum_1_io_result; // @[package.scala 94:16:@37530.4]
  assign RetimeWrapper_23_clock = clock; // @[:@37537.4]
  assign RetimeWrapper_23_reset = reset; // @[:@37538.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37540.4]
  assign RetimeWrapper_23_io_in = x1058_x540_D1_0_number[47:40]; // @[package.scala 94:16:@37539.4]
  assign RetimeWrapper_24_clock = clock; // @[:@37550.4]
  assign RetimeWrapper_24_reset = reset; // @[:@37551.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37553.4]
  assign RetimeWrapper_24_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37552.4]
  assign x606_sum_1_clock = clock; // @[:@37573.4]
  assign x606_sum_1_reset = reset; // @[:@37574.4]
  assign x606_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@37575.4]
  assign x606_sum_1_io_b = {_T_443,_T_444}; // @[Math.scala 152:17:@37576.4]
  assign x606_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37577.4]
  assign RetimeWrapper_25_clock = clock; // @[:@37583.4]
  assign RetimeWrapper_25_reset = reset; // @[:@37584.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37586.4]
  assign RetimeWrapper_25_io_in = x606_sum_1_io_result; // @[package.scala 94:16:@37585.4]
  assign RetimeWrapper_26_clock = clock; // @[:@37592.4]
  assign RetimeWrapper_26_reset = reset; // @[:@37593.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37595.4]
  assign RetimeWrapper_26_io_in = x1058_x540_D1_0_number[55:48]; // @[package.scala 94:16:@37594.4]
  assign RetimeWrapper_27_clock = clock; // @[:@37605.4]
  assign RetimeWrapper_27_reset = reset; // @[:@37606.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37608.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37607.4]
  assign x611_sum_1_clock = clock; // @[:@37628.4]
  assign x611_sum_1_reset = reset; // @[:@37629.4]
  assign x611_sum_1_io_a = {_T_610,_T_611}; // @[Math.scala 151:17:@37630.4]
  assign x611_sum_1_io_b = {_T_488,_T_489}; // @[Math.scala 152:17:@37631.4]
  assign x611_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37632.4]
  assign RetimeWrapper_28_clock = clock; // @[:@37638.4]
  assign RetimeWrapper_28_reset = reset; // @[:@37639.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37641.4]
  assign RetimeWrapper_28_io_in = x1058_x540_D1_0_number[63:56]; // @[package.scala 94:16:@37640.4]
  assign RetimeWrapper_29_clock = clock; // @[:@37647.4]
  assign RetimeWrapper_29_reset = reset; // @[:@37648.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37650.4]
  assign RetimeWrapper_29_io_in = x611_sum_1_io_result; // @[package.scala 94:16:@37649.4]
  assign RetimeWrapper_30_clock = clock; // @[:@37660.4]
  assign RetimeWrapper_30_reset = reset; // @[:@37661.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37663.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37662.4]
  assign RetimeWrapper_31_clock = clock; // @[:@37681.4]
  assign RetimeWrapper_31_reset = reset; // @[:@37682.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37684.4]
  assign RetimeWrapper_31_io_in = x586_rdrow_1_io_result; // @[package.scala 94:16:@37683.4]
  assign RetimeWrapper_32_clock = clock; // @[:@37708.4]
  assign RetimeWrapper_32_reset = reset; // @[:@37709.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37711.4]
  assign RetimeWrapper_32_io_in = x577_rdcol_1_io_result; // @[package.scala 94:16:@37710.4]
  assign RetimeWrapper_33_clock = clock; // @[:@37750.4]
  assign RetimeWrapper_33_reset = reset; // @[:@37751.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37753.4]
  assign RetimeWrapper_33_io_in = {_T_488,_T_489}; // @[package.scala 94:16:@37752.4]
  assign x623_sum_1_clock = clock; // @[:@37759.4]
  assign x623_sum_1_reset = reset; // @[:@37760.4]
  assign x623_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@37761.4]
  assign x623_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@37762.4]
  assign x623_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37763.4]
  assign RetimeWrapper_34_clock = clock; // @[:@37769.4]
  assign RetimeWrapper_34_reset = reset; // @[:@37770.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37772.4]
  assign RetimeWrapper_34_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@37771.4]
  assign RetimeWrapper_35_clock = clock; // @[:@37778.4]
  assign RetimeWrapper_35_reset = reset; // @[:@37779.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37781.4]
  assign RetimeWrapper_35_io_in = $unsigned(_T_778); // @[package.scala 94:16:@37780.4]
  assign RetimeWrapper_36_clock = clock; // @[:@37787.4]
  assign RetimeWrapper_36_reset = reset; // @[:@37788.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37790.4]
  assign RetimeWrapper_36_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@37789.4]
  assign RetimeWrapper_37_clock = clock; // @[:@37796.4]
  assign RetimeWrapper_37_reset = reset; // @[:@37797.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37799.4]
  assign RetimeWrapper_37_io_in = ~ x619; // @[package.scala 94:16:@37798.4]
  assign RetimeWrapper_38_clock = clock; // @[:@37810.4]
  assign RetimeWrapper_38_reset = reset; // @[:@37811.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37813.4]
  assign RetimeWrapper_38_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37812.4]
  assign RetimeWrapper_39_clock = clock; // @[:@37831.4]
  assign RetimeWrapper_39_reset = reset; // @[:@37832.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37834.4]
  assign RetimeWrapper_39_io_in = x568_rdcol_1_io_result; // @[package.scala 94:16:@37833.4]
  assign RetimeWrapper_40_clock = clock; // @[:@37853.4]
  assign RetimeWrapper_40_reset = reset; // @[:@37854.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37856.4]
  assign RetimeWrapper_40_io_in = {_T_443,_T_444}; // @[package.scala 94:16:@37855.4]
  assign x632_sum_1_clock = clock; // @[:@37862.4]
  assign x632_sum_1_reset = reset; // @[:@37863.4]
  assign x632_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@37864.4]
  assign x632_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@37865.4]
  assign x632_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37866.4]
  assign RetimeWrapper_41_clock = clock; // @[:@37872.4]
  assign RetimeWrapper_41_reset = reset; // @[:@37873.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37875.4]
  assign RetimeWrapper_41_io_in = ~ x630; // @[package.scala 94:16:@37874.4]
  assign RetimeWrapper_42_clock = clock; // @[:@37886.4]
  assign RetimeWrapper_42_reset = reset; // @[:@37887.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37889.4]
  assign RetimeWrapper_42_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37888.4]
  assign RetimeWrapper_43_clock = clock; // @[:@37907.4]
  assign RetimeWrapper_43_reset = reset; // @[:@37908.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37910.4]
  assign RetimeWrapper_43_io_in = x559_rdcol_1_io_result; // @[package.scala 94:16:@37909.4]
  assign RetimeWrapper_44_clock = clock; // @[:@37931.4]
  assign RetimeWrapper_44_reset = reset; // @[:@37932.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37934.4]
  assign RetimeWrapper_44_io_in = {_T_395,_T_396}; // @[package.scala 94:16:@37933.4]
  assign x640_sum_1_clock = clock; // @[:@37940.4]
  assign x640_sum_1_reset = reset; // @[:@37941.4]
  assign x640_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@37942.4]
  assign x640_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@37943.4]
  assign x640_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@37944.4]
  assign RetimeWrapper_45_clock = clock; // @[:@37950.4]
  assign RetimeWrapper_45_reset = reset; // @[:@37951.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37953.4]
  assign RetimeWrapper_45_io_in = ~ x638; // @[package.scala 94:16:@37952.4]
  assign RetimeWrapper_46_clock = clock; // @[:@37964.4]
  assign RetimeWrapper_46_reset = reset; // @[:@37965.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37967.4]
  assign RetimeWrapper_46_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@37966.4]
  assign RetimeWrapper_47_clock = clock; // @[:@37985.4]
  assign RetimeWrapper_47_reset = reset; // @[:@37986.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@37988.4]
  assign RetimeWrapper_47_io_in = __1_io_result; // @[package.scala 94:16:@37987.4]
  assign RetimeWrapper_48_clock = clock; // @[:@38001.4]
  assign RetimeWrapper_48_reset = reset; // @[:@38002.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38004.4]
  assign RetimeWrapper_48_io_in = $signed(_T_935) < $signed(32'sh0); // @[package.scala 94:16:@38003.4]
  assign RetimeWrapper_49_clock = clock; // @[:@38016.4]
  assign RetimeWrapper_49_reset = reset; // @[:@38017.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38019.4]
  assign RetimeWrapper_49_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@38018.4]
  assign x648_sum_1_clock = clock; // @[:@38025.4]
  assign x648_sum_1_reset = reset; // @[:@38026.4]
  assign x648_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@38027.4]
  assign x648_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@38028.4]
  assign x648_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38029.4]
  assign RetimeWrapper_50_clock = clock; // @[:@38035.4]
  assign RetimeWrapper_50_reset = reset; // @[:@38036.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38038.4]
  assign RetimeWrapper_50_io_in = ~ x646; // @[package.scala 94:16:@38037.4]
  assign RetimeWrapper_51_clock = clock; // @[:@38049.4]
  assign RetimeWrapper_51_reset = reset; // @[:@38050.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38052.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38051.4]
  assign x653_rdcol_1_clock = clock; // @[:@38072.4]
  assign x653_rdcol_1_reset = reset; // @[:@38073.4]
  assign x653_rdcol_1_io_a = RetimeWrapper_47_io_out; // @[Math.scala 151:17:@38074.4]
  assign x653_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@38075.4]
  assign x653_rdcol_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38076.4]
  assign x659_sum_1_clock = clock; // @[:@38104.4]
  assign x659_sum_1_reset = reset; // @[:@38105.4]
  assign x659_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@38106.4]
  assign x659_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@38107.4]
  assign x659_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38108.4]
  assign RetimeWrapper_52_clock = clock; // @[:@38114.4]
  assign RetimeWrapper_52_reset = reset; // @[:@38115.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38117.4]
  assign RetimeWrapper_52_io_in = ~ x655; // @[package.scala 94:16:@38116.4]
  assign RetimeWrapper_53_clock = clock; // @[:@38128.4]
  assign RetimeWrapper_53_reset = reset; // @[:@38129.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38131.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38130.4]
  assign x665_rdcol_1_clock = clock; // @[:@38151.4]
  assign x665_rdcol_1_reset = reset; // @[:@38152.4]
  assign x665_rdcol_1_io_a = RetimeWrapper_47_io_out; // @[Math.scala 151:17:@38153.4]
  assign x665_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@38154.4]
  assign x665_rdcol_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38155.4]
  assign x671_sum_1_clock = clock; // @[:@38183.4]
  assign x671_sum_1_reset = reset; // @[:@38184.4]
  assign x671_sum_1_io_a = {_T_787,_T_788}; // @[Math.scala 151:17:@38185.4]
  assign x671_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@38186.4]
  assign x671_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38187.4]
  assign RetimeWrapper_54_clock = clock; // @[:@38193.4]
  assign RetimeWrapper_54_reset = reset; // @[:@38194.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38196.4]
  assign RetimeWrapper_54_io_in = ~ x667; // @[package.scala 94:16:@38195.4]
  assign RetimeWrapper_55_clock = clock; // @[:@38207.4]
  assign RetimeWrapper_55_reset = reset; // @[:@38208.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38210.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38209.4]
  assign RetimeWrapper_56_clock = clock; // @[:@38228.4]
  assign RetimeWrapper_56_reset = reset; // @[:@38229.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38231.4]
  assign RetimeWrapper_56_io_in = __io_result; // @[package.scala 94:16:@38230.4]
  assign RetimeWrapper_57_clock = clock; // @[:@38255.4]
  assign RetimeWrapper_57_reset = reset; // @[:@38256.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38258.4]
  assign RetimeWrapper_57_io_in = $signed(_T_1103) < $signed(32'sh0); // @[package.scala 94:16:@38257.4]
  assign RetimeWrapper_58_clock = clock; // @[:@38290.4]
  assign RetimeWrapper_58_reset = reset; // @[:@38291.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38293.4]
  assign RetimeWrapper_58_io_in = {_T_1142,_T_1143}; // @[package.scala 94:16:@38292.4]
  assign x683_sum_1_clock = clock; // @[:@38299.4]
  assign x683_sum_1_reset = reset; // @[:@38300.4]
  assign x683_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@38301.4]
  assign x683_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@38302.4]
  assign x683_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38303.4]
  assign RetimeWrapper_59_clock = clock; // @[:@38309.4]
  assign RetimeWrapper_59_reset = reset; // @[:@38310.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38312.4]
  assign RetimeWrapper_59_io_in = ~ x679; // @[package.scala 94:16:@38311.4]
  assign RetimeWrapper_60_clock = clock; // @[:@38318.4]
  assign RetimeWrapper_60_reset = reset; // @[:@38319.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38321.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1133); // @[package.scala 94:16:@38320.4]
  assign RetimeWrapper_61_clock = clock; // @[:@38332.4]
  assign RetimeWrapper_61_reset = reset; // @[:@38333.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38335.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38334.4]
  assign x691_sum_1_clock = clock; // @[:@38361.4]
  assign x691_sum_1_reset = reset; // @[:@38362.4]
  assign x691_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@38363.4]
  assign x691_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@38364.4]
  assign x691_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38365.4]
  assign RetimeWrapper_62_clock = clock; // @[:@38371.4]
  assign RetimeWrapper_62_reset = reset; // @[:@38372.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38374.4]
  assign RetimeWrapper_62_io_in = ~ x689; // @[package.scala 94:16:@38373.4]
  assign RetimeWrapper_63_clock = clock; // @[:@38385.4]
  assign RetimeWrapper_63_reset = reset; // @[:@38386.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38388.4]
  assign RetimeWrapper_63_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38387.4]
  assign x698_sum_1_clock = clock; // @[:@38412.4]
  assign x698_sum_1_reset = reset; // @[:@38413.4]
  assign x698_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@38414.4]
  assign x698_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@38415.4]
  assign x698_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38416.4]
  assign RetimeWrapper_64_clock = clock; // @[:@38422.4]
  assign RetimeWrapper_64_reset = reset; // @[:@38423.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38425.4]
  assign RetimeWrapper_64_io_in = ~ x696; // @[package.scala 94:16:@38424.4]
  assign RetimeWrapper_65_clock = clock; // @[:@38436.4]
  assign RetimeWrapper_65_reset = reset; // @[:@38437.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38439.4]
  assign RetimeWrapper_65_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38438.4]
  assign RetimeWrapper_66_clock = clock; // @[:@38463.4]
  assign RetimeWrapper_66_reset = reset; // @[:@38464.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38466.4]
  assign RetimeWrapper_66_io_in = {_T_341,_T_342}; // @[package.scala 94:16:@38465.4]
  assign x705_sum_1_clock = clock; // @[:@38472.4]
  assign x705_sum_1_reset = reset; // @[:@38473.4]
  assign x705_sum_1_io_a = {_T_1142,_T_1143}; // @[Math.scala 151:17:@38474.4]
  assign x705_sum_1_io_b = RetimeWrapper_66_io_out; // @[Math.scala 152:17:@38475.4]
  assign x705_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38476.4]
  assign RetimeWrapper_67_clock = clock; // @[:@38482.4]
  assign RetimeWrapper_67_reset = reset; // @[:@38483.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38485.4]
  assign RetimeWrapper_67_io_in = ~ x703; // @[package.scala 94:16:@38484.4]
  assign RetimeWrapper_68_clock = clock; // @[:@38491.4]
  assign RetimeWrapper_68_reset = reset; // @[:@38492.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38494.4]
  assign RetimeWrapper_68_io_in = x705_sum_1_io_result; // @[package.scala 94:16:@38493.4]
  assign RetimeWrapper_69_clock = clock; // @[:@38505.4]
  assign RetimeWrapper_69_reset = reset; // @[:@38506.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38508.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38507.4]
  assign x712_sum_1_clock = clock; // @[:@38532.4]
  assign x712_sum_1_reset = reset; // @[:@38533.4]
  assign x712_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@38534.4]
  assign x712_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@38535.4]
  assign x712_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38536.4]
  assign RetimeWrapper_70_clock = clock; // @[:@38542.4]
  assign RetimeWrapper_70_reset = reset; // @[:@38543.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38545.4]
  assign RetimeWrapper_70_io_in = ~ x710; // @[package.scala 94:16:@38544.4]
  assign RetimeWrapper_71_clock = clock; // @[:@38556.4]
  assign RetimeWrapper_71_reset = reset; // @[:@38557.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38559.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38558.4]
  assign x719_sum_1_clock = clock; // @[:@38583.4]
  assign x719_sum_1_reset = reset; // @[:@38584.4]
  assign x719_sum_1_io_a = RetimeWrapper_58_io_out; // @[Math.scala 151:17:@38585.4]
  assign x719_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@38586.4]
  assign x719_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38587.4]
  assign RetimeWrapper_72_clock = clock; // @[:@38593.4]
  assign RetimeWrapper_72_reset = reset; // @[:@38594.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38596.4]
  assign RetimeWrapper_72_io_in = ~ x717; // @[package.scala 94:16:@38595.4]
  assign RetimeWrapper_73_clock = clock; // @[:@38607.4]
  assign RetimeWrapper_73_reset = reset; // @[:@38608.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38610.4]
  assign RetimeWrapper_73_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38609.4]
  assign x724_rdrow_1_clock = clock; // @[:@38630.4]
  assign x724_rdrow_1_reset = reset; // @[:@38631.4]
  assign x724_rdrow_1_io_a = RetimeWrapper_56_io_out; // @[Math.scala 151:17:@38632.4]
  assign x724_rdrow_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@38633.4]
  assign x724_rdrow_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38634.4]
  assign x731_sum_1_clock = clock; // @[:@38684.4]
  assign x731_sum_1_reset = reset; // @[:@38685.4]
  assign x731_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@38686.4]
  assign x731_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@38687.4]
  assign x731_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38688.4]
  assign RetimeWrapper_74_clock = clock; // @[:@38694.4]
  assign RetimeWrapper_74_reset = reset; // @[:@38695.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38697.4]
  assign RetimeWrapper_74_io_in = $unsigned(_T_1394); // @[package.scala 94:16:@38696.4]
  assign RetimeWrapper_75_clock = clock; // @[:@38703.4]
  assign RetimeWrapper_75_reset = reset; // @[:@38704.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38706.4]
  assign RetimeWrapper_75_io_in = ~ x727; // @[package.scala 94:16:@38705.4]
  assign RetimeWrapper_76_clock = clock; // @[:@38717.4]
  assign RetimeWrapper_76_reset = reset; // @[:@38718.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38720.4]
  assign RetimeWrapper_76_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38719.4]
  assign x739_sum_1_clock = clock; // @[:@38746.4]
  assign x739_sum_1_reset = reset; // @[:@38747.4]
  assign x739_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@38748.4]
  assign x739_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@38749.4]
  assign x739_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38750.4]
  assign RetimeWrapper_77_clock = clock; // @[:@38756.4]
  assign RetimeWrapper_77_reset = reset; // @[:@38757.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38759.4]
  assign RetimeWrapper_77_io_in = ~ x737; // @[package.scala 94:16:@38758.4]
  assign RetimeWrapper_78_clock = clock; // @[:@38770.4]
  assign RetimeWrapper_78_reset = reset; // @[:@38771.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38773.4]
  assign RetimeWrapper_78_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38772.4]
  assign x746_sum_1_clock = clock; // @[:@38797.4]
  assign x746_sum_1_reset = reset; // @[:@38798.4]
  assign x746_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@38799.4]
  assign x746_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@38800.4]
  assign x746_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38801.4]
  assign RetimeWrapper_79_clock = clock; // @[:@38807.4]
  assign RetimeWrapper_79_reset = reset; // @[:@38808.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38810.4]
  assign RetimeWrapper_79_io_in = ~ x744; // @[package.scala 94:16:@38809.4]
  assign RetimeWrapper_80_clock = clock; // @[:@38821.4]
  assign RetimeWrapper_80_reset = reset; // @[:@38822.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38824.4]
  assign RetimeWrapper_80_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38823.4]
  assign x753_sum_1_clock = clock; // @[:@38848.4]
  assign x753_sum_1_reset = reset; // @[:@38849.4]
  assign x753_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@38850.4]
  assign x753_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@38851.4]
  assign x753_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38852.4]
  assign RetimeWrapper_81_clock = clock; // @[:@38858.4]
  assign RetimeWrapper_81_reset = reset; // @[:@38859.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38861.4]
  assign RetimeWrapper_81_io_in = ~ x751; // @[package.scala 94:16:@38860.4]
  assign RetimeWrapper_82_clock = clock; // @[:@38872.4]
  assign RetimeWrapper_82_reset = reset; // @[:@38873.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38875.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38874.4]
  assign x760_sum_1_clock = clock; // @[:@38899.4]
  assign x760_sum_1_reset = reset; // @[:@38900.4]
  assign x760_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@38901.4]
  assign x760_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@38902.4]
  assign x760_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38903.4]
  assign RetimeWrapper_83_clock = clock; // @[:@38909.4]
  assign RetimeWrapper_83_reset = reset; // @[:@38910.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38912.4]
  assign RetimeWrapper_83_io_in = ~ x758; // @[package.scala 94:16:@38911.4]
  assign RetimeWrapper_84_clock = clock; // @[:@38923.4]
  assign RetimeWrapper_84_reset = reset; // @[:@38924.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38926.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38925.4]
  assign x767_sum_1_clock = clock; // @[:@38950.4]
  assign x767_sum_1_reset = reset; // @[:@38951.4]
  assign x767_sum_1_io_a = {_T_1403,_T_1404}; // @[Math.scala 151:17:@38952.4]
  assign x767_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@38953.4]
  assign x767_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@38954.4]
  assign RetimeWrapper_85_clock = clock; // @[:@38960.4]
  assign RetimeWrapper_85_reset = reset; // @[:@38961.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38963.4]
  assign RetimeWrapper_85_io_in = ~ x765; // @[package.scala 94:16:@38962.4]
  assign RetimeWrapper_86_clock = clock; // @[:@38974.4]
  assign RetimeWrapper_86_reset = reset; // @[:@38975.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38977.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38976.4]
  assign x772_rdrow_1_clock = clock; // @[:@38997.4]
  assign x772_rdrow_1_reset = reset; // @[:@38998.4]
  assign x772_rdrow_1_io_a = RetimeWrapper_56_io_out; // @[Math.scala 151:17:@38999.4]
  assign x772_rdrow_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@39000.4]
  assign x772_rdrow_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39001.4]
  assign x779_sum_1_clock = clock; // @[:@39051.4]
  assign x779_sum_1_reset = reset; // @[:@39052.4]
  assign x779_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@39053.4]
  assign x779_sum_1_io_b = RetimeWrapper_33_io_out; // @[Math.scala 152:17:@39054.4]
  assign x779_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39055.4]
  assign RetimeWrapper_87_clock = clock; // @[:@39061.4]
  assign RetimeWrapper_87_reset = reset; // @[:@39062.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39064.4]
  assign RetimeWrapper_87_io_in = $unsigned(_T_1646); // @[package.scala 94:16:@39063.4]
  assign RetimeWrapper_88_clock = clock; // @[:@39070.4]
  assign RetimeWrapper_88_reset = reset; // @[:@39071.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39073.4]
  assign RetimeWrapper_88_io_in = ~ x775; // @[package.scala 94:16:@39072.4]
  assign RetimeWrapper_89_clock = clock; // @[:@39084.4]
  assign RetimeWrapper_89_reset = reset; // @[:@39085.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39087.4]
  assign RetimeWrapper_89_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39086.4]
  assign x787_sum_1_clock = clock; // @[:@39111.4]
  assign x787_sum_1_reset = reset; // @[:@39112.4]
  assign x787_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@39113.4]
  assign x787_sum_1_io_b = RetimeWrapper_40_io_out; // @[Math.scala 152:17:@39114.4]
  assign x787_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39115.4]
  assign RetimeWrapper_90_clock = clock; // @[:@39121.4]
  assign RetimeWrapper_90_reset = reset; // @[:@39122.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39124.4]
  assign RetimeWrapper_90_io_in = ~ x785; // @[package.scala 94:16:@39123.4]
  assign RetimeWrapper_91_clock = clock; // @[:@39135.4]
  assign RetimeWrapper_91_reset = reset; // @[:@39136.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39138.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39137.4]
  assign x794_sum_1_clock = clock; // @[:@39164.4]
  assign x794_sum_1_reset = reset; // @[:@39165.4]
  assign x794_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@39166.4]
  assign x794_sum_1_io_b = RetimeWrapper_44_io_out; // @[Math.scala 152:17:@39167.4]
  assign x794_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39168.4]
  assign RetimeWrapper_92_clock = clock; // @[:@39174.4]
  assign RetimeWrapper_92_reset = reset; // @[:@39175.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39177.4]
  assign RetimeWrapper_92_io_in = ~ x792; // @[package.scala 94:16:@39176.4]
  assign RetimeWrapper_93_clock = clock; // @[:@39188.4]
  assign RetimeWrapper_93_reset = reset; // @[:@39189.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39191.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39190.4]
  assign x801_sum_1_clock = clock; // @[:@39215.4]
  assign x801_sum_1_reset = reset; // @[:@39216.4]
  assign x801_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@39217.4]
  assign x801_sum_1_io_b = RetimeWrapper_49_io_out; // @[Math.scala 152:17:@39218.4]
  assign x801_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39219.4]
  assign RetimeWrapper_94_clock = clock; // @[:@39225.4]
  assign RetimeWrapper_94_reset = reset; // @[:@39226.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39228.4]
  assign RetimeWrapper_94_io_in = ~ x799; // @[package.scala 94:16:@39227.4]
  assign RetimeWrapper_95_clock = clock; // @[:@39239.4]
  assign RetimeWrapper_95_reset = reset; // @[:@39240.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39242.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39241.4]
  assign x808_sum_1_clock = clock; // @[:@39266.4]
  assign x808_sum_1_reset = reset; // @[:@39267.4]
  assign x808_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@39268.4]
  assign x808_sum_1_io_b = {_T_1003,_T_1004}; // @[Math.scala 152:17:@39269.4]
  assign x808_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39270.4]
  assign RetimeWrapper_96_clock = clock; // @[:@39276.4]
  assign RetimeWrapper_96_reset = reset; // @[:@39277.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39279.4]
  assign RetimeWrapper_96_io_in = ~ x806; // @[package.scala 94:16:@39278.4]
  assign RetimeWrapper_97_clock = clock; // @[:@39290.4]
  assign RetimeWrapper_97_reset = reset; // @[:@39291.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39293.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39292.4]
  assign x815_sum_1_clock = clock; // @[:@39317.4]
  assign x815_sum_1_reset = reset; // @[:@39318.4]
  assign x815_sum_1_io_a = {_T_1655,_T_1656}; // @[Math.scala 151:17:@39319.4]
  assign x815_sum_1_io_b = {_T_1061,_T_1062}; // @[Math.scala 152:17:@39320.4]
  assign x815_sum_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39321.4]
  assign RetimeWrapper_98_clock = clock; // @[:@39327.4]
  assign RetimeWrapper_98_reset = reset; // @[:@39328.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39330.4]
  assign RetimeWrapper_98_io_in = ~ x813; // @[package.scala 94:16:@39329.4]
  assign RetimeWrapper_99_clock = clock; // @[:@39341.4]
  assign RetimeWrapper_99_reset = reset; // @[:@39342.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39344.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@39343.4]
  assign x825_x17_1_clock = clock; // @[:@39387.4]
  assign x825_x17_1_reset = reset; // @[:@39388.4]
  assign x825_x17_1_io_a = x539_lb_0_io_rPort_17_output_0; // @[Math.scala 151:17:@39389.4]
  assign x825_x17_1_io_b = _T_1860[7:0]; // @[Math.scala 152:17:@39390.4]
  assign x825_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39391.4]
  assign x826_x18_1_clock = clock; // @[:@39397.4]
  assign x826_x18_1_reset = reset; // @[:@39398.4]
  assign x826_x18_1_io_a = x539_lb_0_io_rPort_16_output_0; // @[Math.scala 151:17:@39399.4]
  assign x826_x18_1_io_b = _T_1864[7:0]; // @[Math.scala 152:17:@39400.4]
  assign x826_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39401.4]
  assign x827_x17_1_clock = clock; // @[:@39407.4]
  assign x827_x17_1_reset = reset; // @[:@39408.4]
  assign x827_x17_1_io_a = _T_1868[7:0]; // @[Math.scala 151:17:@39409.4]
  assign x827_x17_1_io_b = _T_1872[7:0]; // @[Math.scala 152:17:@39410.4]
  assign x827_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39411.4]
  assign x828_x18_1_clock = clock; // @[:@39417.4]
  assign x828_x18_1_reset = reset; // @[:@39418.4]
  assign x828_x18_1_io_a = x539_lb_0_io_rPort_21_output_0; // @[Math.scala 151:17:@39419.4]
  assign x828_x18_1_io_b = _T_1876[7:0]; // @[Math.scala 152:17:@39420.4]
  assign x828_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39421.4]
  assign x829_x17_1_io_a = x825_x17_1_io_result; // @[Math.scala 151:17:@39429.4]
  assign x829_x17_1_io_b = x826_x18_1_io_result; // @[Math.scala 152:17:@39430.4]
  assign x830_x18_1_io_a = x827_x17_1_io_result; // @[Math.scala 151:17:@39439.4]
  assign x830_x18_1_io_b = x828_x18_1_io_result; // @[Math.scala 152:17:@39440.4]
  assign x831_x17_1_io_a = x829_x17_1_io_result; // @[Math.scala 151:17:@39449.4]
  assign x831_x17_1_io_b = x830_x18_1_io_result; // @[Math.scala 152:17:@39450.4]
  assign RetimeWrapper_100_clock = clock; // @[:@39457.4]
  assign RetimeWrapper_100_reset = reset; // @[:@39458.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39460.4]
  assign RetimeWrapper_100_io_in = x539_lb_0_io_rPort_15_output_0; // @[package.scala 94:16:@39459.4]
  assign x832_sum_1_io_a = x831_x17_1_io_result; // @[Math.scala 151:17:@39468.4]
  assign x832_sum_1_io_b = RetimeWrapper_100_io_out; // @[Math.scala 152:17:@39469.4]
  assign RetimeWrapper_101_clock = clock; // @[:@39480.4]
  assign RetimeWrapper_101_reset = reset; // @[:@39481.4]
  assign RetimeWrapper_101_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@39483.4]
  assign RetimeWrapper_101_io_in = {4'h0,_T_1912}; // @[package.scala 94:16:@39482.4]
  assign RetimeWrapper_102_clock = clock; // @[:@39490.4]
  assign RetimeWrapper_102_reset = reset; // @[:@39491.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39493.4]
  assign RetimeWrapper_102_io_in = x539_lb_0_io_rPort_17_output_0; // @[package.scala 94:16:@39492.4]
  assign x834_sub_1_io_a = RetimeWrapper_102_io_out; // @[Math.scala 192:17:@39501.4]
  assign x834_sub_1_io_b = RetimeWrapper_101_io_out; // @[Math.scala 193:17:@39502.4]
  assign RetimeWrapper_103_clock = clock; // @[:@39524.4]
  assign RetimeWrapper_103_reset = reset; // @[:@39525.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39527.4]
  assign RetimeWrapper_103_io_in = x835 ? x834_sub_number : 8'h0; // @[package.scala 94:16:@39526.4]
  assign x838_div_1_clock = clock; // @[:@39535.4]
  assign x838_div_1_reset = reset; // @[:@39536.4]
  assign x838_div_1_io_a = RetimeWrapper_103_io_out; // @[Math.scala 328:17:@39537.4]
  assign x838_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@39539.4]
  assign RetimeWrapper_104_clock = clock; // @[:@39545.4]
  assign RetimeWrapper_104_reset = reset; // @[:@39546.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39548.4]
  assign RetimeWrapper_104_io_in = x539_lb_0_io_rPort_17_output_0; // @[package.scala 94:16:@39547.4]
  assign x839_sum_1_io_a = RetimeWrapper_104_io_out; // @[Math.scala 151:17:@39556.4]
  assign x839_sum_1_io_b = x838_div_1_io_result; // @[Math.scala 152:17:@39557.4]
  assign RetimeWrapper_105_clock = clock; // @[:@39564.4]
  assign RetimeWrapper_105_reset = reset; // @[:@39565.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39567.4]
  assign RetimeWrapper_105_io_in = RetimeWrapper_101_io_out; // @[package.scala 94:16:@39566.4]
  assign RetimeWrapper_106_clock = clock; // @[:@39573.4]
  assign RetimeWrapper_106_reset = reset; // @[:@39574.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39576.4]
  assign RetimeWrapper_106_io_in = x833_number == 8'h0; // @[package.scala 94:16:@39575.4]
  assign x846_x17_1_clock = clock; // @[:@39612.4]
  assign x846_x17_1_reset = reset; // @[:@39613.4]
  assign x846_x17_1_io_a = x539_lb_0_io_rPort_22_output_0; // @[Math.scala 151:17:@39614.4]
  assign x846_x17_1_io_b = _T_1969[7:0]; // @[Math.scala 152:17:@39615.4]
  assign x846_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39616.4]
  assign x847_x18_1_clock = clock; // @[:@39622.4]
  assign x847_x18_1_reset = reset; // @[:@39623.4]
  assign x847_x18_1_io_a = x539_lb_0_io_rPort_2_output_0; // @[Math.scala 151:17:@39624.4]
  assign x847_x18_1_io_b = _T_1973[7:0]; // @[Math.scala 152:17:@39625.4]
  assign x847_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39626.4]
  assign x848_x17_1_clock = clock; // @[:@39632.4]
  assign x848_x17_1_reset = reset; // @[:@39633.4]
  assign x848_x17_1_io_a = _T_1977[7:0]; // @[Math.scala 151:17:@39634.4]
  assign x848_x17_1_io_b = _T_1981[7:0]; // @[Math.scala 152:17:@39635.4]
  assign x848_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39636.4]
  assign x849_x18_1_clock = clock; // @[:@39642.4]
  assign x849_x18_1_reset = reset; // @[:@39643.4]
  assign x849_x18_1_io_a = x539_lb_0_io_rPort_6_output_0; // @[Math.scala 151:17:@39644.4]
  assign x849_x18_1_io_b = _T_1985[7:0]; // @[Math.scala 152:17:@39645.4]
  assign x849_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39646.4]
  assign x850_x17_1_io_a = x846_x17_1_io_result; // @[Math.scala 151:17:@39654.4]
  assign x850_x17_1_io_b = x847_x18_1_io_result; // @[Math.scala 152:17:@39655.4]
  assign x851_x18_1_io_a = x848_x17_1_io_result; // @[Math.scala 151:17:@39664.4]
  assign x851_x18_1_io_b = x849_x18_1_io_result; // @[Math.scala 152:17:@39665.4]
  assign x852_x17_1_io_a = x850_x17_1_io_result; // @[Math.scala 151:17:@39674.4]
  assign x852_x17_1_io_b = x851_x18_1_io_result; // @[Math.scala 152:17:@39675.4]
  assign RetimeWrapper_107_clock = clock; // @[:@39682.4]
  assign RetimeWrapper_107_reset = reset; // @[:@39683.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39685.4]
  assign RetimeWrapper_107_io_in = x539_lb_0_io_rPort_4_output_0; // @[package.scala 94:16:@39684.4]
  assign x853_sum_1_io_a = x852_x17_1_io_result; // @[Math.scala 151:17:@39693.4]
  assign x853_sum_1_io_b = RetimeWrapper_107_io_out; // @[Math.scala 152:17:@39694.4]
  assign RetimeWrapper_108_clock = clock; // @[:@39705.4]
  assign RetimeWrapper_108_reset = reset; // @[:@39706.4]
  assign RetimeWrapper_108_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@39708.4]
  assign RetimeWrapper_108_io_in = {4'h0,_T_2021}; // @[package.scala 94:16:@39707.4]
  assign RetimeWrapper_109_clock = clock; // @[:@39715.4]
  assign RetimeWrapper_109_reset = reset; // @[:@39716.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39718.4]
  assign RetimeWrapper_109_io_in = x539_lb_0_io_rPort_22_output_0; // @[package.scala 94:16:@39717.4]
  assign x855_sub_1_io_a = RetimeWrapper_109_io_out; // @[Math.scala 192:17:@39726.4]
  assign x855_sub_1_io_b = RetimeWrapper_108_io_out; // @[Math.scala 193:17:@39727.4]
  assign RetimeWrapper_110_clock = clock; // @[:@39749.4]
  assign RetimeWrapper_110_reset = reset; // @[:@39750.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39752.4]
  assign RetimeWrapper_110_io_in = x856 ? x855_sub_number : 8'h0; // @[package.scala 94:16:@39751.4]
  assign x859_div_1_clock = clock; // @[:@39760.4]
  assign x859_div_1_reset = reset; // @[:@39761.4]
  assign x859_div_1_io_a = RetimeWrapper_110_io_out; // @[Math.scala 328:17:@39762.4]
  assign x859_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@39764.4]
  assign RetimeWrapper_111_clock = clock; // @[:@39770.4]
  assign RetimeWrapper_111_reset = reset; // @[:@39771.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39773.4]
  assign RetimeWrapper_111_io_in = x539_lb_0_io_rPort_22_output_0; // @[package.scala 94:16:@39772.4]
  assign x860_sum_1_io_a = RetimeWrapper_111_io_out; // @[Math.scala 151:17:@39781.4]
  assign x860_sum_1_io_b = x859_div_1_io_result; // @[Math.scala 152:17:@39782.4]
  assign RetimeWrapper_112_clock = clock; // @[:@39789.4]
  assign RetimeWrapper_112_reset = reset; // @[:@39790.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39792.4]
  assign RetimeWrapper_112_io_in = RetimeWrapper_108_io_out; // @[package.scala 94:16:@39791.4]
  assign RetimeWrapper_113_clock = clock; // @[:@39798.4]
  assign RetimeWrapper_113_reset = reset; // @[:@39799.4]
  assign RetimeWrapper_113_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39801.4]
  assign RetimeWrapper_113_io_in = x854_number == 8'h0; // @[package.scala 94:16:@39800.4]
  assign x866_x17_1_clock = clock; // @[:@39830.4]
  assign x866_x17_1_reset = reset; // @[:@39831.4]
  assign x866_x17_1_io_a = x539_lb_0_io_rPort_16_output_0; // @[Math.scala 151:17:@39832.4]
  assign x866_x17_1_io_b = _T_2076[7:0]; // @[Math.scala 152:17:@39833.4]
  assign x866_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39834.4]
  assign x867_x18_1_clock = clock; // @[:@39840.4]
  assign x867_x18_1_reset = reset; // @[:@39841.4]
  assign x867_x18_1_io_a = x539_lb_0_io_rPort_14_output_0; // @[Math.scala 151:17:@39842.4]
  assign x867_x18_1_io_b = _T_1872[7:0]; // @[Math.scala 152:17:@39843.4]
  assign x867_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39844.4]
  assign x868_x17_1_clock = clock; // @[:@39850.4]
  assign x868_x17_1_reset = reset; // @[:@39851.4]
  assign x868_x17_1_io_a = _T_2080[7:0]; // @[Math.scala 151:17:@39852.4]
  assign x868_x17_1_io_b = _T_2084[7:0]; // @[Math.scala 152:17:@39853.4]
  assign x868_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39854.4]
  assign x869_x18_1_clock = clock; // @[:@39860.4]
  assign x869_x18_1_reset = reset; // @[:@39861.4]
  assign x869_x18_1_io_a = x539_lb_0_io_rPort_15_output_0; // @[Math.scala 151:17:@39862.4]
  assign x869_x18_1_io_b = _T_2088[7:0]; // @[Math.scala 152:17:@39863.4]
  assign x869_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@39864.4]
  assign x870_x17_1_io_a = x866_x17_1_io_result; // @[Math.scala 151:17:@39872.4]
  assign x870_x17_1_io_b = x867_x18_1_io_result; // @[Math.scala 152:17:@39873.4]
  assign x871_x18_1_io_a = x868_x17_1_io_result; // @[Math.scala 151:17:@39882.4]
  assign x871_x18_1_io_b = x869_x18_1_io_result; // @[Math.scala 152:17:@39883.4]
  assign x872_x17_1_io_a = x870_x17_1_io_result; // @[Math.scala 151:17:@39892.4]
  assign x872_x17_1_io_b = x871_x18_1_io_result; // @[Math.scala 152:17:@39893.4]
  assign RetimeWrapper_114_clock = clock; // @[:@39900.4]
  assign RetimeWrapper_114_reset = reset; // @[:@39901.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39903.4]
  assign RetimeWrapper_114_io_in = x539_lb_0_io_rPort_18_output_0; // @[package.scala 94:16:@39902.4]
  assign x873_sum_1_io_a = x872_x17_1_io_result; // @[Math.scala 151:17:@39911.4]
  assign x873_sum_1_io_b = RetimeWrapper_114_io_out; // @[Math.scala 152:17:@39912.4]
  assign RetimeWrapper_115_clock = clock; // @[:@39923.4]
  assign RetimeWrapper_115_reset = reset; // @[:@39924.4]
  assign RetimeWrapper_115_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@39926.4]
  assign RetimeWrapper_115_io_in = {4'h0,_T_2124}; // @[package.scala 94:16:@39925.4]
  assign RetimeWrapper_116_clock = clock; // @[:@39933.4]
  assign RetimeWrapper_116_reset = reset; // @[:@39934.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39936.4]
  assign RetimeWrapper_116_io_in = x539_lb_0_io_rPort_16_output_0; // @[package.scala 94:16:@39935.4]
  assign x875_sub_1_io_a = RetimeWrapper_116_io_out; // @[Math.scala 192:17:@39944.4]
  assign x875_sub_1_io_b = RetimeWrapper_115_io_out; // @[Math.scala 193:17:@39945.4]
  assign RetimeWrapper_117_clock = clock; // @[:@39967.4]
  assign RetimeWrapper_117_reset = reset; // @[:@39968.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39970.4]
  assign RetimeWrapper_117_io_in = x876 ? x875_sub_number : 8'h0; // @[package.scala 94:16:@39969.4]
  assign x879_div_1_clock = clock; // @[:@39978.4]
  assign x879_div_1_reset = reset; // @[:@39979.4]
  assign x879_div_1_io_a = RetimeWrapper_117_io_out; // @[Math.scala 328:17:@39980.4]
  assign x879_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@39982.4]
  assign RetimeWrapper_118_clock = clock; // @[:@39988.4]
  assign RetimeWrapper_118_reset = reset; // @[:@39989.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@39991.4]
  assign RetimeWrapper_118_io_in = x539_lb_0_io_rPort_16_output_0; // @[package.scala 94:16:@39990.4]
  assign x880_sum_1_io_a = RetimeWrapper_118_io_out; // @[Math.scala 151:17:@40001.4]
  assign x880_sum_1_io_b = x879_div_1_io_result; // @[Math.scala 152:17:@40002.4]
  assign RetimeWrapper_119_clock = clock; // @[:@40009.4]
  assign RetimeWrapper_119_reset = reset; // @[:@40010.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40012.4]
  assign RetimeWrapper_119_io_in = RetimeWrapper_115_io_out; // @[package.scala 94:16:@40011.4]
  assign RetimeWrapper_120_clock = clock; // @[:@40018.4]
  assign RetimeWrapper_120_reset = reset; // @[:@40019.4]
  assign RetimeWrapper_120_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40021.4]
  assign RetimeWrapper_120_io_in = x874_number == 8'h0; // @[package.scala 94:16:@40020.4]
  assign x886_x17_1_clock = clock; // @[:@40050.4]
  assign x886_x17_1_reset = reset; // @[:@40051.4]
  assign x886_x17_1_io_a = x539_lb_0_io_rPort_2_output_0; // @[Math.scala 151:17:@40052.4]
  assign x886_x17_1_io_b = _T_2181[7:0]; // @[Math.scala 152:17:@40053.4]
  assign x886_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40054.4]
  assign x887_x18_1_clock = clock; // @[:@40060.4]
  assign x887_x18_1_reset = reset; // @[:@40061.4]
  assign x887_x18_1_io_a = x539_lb_0_io_rPort_13_output_0; // @[Math.scala 151:17:@40062.4]
  assign x887_x18_1_io_b = _T_1981[7:0]; // @[Math.scala 152:17:@40063.4]
  assign x887_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40064.4]
  assign x888_x17_1_clock = clock; // @[:@40070.4]
  assign x888_x17_1_reset = reset; // @[:@40071.4]
  assign x888_x17_1_io_a = _T_2185[7:0]; // @[Math.scala 151:17:@40072.4]
  assign x888_x17_1_io_b = _T_2189[7:0]; // @[Math.scala 152:17:@40073.4]
  assign x888_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40074.4]
  assign x889_x18_1_clock = clock; // @[:@40080.4]
  assign x889_x18_1_reset = reset; // @[:@40081.4]
  assign x889_x18_1_io_a = x539_lb_0_io_rPort_4_output_0; // @[Math.scala 151:17:@40082.4]
  assign x889_x18_1_io_b = _T_2193[7:0]; // @[Math.scala 152:17:@40083.4]
  assign x889_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40084.4]
  assign x890_x17_1_io_a = x886_x17_1_io_result; // @[Math.scala 151:17:@40092.4]
  assign x890_x17_1_io_b = x887_x18_1_io_result; // @[Math.scala 152:17:@40093.4]
  assign x891_x18_1_io_a = x888_x17_1_io_result; // @[Math.scala 151:17:@40102.4]
  assign x891_x18_1_io_b = x889_x18_1_io_result; // @[Math.scala 152:17:@40103.4]
  assign x892_x17_1_io_a = x890_x17_1_io_result; // @[Math.scala 151:17:@40112.4]
  assign x892_x17_1_io_b = x891_x18_1_io_result; // @[Math.scala 152:17:@40113.4]
  assign RetimeWrapper_121_clock = clock; // @[:@40120.4]
  assign RetimeWrapper_121_reset = reset; // @[:@40121.4]
  assign RetimeWrapper_121_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40123.4]
  assign RetimeWrapper_121_io_in = x539_lb_0_io_rPort_3_output_0; // @[package.scala 94:16:@40122.4]
  assign x893_sum_1_io_a = x892_x17_1_io_result; // @[Math.scala 151:17:@40131.4]
  assign x893_sum_1_io_b = RetimeWrapper_121_io_out; // @[Math.scala 152:17:@40132.4]
  assign RetimeWrapper_122_clock = clock; // @[:@40143.4]
  assign RetimeWrapper_122_reset = reset; // @[:@40144.4]
  assign RetimeWrapper_122_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@40146.4]
  assign RetimeWrapper_122_io_in = {4'h0,_T_2229}; // @[package.scala 94:16:@40145.4]
  assign RetimeWrapper_123_clock = clock; // @[:@40153.4]
  assign RetimeWrapper_123_reset = reset; // @[:@40154.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40156.4]
  assign RetimeWrapper_123_io_in = x539_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@40155.4]
  assign x895_sub_1_io_a = RetimeWrapper_123_io_out; // @[Math.scala 192:17:@40164.4]
  assign x895_sub_1_io_b = RetimeWrapper_122_io_out; // @[Math.scala 193:17:@40165.4]
  assign RetimeWrapper_124_clock = clock; // @[:@40187.4]
  assign RetimeWrapper_124_reset = reset; // @[:@40188.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40190.4]
  assign RetimeWrapper_124_io_in = x896 ? x895_sub_number : 8'h0; // @[package.scala 94:16:@40189.4]
  assign x899_div_1_clock = clock; // @[:@40198.4]
  assign x899_div_1_reset = reset; // @[:@40199.4]
  assign x899_div_1_io_a = RetimeWrapper_124_io_out; // @[Math.scala 328:17:@40200.4]
  assign x899_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@40202.4]
  assign RetimeWrapper_125_clock = clock; // @[:@40208.4]
  assign RetimeWrapper_125_reset = reset; // @[:@40209.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40211.4]
  assign RetimeWrapper_125_io_in = x539_lb_0_io_rPort_2_output_0; // @[package.scala 94:16:@40210.4]
  assign x900_sum_1_io_a = RetimeWrapper_125_io_out; // @[Math.scala 151:17:@40219.4]
  assign x900_sum_1_io_b = x899_div_1_io_result; // @[Math.scala 152:17:@40220.4]
  assign RetimeWrapper_126_clock = clock; // @[:@40227.4]
  assign RetimeWrapper_126_reset = reset; // @[:@40228.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40230.4]
  assign RetimeWrapper_126_io_in = RetimeWrapper_122_io_out; // @[package.scala 94:16:@40229.4]
  assign RetimeWrapper_127_clock = clock; // @[:@40236.4]
  assign RetimeWrapper_127_reset = reset; // @[:@40237.4]
  assign RetimeWrapper_127_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40239.4]
  assign RetimeWrapper_127_io_in = x894_number == 8'h0; // @[package.scala 94:16:@40238.4]
  assign x905_x17_1_clock = clock; // @[:@40263.4]
  assign x905_x17_1_reset = reset; // @[:@40264.4]
  assign x905_x17_1_io_a = x539_lb_0_io_rPort_5_output_0; // @[Math.scala 151:17:@40265.4]
  assign x905_x17_1_io_b = _T_1973[7:0]; // @[Math.scala 152:17:@40266.4]
  assign x905_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40267.4]
  assign x906_x18_1_clock = clock; // @[:@40273.4]
  assign x906_x18_1_reset = reset; // @[:@40274.4]
  assign x906_x18_1_io_a = x539_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@40275.4]
  assign x906_x18_1_io_b = _T_2284[7:0]; // @[Math.scala 152:17:@40276.4]
  assign x906_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40277.4]
  assign x907_x17_1_clock = clock; // @[:@40283.4]
  assign x907_x17_1_reset = reset; // @[:@40284.4]
  assign x907_x17_1_io_a = _T_2288[7:0]; // @[Math.scala 151:17:@40285.4]
  assign x907_x17_1_io_b = _T_1985[7:0]; // @[Math.scala 152:17:@40286.4]
  assign x907_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40287.4]
  assign x908_x18_1_clock = clock; // @[:@40293.4]
  assign x908_x18_1_reset = reset; // @[:@40294.4]
  assign x908_x18_1_io_a = x539_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@40295.4]
  assign x908_x18_1_io_b = _T_2292[7:0]; // @[Math.scala 152:17:@40296.4]
  assign x908_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40297.4]
  assign x909_x17_1_io_a = x905_x17_1_io_result; // @[Math.scala 151:17:@40305.4]
  assign x909_x17_1_io_b = x906_x18_1_io_result; // @[Math.scala 152:17:@40306.4]
  assign x910_x18_1_io_a = x907_x17_1_io_result; // @[Math.scala 151:17:@40315.4]
  assign x910_x18_1_io_b = x908_x18_1_io_result; // @[Math.scala 152:17:@40316.4]
  assign x911_x17_1_io_a = x909_x17_1_io_result; // @[Math.scala 151:17:@40325.4]
  assign x911_x17_1_io_b = x910_x18_1_io_result; // @[Math.scala 152:17:@40326.4]
  assign RetimeWrapper_128_clock = clock; // @[:@40333.4]
  assign RetimeWrapper_128_reset = reset; // @[:@40334.4]
  assign RetimeWrapper_128_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40336.4]
  assign RetimeWrapper_128_io_in = x539_lb_0_io_rPort_0_output_0; // @[package.scala 94:16:@40335.4]
  assign x912_sum_1_io_a = x911_x17_1_io_result; // @[Math.scala 151:17:@40344.4]
  assign x912_sum_1_io_b = RetimeWrapper_128_io_out; // @[Math.scala 152:17:@40345.4]
  assign RetimeWrapper_129_clock = clock; // @[:@40356.4]
  assign RetimeWrapper_129_reset = reset; // @[:@40357.4]
  assign RetimeWrapper_129_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@40359.4]
  assign RetimeWrapper_129_io_in = {4'h0,_T_2328}; // @[package.scala 94:16:@40358.4]
  assign RetimeWrapper_130_clock = clock; // @[:@40366.4]
  assign RetimeWrapper_130_reset = reset; // @[:@40367.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40369.4]
  assign RetimeWrapper_130_io_in = x539_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@40368.4]
  assign x914_sub_1_io_a = RetimeWrapper_130_io_out; // @[Math.scala 192:17:@40377.4]
  assign x914_sub_1_io_b = RetimeWrapper_129_io_out; // @[Math.scala 193:17:@40378.4]
  assign RetimeWrapper_131_clock = clock; // @[:@40400.4]
  assign RetimeWrapper_131_reset = reset; // @[:@40401.4]
  assign RetimeWrapper_131_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40403.4]
  assign RetimeWrapper_131_io_in = x915 ? x914_sub_number : 8'h0; // @[package.scala 94:16:@40402.4]
  assign x918_div_1_clock = clock; // @[:@40413.4]
  assign x918_div_1_reset = reset; // @[:@40414.4]
  assign x918_div_1_io_a = RetimeWrapper_131_io_out; // @[Math.scala 328:17:@40415.4]
  assign x918_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@40417.4]
  assign RetimeWrapper_132_clock = clock; // @[:@40423.4]
  assign RetimeWrapper_132_reset = reset; // @[:@40424.4]
  assign RetimeWrapper_132_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40426.4]
  assign RetimeWrapper_132_io_in = x539_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@40425.4]
  assign x919_sum_1_io_a = RetimeWrapper_132_io_out; // @[Math.scala 151:17:@40434.4]
  assign x919_sum_1_io_b = x918_div_1_io_result; // @[Math.scala 152:17:@40435.4]
  assign RetimeWrapper_133_clock = clock; // @[:@40442.4]
  assign RetimeWrapper_133_reset = reset; // @[:@40443.4]
  assign RetimeWrapper_133_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40445.4]
  assign RetimeWrapper_133_io_in = x913_number == 8'h0; // @[package.scala 94:16:@40444.4]
  assign RetimeWrapper_134_clock = clock; // @[:@40451.4]
  assign RetimeWrapper_134_reset = reset; // @[:@40452.4]
  assign RetimeWrapper_134_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40454.4]
  assign RetimeWrapper_134_io_in = RetimeWrapper_129_io_out; // @[package.scala 94:16:@40453.4]
  assign x923_x17_1_clock = clock; // @[:@40473.4]
  assign x923_x17_1_reset = reset; // @[:@40474.4]
  assign x923_x17_1_io_a = x539_lb_0_io_rPort_9_output_0; // @[Math.scala 151:17:@40475.4]
  assign x923_x17_1_io_b = _T_1872[7:0]; // @[Math.scala 152:17:@40476.4]
  assign x923_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40477.4]
  assign x924_x18_1_clock = clock; // @[:@40483.4]
  assign x924_x18_1_reset = reset; // @[:@40484.4]
  assign x924_x18_1_io_a = x539_lb_0_io_rPort_23_output_0; // @[Math.scala 151:17:@40485.4]
  assign x924_x18_1_io_b = _T_1876[7:0]; // @[Math.scala 152:17:@40486.4]
  assign x924_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40487.4]
  assign x925_x17_1_clock = clock; // @[:@40493.4]
  assign x925_x17_1_reset = reset; // @[:@40494.4]
  assign x925_x17_1_io_a = _T_2385[7:0]; // @[Math.scala 151:17:@40495.4]
  assign x925_x17_1_io_b = _T_2088[7:0]; // @[Math.scala 152:17:@40496.4]
  assign x925_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40497.4]
  assign x926_x18_1_clock = clock; // @[:@40503.4]
  assign x926_x18_1_reset = reset; // @[:@40504.4]
  assign x926_x18_1_io_a = x539_lb_0_io_rPort_20_output_0; // @[Math.scala 151:17:@40505.4]
  assign x926_x18_1_io_b = _T_2389[7:0]; // @[Math.scala 152:17:@40506.4]
  assign x926_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40507.4]
  assign x927_x17_1_io_a = x923_x17_1_io_result; // @[Math.scala 151:17:@40515.4]
  assign x927_x17_1_io_b = x924_x18_1_io_result; // @[Math.scala 152:17:@40516.4]
  assign x928_x18_1_io_a = x925_x17_1_io_result; // @[Math.scala 151:17:@40525.4]
  assign x928_x18_1_io_b = x926_x18_1_io_result; // @[Math.scala 152:17:@40526.4]
  assign x929_x17_1_io_a = x927_x17_1_io_result; // @[Math.scala 151:17:@40535.4]
  assign x929_x17_1_io_b = x928_x18_1_io_result; // @[Math.scala 152:17:@40536.4]
  assign RetimeWrapper_135_clock = clock; // @[:@40543.4]
  assign RetimeWrapper_135_reset = reset; // @[:@40544.4]
  assign RetimeWrapper_135_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40546.4]
  assign RetimeWrapper_135_io_in = x539_lb_0_io_rPort_10_output_0; // @[package.scala 94:16:@40545.4]
  assign x930_sum_1_io_a = x929_x17_1_io_result; // @[Math.scala 151:17:@40554.4]
  assign x930_sum_1_io_b = RetimeWrapper_135_io_out; // @[Math.scala 152:17:@40555.4]
  assign RetimeWrapper_136_clock = clock; // @[:@40566.4]
  assign RetimeWrapper_136_reset = reset; // @[:@40567.4]
  assign RetimeWrapper_136_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@40569.4]
  assign RetimeWrapper_136_io_in = {4'h0,_T_2425}; // @[package.scala 94:16:@40568.4]
  assign RetimeWrapper_137_clock = clock; // @[:@40576.4]
  assign RetimeWrapper_137_reset = reset; // @[:@40577.4]
  assign RetimeWrapper_137_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40579.4]
  assign RetimeWrapper_137_io_in = x539_lb_0_io_rPort_9_output_0; // @[package.scala 94:16:@40578.4]
  assign x932_sub_1_io_a = RetimeWrapper_137_io_out; // @[Math.scala 192:17:@40587.4]
  assign x932_sub_1_io_b = RetimeWrapper_136_io_out; // @[Math.scala 193:17:@40588.4]
  assign RetimeWrapper_138_clock = clock; // @[:@40610.4]
  assign RetimeWrapper_138_reset = reset; // @[:@40611.4]
  assign RetimeWrapper_138_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40613.4]
  assign RetimeWrapper_138_io_in = x933 ? x932_sub_number : 8'h0; // @[package.scala 94:16:@40612.4]
  assign x936_div_1_clock = clock; // @[:@40621.4]
  assign x936_div_1_reset = reset; // @[:@40622.4]
  assign x936_div_1_io_a = RetimeWrapper_138_io_out; // @[Math.scala 328:17:@40623.4]
  assign x936_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@40625.4]
  assign RetimeWrapper_139_clock = clock; // @[:@40631.4]
  assign RetimeWrapper_139_reset = reset; // @[:@40632.4]
  assign RetimeWrapper_139_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40634.4]
  assign RetimeWrapper_139_io_in = x539_lb_0_io_rPort_9_output_0; // @[package.scala 94:16:@40633.4]
  assign x937_sum_1_io_a = RetimeWrapper_139_io_out; // @[Math.scala 151:17:@40642.4]
  assign x937_sum_1_io_b = x936_div_1_io_result; // @[Math.scala 152:17:@40643.4]
  assign RetimeWrapper_140_clock = clock; // @[:@40650.4]
  assign RetimeWrapper_140_reset = reset; // @[:@40651.4]
  assign RetimeWrapper_140_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40653.4]
  assign RetimeWrapper_140_io_in = x931_number == 8'h0; // @[package.scala 94:16:@40652.4]
  assign RetimeWrapper_141_clock = clock; // @[:@40659.4]
  assign RetimeWrapper_141_reset = reset; // @[:@40660.4]
  assign RetimeWrapper_141_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40662.4]
  assign RetimeWrapper_141_io_in = RetimeWrapper_136_io_out; // @[package.scala 94:16:@40661.4]
  assign x941_x17_1_clock = clock; // @[:@40681.4]
  assign x941_x17_1_reset = reset; // @[:@40682.4]
  assign x941_x17_1_io_a = x539_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@40683.4]
  assign x941_x17_1_io_b = _T_1981[7:0]; // @[Math.scala 152:17:@40684.4]
  assign x941_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40685.4]
  assign x942_x18_1_clock = clock; // @[:@40691.4]
  assign x942_x18_1_reset = reset; // @[:@40692.4]
  assign x942_x18_1_io_a = x539_lb_0_io_rPort_1_output_0; // @[Math.scala 151:17:@40693.4]
  assign x942_x18_1_io_b = _T_1985[7:0]; // @[Math.scala 152:17:@40694.4]
  assign x942_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40695.4]
  assign x943_x17_1_clock = clock; // @[:@40701.4]
  assign x943_x17_1_reset = reset; // @[:@40702.4]
  assign x943_x17_1_io_a = _T_2480[7:0]; // @[Math.scala 151:17:@40703.4]
  assign x943_x17_1_io_b = _T_2193[7:0]; // @[Math.scala 152:17:@40704.4]
  assign x943_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40705.4]
  assign x944_x18_1_clock = clock; // @[:@40711.4]
  assign x944_x18_1_reset = reset; // @[:@40712.4]
  assign x944_x18_1_io_a = x539_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@40713.4]
  assign x944_x18_1_io_b = _T_2484[7:0]; // @[Math.scala 152:17:@40714.4]
  assign x944_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40715.4]
  assign x945_x17_1_io_a = x941_x17_1_io_result; // @[Math.scala 151:17:@40723.4]
  assign x945_x17_1_io_b = x942_x18_1_io_result; // @[Math.scala 152:17:@40724.4]
  assign x946_x18_1_io_a = x943_x17_1_io_result; // @[Math.scala 151:17:@40733.4]
  assign x946_x18_1_io_b = x944_x18_1_io_result; // @[Math.scala 152:17:@40734.4]
  assign x947_x17_1_io_a = x945_x17_1_io_result; // @[Math.scala 151:17:@40743.4]
  assign x947_x17_1_io_b = x946_x18_1_io_result; // @[Math.scala 152:17:@40744.4]
  assign RetimeWrapper_142_clock = clock; // @[:@40751.4]
  assign RetimeWrapper_142_reset = reset; // @[:@40752.4]
  assign RetimeWrapper_142_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40754.4]
  assign RetimeWrapper_142_io_in = x539_lb_0_io_rPort_11_output_0; // @[package.scala 94:16:@40753.4]
  assign x948_sum_1_io_a = x947_x17_1_io_result; // @[Math.scala 151:17:@40762.4]
  assign x948_sum_1_io_b = RetimeWrapper_142_io_out; // @[Math.scala 152:17:@40763.4]
  assign RetimeWrapper_143_clock = clock; // @[:@40774.4]
  assign RetimeWrapper_143_reset = reset; // @[:@40775.4]
  assign RetimeWrapper_143_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@40777.4]
  assign RetimeWrapper_143_io_in = {4'h0,_T_2520}; // @[package.scala 94:16:@40776.4]
  assign RetimeWrapper_144_clock = clock; // @[:@40784.4]
  assign RetimeWrapper_144_reset = reset; // @[:@40785.4]
  assign RetimeWrapper_144_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40787.4]
  assign RetimeWrapper_144_io_in = x539_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@40786.4]
  assign x950_sub_1_io_a = RetimeWrapper_144_io_out; // @[Math.scala 192:17:@40795.4]
  assign x950_sub_1_io_b = RetimeWrapper_143_io_out; // @[Math.scala 193:17:@40796.4]
  assign RetimeWrapper_145_clock = clock; // @[:@40818.4]
  assign RetimeWrapper_145_reset = reset; // @[:@40819.4]
  assign RetimeWrapper_145_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40821.4]
  assign RetimeWrapper_145_io_in = x951 ? x950_sub_number : 8'h0; // @[package.scala 94:16:@40820.4]
  assign x954_div_1_clock = clock; // @[:@40829.4]
  assign x954_div_1_reset = reset; // @[:@40830.4]
  assign x954_div_1_io_a = RetimeWrapper_145_io_out; // @[Math.scala 328:17:@40831.4]
  assign x954_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@40833.4]
  assign RetimeWrapper_146_clock = clock; // @[:@40839.4]
  assign RetimeWrapper_146_reset = reset; // @[:@40840.4]
  assign RetimeWrapper_146_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40842.4]
  assign RetimeWrapper_146_io_in = x539_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@40841.4]
  assign x955_sum_1_io_a = RetimeWrapper_146_io_out; // @[Math.scala 151:17:@40852.4]
  assign x955_sum_1_io_b = x954_div_1_io_result; // @[Math.scala 152:17:@40853.4]
  assign RetimeWrapper_147_clock = clock; // @[:@40860.4]
  assign RetimeWrapper_147_reset = reset; // @[:@40861.4]
  assign RetimeWrapper_147_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40863.4]
  assign RetimeWrapper_147_io_in = x949_number == 8'h0; // @[package.scala 94:16:@40862.4]
  assign RetimeWrapper_148_clock = clock; // @[:@40869.4]
  assign RetimeWrapper_148_reset = reset; // @[:@40870.4]
  assign RetimeWrapper_148_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40872.4]
  assign RetimeWrapper_148_io_in = RetimeWrapper_143_io_out; // @[package.scala 94:16:@40871.4]
  assign x960_x17_1_clock = clock; // @[:@40896.4]
  assign x960_x17_1_reset = reset; // @[:@40897.4]
  assign x960_x17_1_io_a = x539_lb_0_io_rPort_23_output_0; // @[Math.scala 151:17:@40898.4]
  assign x960_x17_1_io_b = _T_2084[7:0]; // @[Math.scala 152:17:@40899.4]
  assign x960_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40900.4]
  assign x961_x18_1_clock = clock; // @[:@40906.4]
  assign x961_x18_1_reset = reset; // @[:@40907.4]
  assign x961_x18_1_io_a = x539_lb_0_io_rPort_12_output_0; // @[Math.scala 151:17:@40908.4]
  assign x961_x18_1_io_b = _T_2088[7:0]; // @[Math.scala 152:17:@40909.4]
  assign x961_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40910.4]
  assign x962_x17_1_clock = clock; // @[:@40916.4]
  assign x962_x17_1_reset = reset; // @[:@40917.4]
  assign x962_x17_1_io_a = _T_2577[7:0]; // @[Math.scala 151:17:@40918.4]
  assign x962_x17_1_io_b = _T_2581[7:0]; // @[Math.scala 152:17:@40919.4]
  assign x962_x17_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40920.4]
  assign x963_x18_1_clock = clock; // @[:@40926.4]
  assign x963_x18_1_reset = reset; // @[:@40927.4]
  assign x963_x18_1_io_a = x539_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@40928.4]
  assign x963_x18_1_io_b = _T_2585[7:0]; // @[Math.scala 152:17:@40929.4]
  assign x963_x18_1_io_flow = io_in_x527_TREADY; // @[Math.scala 153:20:@40930.4]
  assign x964_x17_1_io_a = x960_x17_1_io_result; // @[Math.scala 151:17:@40938.4]
  assign x964_x17_1_io_b = x961_x18_1_io_result; // @[Math.scala 152:17:@40939.4]
  assign x965_x18_1_io_a = x962_x17_1_io_result; // @[Math.scala 151:17:@40948.4]
  assign x965_x18_1_io_b = x963_x18_1_io_result; // @[Math.scala 152:17:@40949.4]
  assign x966_x17_1_io_a = x964_x17_1_io_result; // @[Math.scala 151:17:@40958.4]
  assign x966_x17_1_io_b = x965_x18_1_io_result; // @[Math.scala 152:17:@40959.4]
  assign RetimeWrapper_149_clock = clock; // @[:@40966.4]
  assign RetimeWrapper_149_reset = reset; // @[:@40967.4]
  assign RetimeWrapper_149_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@40969.4]
  assign RetimeWrapper_149_io_in = x539_lb_0_io_rPort_19_output_0; // @[package.scala 94:16:@40968.4]
  assign x967_sum_1_io_a = x966_x17_1_io_result; // @[Math.scala 151:17:@40977.4]
  assign x967_sum_1_io_b = RetimeWrapper_149_io_out; // @[Math.scala 152:17:@40978.4]
  assign RetimeWrapper_150_clock = clock; // @[:@40989.4]
  assign RetimeWrapper_150_reset = reset; // @[:@40990.4]
  assign RetimeWrapper_150_io_flow = io_in_x527_TREADY; // @[package.scala 95:18:@40992.4]
  assign RetimeWrapper_150_io_in = {4'h0,_T_2621}; // @[package.scala 94:16:@40991.4]
  assign RetimeWrapper_151_clock = clock; // @[:@40999.4]
  assign RetimeWrapper_151_reset = reset; // @[:@41000.4]
  assign RetimeWrapper_151_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41002.4]
  assign RetimeWrapper_151_io_in = x539_lb_0_io_rPort_23_output_0; // @[package.scala 94:16:@41001.4]
  assign x969_sub_1_io_a = RetimeWrapper_151_io_out; // @[Math.scala 192:17:@41010.4]
  assign x969_sub_1_io_b = RetimeWrapper_150_io_out; // @[Math.scala 193:17:@41011.4]
  assign RetimeWrapper_152_clock = clock; // @[:@41033.4]
  assign RetimeWrapper_152_reset = reset; // @[:@41034.4]
  assign RetimeWrapper_152_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41036.4]
  assign RetimeWrapper_152_io_in = x970 ? x969_sub_number : 8'h0; // @[package.scala 94:16:@41035.4]
  assign x973_div_1_clock = clock; // @[:@41044.4]
  assign x973_div_1_reset = reset; // @[:@41045.4]
  assign x973_div_1_io_a = RetimeWrapper_152_io_out; // @[Math.scala 328:17:@41046.4]
  assign x973_div_1_io_flow = io_in_x527_TREADY; // @[Math.scala 330:20:@41048.4]
  assign RetimeWrapper_153_clock = clock; // @[:@41054.4]
  assign RetimeWrapper_153_reset = reset; // @[:@41055.4]
  assign RetimeWrapper_153_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41057.4]
  assign RetimeWrapper_153_io_in = x539_lb_0_io_rPort_23_output_0; // @[package.scala 94:16:@41056.4]
  assign x974_sum_1_io_a = RetimeWrapper_153_io_out; // @[Math.scala 151:17:@41065.4]
  assign x974_sum_1_io_b = x973_div_1_io_result; // @[Math.scala 152:17:@41066.4]
  assign RetimeWrapper_154_clock = clock; // @[:@41073.4]
  assign RetimeWrapper_154_reset = reset; // @[:@41074.4]
  assign RetimeWrapper_154_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41076.4]
  assign RetimeWrapper_154_io_in = x968_number == 8'h0; // @[package.scala 94:16:@41075.4]
  assign RetimeWrapper_155_clock = clock; // @[:@41082.4]
  assign RetimeWrapper_155_reset = reset; // @[:@41083.4]
  assign RetimeWrapper_155_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41085.4]
  assign RetimeWrapper_155_io_in = RetimeWrapper_150_io_out; // @[package.scala 94:16:@41084.4]
  assign RetimeWrapper_156_clock = clock; // @[:@41112.4]
  assign RetimeWrapper_156_reset = reset; // @[:@41113.4]
  assign RetimeWrapper_156_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41115.4]
  assign RetimeWrapper_156_io_in = {_T_2693,_T_2690}; // @[package.scala 94:16:@41114.4]
  assign RetimeWrapper_157_clock = clock; // @[:@41121.4]
  assign RetimeWrapper_157_reset = reset; // @[:@41122.4]
  assign RetimeWrapper_157_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41124.4]
  assign RetimeWrapper_157_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@41123.4]
  assign RetimeWrapper_158_clock = clock; // @[:@41130.4]
  assign RetimeWrapper_158_reset = reset; // @[:@41131.4]
  assign RetimeWrapper_158_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41133.4]
  assign RetimeWrapper_158_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@41132.4]
  assign RetimeWrapper_159_clock = clock; // @[:@41139.4]
  assign RetimeWrapper_159_reset = reset; // @[:@41140.4]
  assign RetimeWrapper_159_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@41142.4]
  assign RetimeWrapper_159_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@41141.4]
endmodule
module x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1( // @[:@41160.2]
  input          clock, // @[:@41161.4]
  input          reset, // @[:@41162.4]
  output         io_in_x527_TVALID, // @[:@41163.4]
  input          io_in_x527_TREADY, // @[:@41163.4]
  output [255:0] io_in_x527_TDATA, // @[:@41163.4]
  input          io_in_x526_TVALID, // @[:@41163.4]
  output         io_in_x526_TREADY, // @[:@41163.4]
  input  [255:0] io_in_x526_TDATA, // @[:@41163.4]
  input  [7:0]   io_in_x526_TID, // @[:@41163.4]
  input  [7:0]   io_in_x526_TDEST, // @[:@41163.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@41163.4]
  input          io_sigsIn_smChildAcks_0, // @[:@41163.4]
  output         io_sigsOut_smDoneIn_0, // @[:@41163.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@41163.4]
  input          io_rr // @[:@41163.4]
);
  wire  x534_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x534_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x534_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x534_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire [31:0] x534_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire [31:0] x534_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x534_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x534_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x534_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@41173.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41260.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41260.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41260.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41260.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41260.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@41302.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@41302.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@41302.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@41302.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@41302.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@41310.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@41310.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TVALID; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TREADY; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire [255:0] x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TDATA; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TREADY; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire [255:0] x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TDATA; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire [7:0] x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TID; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire [7:0] x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TDEST; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire [31:0] x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire [31:0] x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
  wire  _T_239; // @[package.scala 96:25:@41265.4 package.scala 96:25:@41266.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x981_outr_UnitPipe.scala 68:66:@41271.4]
  wire  _T_252; // @[package.scala 96:25:@41307.4 package.scala 96:25:@41308.4]
  wire  _T_258; // @[package.scala 96:25:@41315.4 package.scala 96:25:@41316.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@41318.4]
  wire  x980_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@41319.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@41327.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@41328.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@41337.4]
  x534_ctrchain x534_ctrchain ( // @[SpatialBlocks.scala 37:22:@41173.4]
    .clock(x534_ctrchain_clock),
    .reset(x534_ctrchain_reset),
    .io_input_reset(x534_ctrchain_io_input_reset),
    .io_input_enable(x534_ctrchain_io_input_enable),
    .io_output_counts_1(x534_ctrchain_io_output_counts_1),
    .io_output_counts_0(x534_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x534_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x534_ctrchain_io_output_oobs_1),
    .io_output_done(x534_ctrchain_io_output_done)
  );
  x980_inr_Foreach_SAMPLER_BOX_sm x980_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 32:18:@41232.4]
    .clock(x980_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x980_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x980_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x980_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x980_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x980_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x980_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x980_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x980_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@41260.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@41302.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@41310.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1 x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1200:24:@41342.4]
    .clock(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x527_TVALID(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TVALID),
    .io_in_x527_TREADY(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TREADY),
    .io_in_x527_TDATA(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TDATA),
    .io_in_x526_TREADY(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TREADY),
    .io_in_x526_TDATA(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TDATA),
    .io_in_x526_TID(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TID),
    .io_in_x526_TDEST(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TDEST),
    .io_sigsIn_backpressure(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@41265.4 package.scala 96:25:@41266.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x526_TVALID | x980_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x981_outr_UnitPipe.scala 68:66:@41271.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@41307.4 package.scala 96:25:@41308.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@41315.4 package.scala 96:25:@41316.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@41318.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@41319.4]
  assign _T_263 = x980_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@41327.4]
  assign _T_264 = ~ x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@41328.4]
  assign _T_269 = x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@41337.4]
  assign io_in_x527_TVALID = x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TVALID; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 48:23:@41400.4]
  assign io_in_x527_TDATA = x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TDATA; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 48:23:@41398.4]
  assign io_in_x526_TREADY = x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TREADY; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 49:23:@41408.4]
  assign io_sigsOut_smDoneIn_0 = x980_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@41325.4]
  assign io_sigsOut_smCtrCopyDone_0 = x980_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@41341.4]
  assign x534_ctrchain_clock = clock; // @[:@41174.4]
  assign x534_ctrchain_reset = reset; // @[:@41175.4]
  assign x534_ctrchain_io_input_reset = x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@41340.4]
  assign x534_ctrchain_io_input_enable = _T_269 & x980_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@41295.4 SpatialBlocks.scala 130:45:@41339.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@41233.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@41234.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_io_enable = x980_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x980_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@41322.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x981_outr_UnitPipe.scala 66:50:@41268.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@41324.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x527_TREADY | x980_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@41296.4]
  assign x980_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x981_outr_UnitPipe.scala 70:48:@41274.4]
  assign RetimeWrapper_clock = clock; // @[:@41261.4]
  assign RetimeWrapper_reset = reset; // @[:@41262.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41264.4]
  assign RetimeWrapper_io_in = x534_ctrchain_io_output_done; // @[package.scala 94:16:@41263.4]
  assign RetimeWrapper_1_clock = clock; // @[:@41303.4]
  assign RetimeWrapper_1_reset = reset; // @[:@41304.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@41306.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@41305.4]
  assign RetimeWrapper_2_clock = clock; // @[:@41311.4]
  assign RetimeWrapper_2_reset = reset; // @[:@41312.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@41314.4]
  assign RetimeWrapper_2_io_in = x980_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@41313.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@41343.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@41344.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x527_TREADY = io_in_x527_TREADY; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 48:23:@41399.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TDATA = io_in_x526_TDATA; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 49:23:@41407.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TID = io_in_x526_TID; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 49:23:@41403.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x526_TDEST = io_in_x526_TDEST; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 49:23:@41402.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x527_TREADY | x980_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41426.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41424.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x980_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41422.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x534_ctrchain_io_output_counts_1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41417.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x534_ctrchain_io_output_counts_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41416.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x534_ctrchain_io_output_oobs_0; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41414.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x534_ctrchain_io_output_oobs_1; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1204:22:@41415.4]
  assign x980_inr_Foreach_SAMPLER_BOX_kernelx980_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x980_inr_Foreach_SAMPLER_BOX.scala 1203:18:@41410.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@41439.2]
  input          clock, // @[:@41440.4]
  input          reset, // @[:@41441.4]
  output         io_in_x527_TVALID, // @[:@41442.4]
  input          io_in_x527_TREADY, // @[:@41442.4]
  output [255:0] io_in_x527_TDATA, // @[:@41442.4]
  input          io_in_x526_TVALID, // @[:@41442.4]
  output         io_in_x526_TREADY, // @[:@41442.4]
  input  [255:0] io_in_x526_TDATA, // @[:@41442.4]
  input  [7:0]   io_in_x526_TID, // @[:@41442.4]
  input  [7:0]   io_in_x526_TDEST, // @[:@41442.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@41442.4]
  input          io_sigsIn_smChildAcks_0, // @[:@41442.4]
  output         io_sigsOut_smDoneIn_0, // @[:@41442.4]
  input          io_rr // @[:@41442.4]
);
  wire  x981_outr_UnitPipe_sm_clock; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_reset; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_enable; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_done; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_parentAck; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_childAck_0; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  x981_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41635.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41635.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41635.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41635.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41635.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@41643.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@41643.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@41643.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@41643.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@41643.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_clock; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_reset; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TVALID; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TREADY; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire [255:0] x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TDATA; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TVALID; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TREADY; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire [255:0] x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TDATA; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire [7:0] x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TID; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire [7:0] x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TDEST; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_rr; // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
  wire  _T_246; // @[package.scala 96:25:@41640.4 package.scala 96:25:@41641.4]
  wire  _T_252; // @[package.scala 96:25:@41648.4 package.scala 96:25:@41649.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@41651.4]
  x981_outr_UnitPipe_sm x981_outr_UnitPipe_sm ( // @[sm_x981_outr_UnitPipe.scala 32:18:@41583.4]
    .clock(x981_outr_UnitPipe_sm_clock),
    .reset(x981_outr_UnitPipe_sm_reset),
    .io_enable(x981_outr_UnitPipe_sm_io_enable),
    .io_done(x981_outr_UnitPipe_sm_io_done),
    .io_parentAck(x981_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x981_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x981_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x981_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x981_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@41635.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@41643.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1 x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1 ( // @[sm_x981_outr_UnitPipe.scala 75:24:@41670.4]
    .clock(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_clock),
    .reset(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_reset),
    .io_in_x527_TVALID(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TVALID),
    .io_in_x527_TREADY(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TREADY),
    .io_in_x527_TDATA(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TDATA),
    .io_in_x526_TVALID(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TVALID),
    .io_in_x526_TREADY(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TREADY),
    .io_in_x526_TDATA(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TDATA),
    .io_in_x526_TID(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TID),
    .io_in_x526_TDEST(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TDEST),
    .io_sigsIn_smEnableOuts_0(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@41640.4 package.scala 96:25:@41641.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@41648.4 package.scala 96:25:@41649.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@41651.4]
  assign io_in_x527_TVALID = x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TVALID; // @[sm_x981_outr_UnitPipe.scala 48:23:@41726.4]
  assign io_in_x527_TDATA = x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TDATA; // @[sm_x981_outr_UnitPipe.scala 48:23:@41724.4]
  assign io_in_x526_TREADY = x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TREADY; // @[sm_x981_outr_UnitPipe.scala 49:23:@41734.4]
  assign io_sigsOut_smDoneIn_0 = x981_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@41658.4]
  assign x981_outr_UnitPipe_sm_clock = clock; // @[:@41584.4]
  assign x981_outr_UnitPipe_sm_reset = reset; // @[:@41585.4]
  assign x981_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@41655.4]
  assign x981_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@41657.4]
  assign x981_outr_UnitPipe_sm_io_doneIn_0 = x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@41627.4]
  assign x981_outr_UnitPipe_sm_io_ctrCopyDone_0 = x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@41669.4]
  assign RetimeWrapper_clock = clock; // @[:@41636.4]
  assign RetimeWrapper_reset = reset; // @[:@41637.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41639.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@41638.4]
  assign RetimeWrapper_1_clock = clock; // @[:@41644.4]
  assign RetimeWrapper_1_reset = reset; // @[:@41645.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@41647.4]
  assign RetimeWrapper_1_io_in = x981_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@41646.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_clock = clock; // @[:@41671.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_reset = reset; // @[:@41672.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x527_TREADY = io_in_x527_TREADY; // @[sm_x981_outr_UnitPipe.scala 48:23:@41725.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TVALID = io_in_x526_TVALID; // @[sm_x981_outr_UnitPipe.scala 49:23:@41735.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TDATA = io_in_x526_TDATA; // @[sm_x981_outr_UnitPipe.scala 49:23:@41733.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TID = io_in_x526_TID; // @[sm_x981_outr_UnitPipe.scala 49:23:@41729.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_in_x526_TDEST = io_in_x526_TDEST; // @[sm_x981_outr_UnitPipe.scala 49:23:@41728.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x981_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x981_outr_UnitPipe.scala 79:22:@41744.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x981_outr_UnitPipe_sm_io_childAck_0; // @[sm_x981_outr_UnitPipe.scala 79:22:@41742.4]
  assign x981_outr_UnitPipe_kernelx981_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x981_outr_UnitPipe.scala 78:18:@41736.4]
endmodule
module AccelUnit( // @[:@41763.2]
  input          clock, // @[:@41764.4]
  input          reset, // @[:@41765.4]
  input          io_enable, // @[:@41766.4]
  output         io_done, // @[:@41766.4]
  input          io_reset, // @[:@41766.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@41766.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@41766.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@41766.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@41766.4]
  output         io_memStreams_loads_0_data_ready, // @[:@41766.4]
  input          io_memStreams_loads_0_data_valid, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@41766.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@41766.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@41766.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@41766.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@41766.4]
  input          io_memStreams_stores_0_data_ready, // @[:@41766.4]
  output         io_memStreams_stores_0_data_valid, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@41766.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@41766.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@41766.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@41766.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@41766.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@41766.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@41766.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@41766.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@41766.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@41766.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@41766.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@41766.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@41766.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@41766.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@41766.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@41766.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@41766.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@41766.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@41766.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@41766.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@41766.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@41766.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@41766.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@41766.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@41766.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@41766.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@41766.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@41766.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@41766.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@41766.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@41766.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@41766.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@41766.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@41766.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@41766.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@41766.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@41766.4]
  output         io_heap_0_req_valid, // @[:@41766.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@41766.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@41766.4]
  input          io_heap_0_resp_valid, // @[:@41766.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@41766.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@41766.4]
  input  [63:0]  io_argIns_0, // @[:@41766.4]
  input  [63:0]  io_argIns_1, // @[:@41766.4]
  input          io_argOuts_0_port_ready, // @[:@41766.4]
  output         io_argOuts_0_port_valid, // @[:@41766.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@41766.4]
  input  [63:0]  io_argOuts_0_echo // @[:@41766.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@41929.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@41929.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@41929.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@41929.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41947.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41947.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41947.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41947.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41947.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@41956.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@41956.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@41956.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@41956.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@41956.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@41956.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@41994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@42026.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@42026.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@42026.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@42026.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@42026.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_in_x527_TVALID; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_in_x527_TREADY; // @[sm_RootController.scala 73:24:@42085.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x527_TDATA; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_in_x526_TVALID; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_in_x526_TREADY; // @[sm_RootController.scala 73:24:@42085.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x526_TDATA; // @[sm_RootController.scala 73:24:@42085.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x526_TID; // @[sm_RootController.scala 73:24:@42085.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x526_TDEST; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@42085.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@42085.4]
  wire  _T_599; // @[package.scala 96:25:@41952.4 package.scala 96:25:@41953.4]
  wire  _T_664; // @[Main.scala 41:50:@42022.4]
  wire  _T_665; // @[Main.scala 41:59:@42023.4]
  wire  _T_677; // @[package.scala 100:49:@42043.4]
  reg  _T_680; // @[package.scala 48:56:@42044.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@41929.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@41947.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@41956.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@41994.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@42026.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@42085.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x527_TVALID(RootController_kernelRootController_concrete1_io_in_x527_TVALID),
    .io_in_x527_TREADY(RootController_kernelRootController_concrete1_io_in_x527_TREADY),
    .io_in_x527_TDATA(RootController_kernelRootController_concrete1_io_in_x527_TDATA),
    .io_in_x526_TVALID(RootController_kernelRootController_concrete1_io_in_x526_TVALID),
    .io_in_x526_TREADY(RootController_kernelRootController_concrete1_io_in_x526_TREADY),
    .io_in_x526_TDATA(RootController_kernelRootController_concrete1_io_in_x526_TDATA),
    .io_in_x526_TID(RootController_kernelRootController_concrete1_io_in_x526_TID),
    .io_in_x526_TDEST(RootController_kernelRootController_concrete1_io_in_x526_TDEST),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@41952.4 package.scala 96:25:@41953.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@42022.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@42023.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@42043.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@42042.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x526_TREADY; // @[sm_RootController.scala 49:23:@42149.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x527_TVALID; // @[sm_RootController.scala 48:23:@42141.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x527_TDATA; // @[sm_RootController.scala 48:23:@42139.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 48:23:@42138.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 48:23:@42137.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 48:23:@42136.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 48:23:@42135.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 48:23:@42134.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 48:23:@42133.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@41930.4]
  assign SingleCounter_reset = reset; // @[:@41931.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@41945.4]
  assign RetimeWrapper_clock = clock; // @[:@41948.4]
  assign RetimeWrapper_reset = reset; // @[:@41949.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41951.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@41950.4]
  assign SRFF_clock = clock; // @[:@41957.4]
  assign SRFF_reset = reset; // @[:@41958.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@42177.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@42040.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@42041.4]
  assign RootController_sm_clock = clock; // @[:@41995.4]
  assign RootController_sm_reset = reset; // @[:@41996.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@42039.4 SpatialBlocks.scala 112:18:@42073.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@42067.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@42047.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@42064.4]
  assign RetimeWrapper_1_clock = clock; // @[:@42027.4]
  assign RetimeWrapper_1_reset = reset; // @[:@42028.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@42030.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@42029.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@42086.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@42087.4]
  assign RootController_kernelRootController_concrete1_io_in_x527_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 48:23:@42140.4]
  assign RootController_kernelRootController_concrete1_io_in_x526_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 49:23:@42150.4]
  assign RootController_kernelRootController_concrete1_io_in_x526_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 49:23:@42148.4]
  assign RootController_kernelRootController_concrete1_io_in_x526_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 49:23:@42144.4]
  assign RootController_kernelRootController_concrete1_io_in_x526_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 49:23:@42143.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@42159.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@42157.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@42151.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@42179.2]
  input         clock, // @[:@42180.4]
  input         reset, // @[:@42181.4]
  input  [31:0] io_raddr, // @[:@42182.4]
  input         io_wen, // @[:@42182.4]
  input  [31:0] io_waddr, // @[:@42182.4]
  input  [63:0] io_wdata, // @[:@42182.4]
  output [63:0] io_rdata // @[:@42182.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@42184.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@42184.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@42184.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@42184.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@42184.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@42184.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@42184.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@42184.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@42184.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@42184.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@42184.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@42184.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@42185.4]
  assign accel_reset = reset; // @[:@42186.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
