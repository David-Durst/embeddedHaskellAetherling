module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module atomTupleCreator_t0Int_t1Int (input [7:0] I0/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O__0/*verilator public*/, output [7:0] O__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O__0 = I0;
assign O__1 = I1;
assign valid_down = valid_up;
endmodule

module coreir_ult #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 < in1;
endmodule

module coreir_term #(parameter width = 1) (input [width-1:0] in/*verilator public*/);

endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_mux #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, input sel/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = sel ? in1 : in0;
endmodule

module coreir_eq #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 == in1;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out/*verilator public*/);
  assign out = value;
endmodule

module coreir_add #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 + in1;
endmodule

module \commonlib_muxn__N2__width1 (input [0:0] in_data_0/*verilator public*/, input [0:0] in_data_1/*verilator public*/, input [0:0] in_sel/*verilator public*/, output [0:0] out/*verilator public*/);
wire [0:0] _join_out;
coreir_mux #(.width(1)) _join(.in0(in_data_0), .in1(in_data_1), .out(_join_out), .sel(in_sel[0]));
assign out = _join_out;
endmodule

module lutN #(parameter N = 1, parameter init = 1) (input [N-1:0] in/*verilator public*/, output out/*verilator public*/);
  assign out = init[in];
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit8 (input [7:0] in/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit (input in/*verilator public*/, output [0:0] out/*verilator public*/);
assign out = in;
endmodule

module Term_Bitt (input I/*verilator public*/);
wire [0:0] dehydrate_tBit_inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBit_inst0_out));
endmodule

module SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] const_0_1_out;
Term_Bitt Term_Bitt_inst0(.I(CE));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
assign O = const_0_1_out;
endmodule

module Mux2xOutBits1 (input [0:0] I0/*verilator public*/, input [0:0] I1/*verilator public*/, output [0:0] O/*verilator public*/, input S/*verilator public*/);
wire [0:0] coreir_commonlib_mux2x1_inst0_out;
\commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(.in_data_0(I0), .in_data_1(I1), .in_sel(S), .out(coreir_commonlib_mux2x1_inst0_out));
assign O = coreir_commonlib_mux2x1_inst0_out;
endmodule

module Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1 (input CE/*verilator public*/, input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [0:0] Mux2xOutBits1_inst0_O;
wire [0:0] const_0_1_out;
wire [0:0] enable_mux_O;
wire [0:0] value_out;
Mux2xOutBits1 Mux2xOutBits1_inst0(.I0(enable_mux_O), .I1(const_0_1_out), .O(Mux2xOutBits1_inst0_O), .S(RESET));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
Mux2xOutBits1 enable_mux(.I0(value_out), .I1(I), .O(enable_mux_O), .S(CE));
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) value(.clk(CLK), .in(Mux2xOutBits1_inst0_O), .out(value_out));
assign O = value_out;
endmodule

module LUT1_2 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h2), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_1 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h1), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_0 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h0), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT_Array_8_Bit_t_1n (input CLK/*verilator public*/, input [0:0] addr/*verilator public*/, output [7:0] data/*verilator public*/);
wire LUT1_0_inst0_O;
wire LUT1_0_inst1_O;
wire LUT1_0_inst2_O;
wire LUT1_0_inst3_O;
wire LUT1_0_inst4_O;
wire LUT1_0_inst5_O;
wire LUT1_1_inst0_O;
wire LUT1_1_inst1_O;
wire [7:0] hydrate_tArray_8_Bit__inst0_out;
LUT1_0 LUT1_0_inst0(.I0(addr[0]), .O(LUT1_0_inst0_O));
LUT1_0 LUT1_0_inst1(.I0(addr[0]), .O(LUT1_0_inst1_O));
LUT1_0 LUT1_0_inst2(.I0(addr[0]), .O(LUT1_0_inst2_O));
LUT1_0 LUT1_0_inst3(.I0(addr[0]), .O(LUT1_0_inst3_O));
LUT1_0 LUT1_0_inst4(.I0(addr[0]), .O(LUT1_0_inst4_O));
LUT1_0 LUT1_0_inst5(.I0(addr[0]), .O(LUT1_0_inst5_O));
LUT1_1 LUT1_1_inst0(.I0(addr[0]), .O(LUT1_1_inst0_O));
LUT1_1 LUT1_1_inst1(.I0(addr[0]), .O(LUT1_1_inst1_O));
\aetherlinglib_hydrate__hydratedTypeBit8 hydrate_tArray_8_Bit__inst0(.in({LUT1_0_inst5_O,LUT1_0_inst4_O,LUT1_0_inst3_O,LUT1_0_inst2_O,LUT1_0_inst1_O,LUT1_1_inst1_O,LUT1_0_inst0_O,LUT1_1_inst0_O}), .out(hydrate_tArray_8_Bit__inst0_out));
assign data = hydrate_tArray_8_Bit__inst0_out;
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Bit_t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8_inst0_O;
Register8 Register8_inst0(.CLK(CLK), .I(I), .O(Register8_inst0_O));
assign O = Register8_inst0_O;
endmodule

module Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst100_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst101_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst102_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst103_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst104_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst105_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst106_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst107_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst108_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst109_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst110_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst111_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst112_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst113_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst114_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst115_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst116_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst117_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst118_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst119_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst120_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst121_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst122_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst123_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst124_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst125_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst126_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst127_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst128_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst129_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst130_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst131_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst132_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst133_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst134_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst135_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst136_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst137_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst138_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst139_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst140_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst141_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst142_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst143_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst144_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst145_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst146_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst147_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst148_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst149_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst150_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst151_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst152_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst153_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst154_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst155_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst156_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst157_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst158_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst159_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst160_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst161_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst162_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst163_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst164_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst165_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst166_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst167_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst168_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst169_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst170_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst171_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst172_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst173_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst174_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst175_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst176_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst177_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst178_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst179_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst180_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst181_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst182_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst183_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst184_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst185_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst186_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst187_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst188_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst189_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst190_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst191_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst192_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst193_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst194_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst195_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst196_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst197_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst198_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst199_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst20_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst21_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst22_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst23_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst24_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst25_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst26_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst27_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst28_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst29_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst30_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst31_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst32_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst33_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst34_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst35_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst36_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst37_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst38_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst39_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst40_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst41_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst42_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst43_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst44_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst45_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst46_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst47_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst48_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst49_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst50_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst51_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst52_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst53_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst54_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst55_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst56_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst57_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst58_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst59_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst60_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst61_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst62_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst63_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst64_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst65_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst66_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst67_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst68_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst69_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst70_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst71_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst72_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst73_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst74_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst75_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst76_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst77_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst78_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst79_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst80_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst81_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst82_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst83_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst84_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst85_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst86_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst87_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst88_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst89_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst90_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst91_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst92_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst93_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst94_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst95_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst96_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst97_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst98_O;
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst99_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I_0), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1(.CLK(CLK), .I(I_1), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10(.CLK(CLK), .I(I_10), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst100(.CLK(CLK), .I(I_100), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst100_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst101(.CLK(CLK), .I(I_101), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst101_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst102(.CLK(CLK), .I(I_102), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst102_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst103(.CLK(CLK), .I(I_103), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst103_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst104(.CLK(CLK), .I(I_104), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst104_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst105(.CLK(CLK), .I(I_105), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst105_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst106(.CLK(CLK), .I(I_106), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst106_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst107(.CLK(CLK), .I(I_107), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst107_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst108(.CLK(CLK), .I(I_108), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst108_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst109(.CLK(CLK), .I(I_109), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst109_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11(.CLK(CLK), .I(I_11), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst110(.CLK(CLK), .I(I_110), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst110_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst111(.CLK(CLK), .I(I_111), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst111_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst112(.CLK(CLK), .I(I_112), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst112_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst113(.CLK(CLK), .I(I_113), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst113_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst114(.CLK(CLK), .I(I_114), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst114_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst115(.CLK(CLK), .I(I_115), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst115_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst116(.CLK(CLK), .I(I_116), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst116_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst117(.CLK(CLK), .I(I_117), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst117_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst118(.CLK(CLK), .I(I_118), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst118_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst119(.CLK(CLK), .I(I_119), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst119_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12(.CLK(CLK), .I(I_12), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst120(.CLK(CLK), .I(I_120), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst120_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst121(.CLK(CLK), .I(I_121), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst121_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst122(.CLK(CLK), .I(I_122), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst122_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst123(.CLK(CLK), .I(I_123), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst123_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst124(.CLK(CLK), .I(I_124), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst124_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst125(.CLK(CLK), .I(I_125), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst125_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst126(.CLK(CLK), .I(I_126), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst126_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst127(.CLK(CLK), .I(I_127), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst127_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst128(.CLK(CLK), .I(I_128), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst128_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst129(.CLK(CLK), .I(I_129), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst129_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13(.CLK(CLK), .I(I_13), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst130(.CLK(CLK), .I(I_130), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst130_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst131(.CLK(CLK), .I(I_131), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst131_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst132(.CLK(CLK), .I(I_132), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst132_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst133(.CLK(CLK), .I(I_133), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst133_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst134(.CLK(CLK), .I(I_134), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst134_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst135(.CLK(CLK), .I(I_135), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst135_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst136(.CLK(CLK), .I(I_136), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst136_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst137(.CLK(CLK), .I(I_137), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst137_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst138(.CLK(CLK), .I(I_138), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst138_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst139(.CLK(CLK), .I(I_139), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst139_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14(.CLK(CLK), .I(I_14), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst140(.CLK(CLK), .I(I_140), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst140_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst141(.CLK(CLK), .I(I_141), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst141_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst142(.CLK(CLK), .I(I_142), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst142_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst143(.CLK(CLK), .I(I_143), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst143_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst144(.CLK(CLK), .I(I_144), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst144_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst145(.CLK(CLK), .I(I_145), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst145_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst146(.CLK(CLK), .I(I_146), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst146_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst147(.CLK(CLK), .I(I_147), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst147_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst148(.CLK(CLK), .I(I_148), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst148_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst149(.CLK(CLK), .I(I_149), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst149_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15(.CLK(CLK), .I(I_15), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst150(.CLK(CLK), .I(I_150), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst150_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst151(.CLK(CLK), .I(I_151), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst151_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst152(.CLK(CLK), .I(I_152), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst152_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst153(.CLK(CLK), .I(I_153), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst153_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst154(.CLK(CLK), .I(I_154), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst154_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst155(.CLK(CLK), .I(I_155), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst155_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst156(.CLK(CLK), .I(I_156), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst156_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst157(.CLK(CLK), .I(I_157), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst157_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst158(.CLK(CLK), .I(I_158), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst158_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst159(.CLK(CLK), .I(I_159), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst159_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16(.CLK(CLK), .I(I_16), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst160(.CLK(CLK), .I(I_160), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst160_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst161(.CLK(CLK), .I(I_161), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst161_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst162(.CLK(CLK), .I(I_162), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst162_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst163(.CLK(CLK), .I(I_163), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst163_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst164(.CLK(CLK), .I(I_164), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst164_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst165(.CLK(CLK), .I(I_165), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst165_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst166(.CLK(CLK), .I(I_166), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst166_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst167(.CLK(CLK), .I(I_167), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst167_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst168(.CLK(CLK), .I(I_168), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst168_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst169(.CLK(CLK), .I(I_169), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst169_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17(.CLK(CLK), .I(I_17), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst170(.CLK(CLK), .I(I_170), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst170_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst171(.CLK(CLK), .I(I_171), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst171_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst172(.CLK(CLK), .I(I_172), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst172_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst173(.CLK(CLK), .I(I_173), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst173_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst174(.CLK(CLK), .I(I_174), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst174_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst175(.CLK(CLK), .I(I_175), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst175_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst176(.CLK(CLK), .I(I_176), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst176_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst177(.CLK(CLK), .I(I_177), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst177_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst178(.CLK(CLK), .I(I_178), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst178_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst179(.CLK(CLK), .I(I_179), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst179_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18(.CLK(CLK), .I(I_18), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst180(.CLK(CLK), .I(I_180), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst180_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst181(.CLK(CLK), .I(I_181), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst181_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst182(.CLK(CLK), .I(I_182), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst182_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst183(.CLK(CLK), .I(I_183), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst183_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst184(.CLK(CLK), .I(I_184), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst184_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst185(.CLK(CLK), .I(I_185), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst185_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst186(.CLK(CLK), .I(I_186), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst186_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst187(.CLK(CLK), .I(I_187), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst187_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst188(.CLK(CLK), .I(I_188), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst188_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst189(.CLK(CLK), .I(I_189), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst189_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19(.CLK(CLK), .I(I_19), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst190(.CLK(CLK), .I(I_190), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst190_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst191(.CLK(CLK), .I(I_191), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst191_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst192(.CLK(CLK), .I(I_192), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst192_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst193(.CLK(CLK), .I(I_193), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst193_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst194(.CLK(CLK), .I(I_194), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst194_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst195(.CLK(CLK), .I(I_195), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst195_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst196(.CLK(CLK), .I(I_196), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst196_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst197(.CLK(CLK), .I(I_197), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst197_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst198(.CLK(CLK), .I(I_198), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst198_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst199(.CLK(CLK), .I(I_199), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst199_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2(.CLK(CLK), .I(I_2), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst20(.CLK(CLK), .I(I_20), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst20_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst21(.CLK(CLK), .I(I_21), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst21_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst22(.CLK(CLK), .I(I_22), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst22_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst23(.CLK(CLK), .I(I_23), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst23_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst24(.CLK(CLK), .I(I_24), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst24_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst25(.CLK(CLK), .I(I_25), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst25_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst26(.CLK(CLK), .I(I_26), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst26_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst27(.CLK(CLK), .I(I_27), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst27_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst28(.CLK(CLK), .I(I_28), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst28_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst29(.CLK(CLK), .I(I_29), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst29_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3(.CLK(CLK), .I(I_3), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst30(.CLK(CLK), .I(I_30), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst30_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst31(.CLK(CLK), .I(I_31), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst31_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst32(.CLK(CLK), .I(I_32), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst32_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst33(.CLK(CLK), .I(I_33), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst33_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst34(.CLK(CLK), .I(I_34), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst34_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst35(.CLK(CLK), .I(I_35), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst35_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst36(.CLK(CLK), .I(I_36), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst36_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst37(.CLK(CLK), .I(I_37), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst37_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst38(.CLK(CLK), .I(I_38), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst38_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst39(.CLK(CLK), .I(I_39), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst39_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4(.CLK(CLK), .I(I_4), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst40(.CLK(CLK), .I(I_40), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst40_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst41(.CLK(CLK), .I(I_41), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst41_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst42(.CLK(CLK), .I(I_42), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst42_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst43(.CLK(CLK), .I(I_43), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst43_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst44(.CLK(CLK), .I(I_44), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst44_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst45(.CLK(CLK), .I(I_45), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst45_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst46(.CLK(CLK), .I(I_46), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst46_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst47(.CLK(CLK), .I(I_47), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst47_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst48(.CLK(CLK), .I(I_48), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst48_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst49(.CLK(CLK), .I(I_49), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst49_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5(.CLK(CLK), .I(I_5), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst50(.CLK(CLK), .I(I_50), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst50_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst51(.CLK(CLK), .I(I_51), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst51_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst52(.CLK(CLK), .I(I_52), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst52_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst53(.CLK(CLK), .I(I_53), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst53_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst54(.CLK(CLK), .I(I_54), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst54_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst55(.CLK(CLK), .I(I_55), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst55_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst56(.CLK(CLK), .I(I_56), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst56_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst57(.CLK(CLK), .I(I_57), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst57_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst58(.CLK(CLK), .I(I_58), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst58_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst59(.CLK(CLK), .I(I_59), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst59_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6(.CLK(CLK), .I(I_6), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst60(.CLK(CLK), .I(I_60), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst60_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst61(.CLK(CLK), .I(I_61), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst61_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst62(.CLK(CLK), .I(I_62), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst62_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst63(.CLK(CLK), .I(I_63), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst63_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst64(.CLK(CLK), .I(I_64), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst64_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst65(.CLK(CLK), .I(I_65), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst65_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst66(.CLK(CLK), .I(I_66), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst66_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst67(.CLK(CLK), .I(I_67), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst67_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst68(.CLK(CLK), .I(I_68), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst68_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst69(.CLK(CLK), .I(I_69), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst69_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7(.CLK(CLK), .I(I_7), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst70(.CLK(CLK), .I(I_70), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst70_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst71(.CLK(CLK), .I(I_71), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst71_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst72(.CLK(CLK), .I(I_72), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst72_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst73(.CLK(CLK), .I(I_73), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst73_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst74(.CLK(CLK), .I(I_74), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst74_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst75(.CLK(CLK), .I(I_75), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst75_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst76(.CLK(CLK), .I(I_76), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst76_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst77(.CLK(CLK), .I(I_77), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst77_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst78(.CLK(CLK), .I(I_78), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst78_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst79(.CLK(CLK), .I(I_79), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst79_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8(.CLK(CLK), .I(I_8), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst80(.CLK(CLK), .I(I_80), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst80_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst81(.CLK(CLK), .I(I_81), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst81_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst82(.CLK(CLK), .I(I_82), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst82_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst83(.CLK(CLK), .I(I_83), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst83_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst84(.CLK(CLK), .I(I_84), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst84_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst85(.CLK(CLK), .I(I_85), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst85_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst86(.CLK(CLK), .I(I_86), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst86_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst87(.CLK(CLK), .I(I_87), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst87_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst88(.CLK(CLK), .I(I_88), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst88_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst89(.CLK(CLK), .I(I_89), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst89_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9(.CLK(CLK), .I(I_9), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst90(.CLK(CLK), .I(I_90), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst90_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst91(.CLK(CLK), .I(I_91), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst91_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst92(.CLK(CLK), .I(I_92), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst92_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst93(.CLK(CLK), .I(I_93), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst93_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst94(.CLK(CLK), .I(I_94), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst94_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst95(.CLK(CLK), .I(I_95), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst95_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst96(.CLK(CLK), .I(I_96), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst96_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst97(.CLK(CLK), .I(I_97), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst97_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst98(.CLK(CLK), .I(I_98), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst98_O));
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst99(.CLK(CLK), .I(I_99), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst99_O));
assign O_0 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
assign O_1 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst1_O;
assign O_10 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst10_O;
assign O_100 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst100_O;
assign O_101 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst101_O;
assign O_102 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst102_O;
assign O_103 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst103_O;
assign O_104 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst104_O;
assign O_105 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst105_O;
assign O_106 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst106_O;
assign O_107 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst107_O;
assign O_108 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst108_O;
assign O_109 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst109_O;
assign O_11 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst11_O;
assign O_110 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst110_O;
assign O_111 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst111_O;
assign O_112 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst112_O;
assign O_113 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst113_O;
assign O_114 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst114_O;
assign O_115 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst115_O;
assign O_116 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst116_O;
assign O_117 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst117_O;
assign O_118 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst118_O;
assign O_119 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst119_O;
assign O_12 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst12_O;
assign O_120 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst120_O;
assign O_121 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst121_O;
assign O_122 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst122_O;
assign O_123 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst123_O;
assign O_124 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst124_O;
assign O_125 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst125_O;
assign O_126 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst126_O;
assign O_127 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst127_O;
assign O_128 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst128_O;
assign O_129 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst129_O;
assign O_13 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst13_O;
assign O_130 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst130_O;
assign O_131 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst131_O;
assign O_132 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst132_O;
assign O_133 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst133_O;
assign O_134 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst134_O;
assign O_135 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst135_O;
assign O_136 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst136_O;
assign O_137 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst137_O;
assign O_138 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst138_O;
assign O_139 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst139_O;
assign O_14 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst14_O;
assign O_140 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst140_O;
assign O_141 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst141_O;
assign O_142 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst142_O;
assign O_143 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst143_O;
assign O_144 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst144_O;
assign O_145 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst145_O;
assign O_146 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst146_O;
assign O_147 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst147_O;
assign O_148 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst148_O;
assign O_149 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst149_O;
assign O_15 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst15_O;
assign O_150 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst150_O;
assign O_151 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst151_O;
assign O_152 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst152_O;
assign O_153 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst153_O;
assign O_154 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst154_O;
assign O_155 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst155_O;
assign O_156 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst156_O;
assign O_157 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst157_O;
assign O_158 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst158_O;
assign O_159 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst159_O;
assign O_16 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst16_O;
assign O_160 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst160_O;
assign O_161 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst161_O;
assign O_162 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst162_O;
assign O_163 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst163_O;
assign O_164 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst164_O;
assign O_165 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst165_O;
assign O_166 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst166_O;
assign O_167 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst167_O;
assign O_168 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst168_O;
assign O_169 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst169_O;
assign O_17 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst17_O;
assign O_170 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst170_O;
assign O_171 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst171_O;
assign O_172 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst172_O;
assign O_173 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst173_O;
assign O_174 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst174_O;
assign O_175 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst175_O;
assign O_176 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst176_O;
assign O_177 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst177_O;
assign O_178 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst178_O;
assign O_179 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst179_O;
assign O_18 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst18_O;
assign O_180 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst180_O;
assign O_181 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst181_O;
assign O_182 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst182_O;
assign O_183 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst183_O;
assign O_184 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst184_O;
assign O_185 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst185_O;
assign O_186 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst186_O;
assign O_187 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst187_O;
assign O_188 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst188_O;
assign O_189 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst189_O;
assign O_19 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst19_O;
assign O_190 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst190_O;
assign O_191 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst191_O;
assign O_192 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst192_O;
assign O_193 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst193_O;
assign O_194 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst194_O;
assign O_195 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst195_O;
assign O_196 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst196_O;
assign O_197 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst197_O;
assign O_198 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst198_O;
assign O_199 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst199_O;
assign O_2 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst2_O;
assign O_20 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst20_O;
assign O_21 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst21_O;
assign O_22 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst22_O;
assign O_23 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst23_O;
assign O_24 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst24_O;
assign O_25 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst25_O;
assign O_26 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst26_O;
assign O_27 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst27_O;
assign O_28 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst28_O;
assign O_29 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst29_O;
assign O_3 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst3_O;
assign O_30 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst30_O;
assign O_31 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst31_O;
assign O_32 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst32_O;
assign O_33 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst33_O;
assign O_34 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst34_O;
assign O_35 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst35_O;
assign O_36 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst36_O;
assign O_37 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst37_O;
assign O_38 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst38_O;
assign O_39 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst39_O;
assign O_4 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst4_O;
assign O_40 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst40_O;
assign O_41 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst41_O;
assign O_42 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst42_O;
assign O_43 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst43_O;
assign O_44 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst44_O;
assign O_45 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst45_O;
assign O_46 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst46_O;
assign O_47 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst47_O;
assign O_48 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst48_O;
assign O_49 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst49_O;
assign O_5 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst5_O;
assign O_50 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst50_O;
assign O_51 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst51_O;
assign O_52 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst52_O;
assign O_53 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst53_O;
assign O_54 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst54_O;
assign O_55 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst55_O;
assign O_56 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst56_O;
assign O_57 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst57_O;
assign O_58 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst58_O;
assign O_59 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst59_O;
assign O_6 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst6_O;
assign O_60 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst60_O;
assign O_61 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst61_O;
assign O_62 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst62_O;
assign O_63 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst63_O;
assign O_64 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst64_O;
assign O_65 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst65_O;
assign O_66 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst66_O;
assign O_67 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst67_O;
assign O_68 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst68_O;
assign O_69 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst69_O;
assign O_7 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst7_O;
assign O_70 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst70_O;
assign O_71 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst71_O;
assign O_72 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst72_O;
assign O_73 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst73_O;
assign O_74 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst74_O;
assign O_75 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst75_O;
assign O_76 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst76_O;
assign O_77 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst77_O;
assign O_78 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst78_O;
assign O_79 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst79_O;
assign O_8 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst8_O;
assign O_80 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst80_O;
assign O_81 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst81_O;
assign O_82 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst82_O;
assign O_83 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst83_O;
assign O_84 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst84_O;
assign O_85 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst85_O;
assign O_86 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst86_O;
assign O_87 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst87_O;
assign O_88 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst88_O;
assign O_89 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst89_O;
assign O_9 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst9_O;
assign O_90 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst90_O;
assign O_91 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst91_O;
assign O_92 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst92_O;
assign O_93 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst93_O;
assign O_94 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst94_O;
assign O_95 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst95_O;
assign O_96 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst96_O;
assign O_97 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst97_O;
assign O_98 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst98_O;
assign O_99 = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst99_O;
endmodule

module Register1 (input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
assign O = DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
endmodule

module Register_Bitt_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] Register1_inst0_O;
Register1 Register1_inst0(.CLK(CLK), .I(I), .O(Register1_inst0_O));
assign O = Register1_inst0_O[0];
endmodule

module FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_100;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_101;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_102;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_103;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_104;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_105;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_106;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_107;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_108;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_109;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_110;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_111;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_112;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_113;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_114;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_115;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_116;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_117;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_118;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_119;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_120;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_121;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_122;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_123;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_124;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_125;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_126;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_127;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_128;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_129;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_130;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_131;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_132;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_133;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_134;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_135;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_136;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_137;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_138;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_139;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_140;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_141;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_142;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_143;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_144;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_145;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_146;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_147;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_148;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_149;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_150;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_151;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_152;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_153;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_154;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_155;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_156;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_157;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_158;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_159;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_160;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_161;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_162;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_163;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_164;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_165;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_166;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_167;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_168;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_169;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_170;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_171;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_172;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_173;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_174;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_175;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_176;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_177;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_178;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_179;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_180;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_181;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_182;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_183;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_184;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_185;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_186;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_187;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_188;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_189;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_190;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_191;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_192;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_193;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_194;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_195;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_196;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_197;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_198;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_199;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_40;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_41;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_42;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_43;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_44;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_45;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_46;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_47;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_48;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_49;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_50;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_51;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_52;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_53;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_54;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_55;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_56;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_57;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_58;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_59;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_60;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_61;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_62;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_63;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_64;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_65;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_66;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_67;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_68;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_69;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_70;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_71;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_72;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_73;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_74;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_75;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_76;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_77;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_78;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_79;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_80;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_81;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_82;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_83;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_84;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_85;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_86;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_87;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_88;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_89;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_90;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_91;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_92;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_93;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_94;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_95;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_96;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_97;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_98;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_99;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_100(I_100), .I_101(I_101), .I_102(I_102), .I_103(I_103), .I_104(I_104), .I_105(I_105), .I_106(I_106), .I_107(I_107), .I_108(I_108), .I_109(I_109), .I_11(I_11), .I_110(I_110), .I_111(I_111), .I_112(I_112), .I_113(I_113), .I_114(I_114), .I_115(I_115), .I_116(I_116), .I_117(I_117), .I_118(I_118), .I_119(I_119), .I_12(I_12), .I_120(I_120), .I_121(I_121), .I_122(I_122), .I_123(I_123), .I_124(I_124), .I_125(I_125), .I_126(I_126), .I_127(I_127), .I_128(I_128), .I_129(I_129), .I_13(I_13), .I_130(I_130), .I_131(I_131), .I_132(I_132), .I_133(I_133), .I_134(I_134), .I_135(I_135), .I_136(I_136), .I_137(I_137), .I_138(I_138), .I_139(I_139), .I_14(I_14), .I_140(I_140), .I_141(I_141), .I_142(I_142), .I_143(I_143), .I_144(I_144), .I_145(I_145), .I_146(I_146), .I_147(I_147), .I_148(I_148), .I_149(I_149), .I_15(I_15), .I_150(I_150), .I_151(I_151), .I_152(I_152), .I_153(I_153), .I_154(I_154), .I_155(I_155), .I_156(I_156), .I_157(I_157), .I_158(I_158), .I_159(I_159), .I_16(I_16), .I_160(I_160), .I_161(I_161), .I_162(I_162), .I_163(I_163), .I_164(I_164), .I_165(I_165), .I_166(I_166), .I_167(I_167), .I_168(I_168), .I_169(I_169), .I_17(I_17), .I_170(I_170), .I_171(I_171), .I_172(I_172), .I_173(I_173), .I_174(I_174), .I_175(I_175), .I_176(I_176), .I_177(I_177), .I_178(I_178), .I_179(I_179), .I_18(I_18), .I_180(I_180), .I_181(I_181), .I_182(I_182), .I_183(I_183), .I_184(I_184), .I_185(I_185), .I_186(I_186), .I_187(I_187), .I_188(I_188), .I_189(I_189), .I_19(I_19), .I_190(I_190), .I_191(I_191), .I_192(I_192), .I_193(I_193), .I_194(I_194), .I_195(I_195), .I_196(I_196), .I_197(I_197), .I_198(I_198), .I_199(I_199), .I_2(I_2), .I_20(I_20), .I_21(I_21), .I_22(I_22), .I_23(I_23), .I_24(I_24), .I_25(I_25), .I_26(I_26), .I_27(I_27), .I_28(I_28), .I_29(I_29), .I_3(I_3), .I_30(I_30), .I_31(I_31), .I_32(I_32), .I_33(I_33), .I_34(I_34), .I_35(I_35), .I_36(I_36), .I_37(I_37), .I_38(I_38), .I_39(I_39), .I_4(I_4), .I_40(I_40), .I_41(I_41), .I_42(I_42), .I_43(I_43), .I_44(I_44), .I_45(I_45), .I_46(I_46), .I_47(I_47), .I_48(I_48), .I_49(I_49), .I_5(I_5), .I_50(I_50), .I_51(I_51), .I_52(I_52), .I_53(I_53), .I_54(I_54), .I_55(I_55), .I_56(I_56), .I_57(I_57), .I_58(I_58), .I_59(I_59), .I_6(I_6), .I_60(I_60), .I_61(I_61), .I_62(I_62), .I_63(I_63), .I_64(I_64), .I_65(I_65), .I_66(I_66), .I_67(I_67), .I_68(I_68), .I_69(I_69), .I_7(I_7), .I_70(I_70), .I_71(I_71), .I_72(I_72), .I_73(I_73), .I_74(I_74), .I_75(I_75), .I_76(I_76), .I_77(I_77), .I_78(I_78), .I_79(I_79), .I_8(I_8), .I_80(I_80), .I_81(I_81), .I_82(I_82), .I_83(I_83), .I_84(I_84), .I_85(I_85), .I_86(I_86), .I_87(I_87), .I_88(I_88), .I_89(I_89), .I_9(I_9), .I_90(I_90), .I_91(I_91), .I_92(I_92), .I_93(I_93), .I_94(I_94), .I_95(I_95), .I_96(I_96), .I_97(I_97), .I_98(I_98), .I_99(I_99), .O_0(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0), .O_1(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1), .O_10(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10), .O_100(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_100), .O_101(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_101), .O_102(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_102), .O_103(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_103), .O_104(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_104), .O_105(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_105), .O_106(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_106), .O_107(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_107), .O_108(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_108), .O_109(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_109), .O_11(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11), .O_110(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_110), .O_111(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_111), .O_112(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_112), .O_113(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_113), .O_114(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_114), .O_115(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_115), .O_116(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_116), .O_117(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_117), .O_118(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_118), .O_119(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_119), .O_12(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12), .O_120(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_120), .O_121(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_121), .O_122(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_122), .O_123(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_123), .O_124(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_124), .O_125(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_125), .O_126(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_126), .O_127(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_127), .O_128(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_128), .O_129(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_129), .O_13(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13), .O_130(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_130), .O_131(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_131), .O_132(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_132), .O_133(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_133), .O_134(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_134), .O_135(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_135), .O_136(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_136), .O_137(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_137), .O_138(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_138), .O_139(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_139), .O_14(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14), .O_140(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_140), .O_141(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_141), .O_142(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_142), .O_143(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_143), .O_144(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_144), .O_145(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_145), .O_146(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_146), .O_147(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_147), .O_148(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_148), .O_149(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_149), .O_15(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15), .O_150(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_150), .O_151(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_151), .O_152(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_152), .O_153(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_153), .O_154(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_154), .O_155(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_155), .O_156(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_156), .O_157(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_157), .O_158(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_158), .O_159(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_159), .O_16(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16), .O_160(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_160), .O_161(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_161), .O_162(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_162), .O_163(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_163), .O_164(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_164), .O_165(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_165), .O_166(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_166), .O_167(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_167), .O_168(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_168), .O_169(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_169), .O_17(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17), .O_170(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_170), .O_171(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_171), .O_172(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_172), .O_173(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_173), .O_174(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_174), .O_175(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_175), .O_176(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_176), .O_177(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_177), .O_178(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_178), .O_179(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_179), .O_18(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18), .O_180(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_180), .O_181(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_181), .O_182(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_182), .O_183(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_183), .O_184(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_184), .O_185(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_185), .O_186(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_186), .O_187(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_187), .O_188(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_188), .O_189(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_189), .O_19(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19), .O_190(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_190), .O_191(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_191), .O_192(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_192), .O_193(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_193), .O_194(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_194), .O_195(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_195), .O_196(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_196), .O_197(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_197), .O_198(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_198), .O_199(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_199), .O_2(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2), .O_20(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20), .O_21(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21), .O_22(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22), .O_23(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23), .O_24(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24), .O_25(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25), .O_26(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26), .O_27(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27), .O_28(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28), .O_29(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29), .O_3(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3), .O_30(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30), .O_31(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31), .O_32(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32), .O_33(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33), .O_34(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34), .O_35(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35), .O_36(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36), .O_37(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37), .O_38(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38), .O_39(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39), .O_4(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4), .O_40(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_40), .O_41(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_41), .O_42(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_42), .O_43(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_43), .O_44(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_44), .O_45(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_45), .O_46(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_46), .O_47(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_47), .O_48(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_48), .O_49(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_49), .O_5(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5), .O_50(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_50), .O_51(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_51), .O_52(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_52), .O_53(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_53), .O_54(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_54), .O_55(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_55), .O_56(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_56), .O_57(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_57), .O_58(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_58), .O_59(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_59), .O_6(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6), .O_60(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_60), .O_61(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_61), .O_62(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_62), .O_63(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_63), .O_64(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_64), .O_65(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_65), .O_66(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_66), .O_67(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_67), .O_68(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_68), .O_69(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_69), .O_7(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7), .O_70(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_70), .O_71(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_71), .O_72(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_72), .O_73(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_73), .O_74(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_74), .O_75(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_75), .O_76(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_76), .O_77(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_77), .O_78(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_78), .O_79(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_79), .O_8(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8), .O_80(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_80), .O_81(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_81), .O_82(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_82), .O_83(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_83), .O_84(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_84), .O_85(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_85), .O_86(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_86), .O_87(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_87), .O_88(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_88), .O_89(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_89), .O_9(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9), .O_90(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_90), .O_91(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_91), .O_92(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_92), .O_93(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_93), .O_94(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_94), .O_95(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_95), .O_96(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_96), .O_97(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_97), .O_98(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_98), .O_99(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_99));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_1 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
assign O_10 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
assign O_100 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_100;
assign O_101 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_101;
assign O_102 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_102;
assign O_103 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_103;
assign O_104 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_104;
assign O_105 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_105;
assign O_106 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_106;
assign O_107 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_107;
assign O_108 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_108;
assign O_109 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_109;
assign O_11 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
assign O_110 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_110;
assign O_111 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_111;
assign O_112 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_112;
assign O_113 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_113;
assign O_114 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_114;
assign O_115 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_115;
assign O_116 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_116;
assign O_117 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_117;
assign O_118 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_118;
assign O_119 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_119;
assign O_12 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
assign O_120 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_120;
assign O_121 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_121;
assign O_122 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_122;
assign O_123 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_123;
assign O_124 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_124;
assign O_125 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_125;
assign O_126 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_126;
assign O_127 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_127;
assign O_128 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_128;
assign O_129 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_129;
assign O_13 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
assign O_130 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_130;
assign O_131 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_131;
assign O_132 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_132;
assign O_133 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_133;
assign O_134 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_134;
assign O_135 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_135;
assign O_136 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_136;
assign O_137 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_137;
assign O_138 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_138;
assign O_139 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_139;
assign O_14 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
assign O_140 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_140;
assign O_141 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_141;
assign O_142 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_142;
assign O_143 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_143;
assign O_144 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_144;
assign O_145 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_145;
assign O_146 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_146;
assign O_147 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_147;
assign O_148 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_148;
assign O_149 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_149;
assign O_15 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
assign O_150 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_150;
assign O_151 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_151;
assign O_152 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_152;
assign O_153 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_153;
assign O_154 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_154;
assign O_155 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_155;
assign O_156 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_156;
assign O_157 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_157;
assign O_158 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_158;
assign O_159 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_159;
assign O_16 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
assign O_160 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_160;
assign O_161 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_161;
assign O_162 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_162;
assign O_163 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_163;
assign O_164 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_164;
assign O_165 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_165;
assign O_166 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_166;
assign O_167 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_167;
assign O_168 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_168;
assign O_169 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_169;
assign O_17 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
assign O_170 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_170;
assign O_171 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_171;
assign O_172 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_172;
assign O_173 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_173;
assign O_174 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_174;
assign O_175 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_175;
assign O_176 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_176;
assign O_177 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_177;
assign O_178 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_178;
assign O_179 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_179;
assign O_18 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
assign O_180 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_180;
assign O_181 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_181;
assign O_182 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_182;
assign O_183 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_183;
assign O_184 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_184;
assign O_185 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_185;
assign O_186 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_186;
assign O_187 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_187;
assign O_188 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_188;
assign O_189 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_189;
assign O_19 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
assign O_190 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_190;
assign O_191 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_191;
assign O_192 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_192;
assign O_193 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_193;
assign O_194 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_194;
assign O_195 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_195;
assign O_196 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_196;
assign O_197 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_197;
assign O_198 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_198;
assign O_199 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_199;
assign O_2 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
assign O_20 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20;
assign O_21 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21;
assign O_22 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22;
assign O_23 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23;
assign O_24 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24;
assign O_25 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25;
assign O_26 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26;
assign O_27 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27;
assign O_28 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28;
assign O_29 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29;
assign O_3 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
assign O_30 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30;
assign O_31 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31;
assign O_32 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32;
assign O_33 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33;
assign O_34 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34;
assign O_35 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35;
assign O_36 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36;
assign O_37 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37;
assign O_38 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38;
assign O_39 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39;
assign O_4 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
assign O_40 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_40;
assign O_41 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_41;
assign O_42 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_42;
assign O_43 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_43;
assign O_44 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_44;
assign O_45 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_45;
assign O_46 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_46;
assign O_47 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_47;
assign O_48 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_48;
assign O_49 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_49;
assign O_5 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
assign O_50 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_50;
assign O_51 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_51;
assign O_52 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_52;
assign O_53 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_53;
assign O_54 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_54;
assign O_55 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_55;
assign O_56 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_56;
assign O_57 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_57;
assign O_58 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_58;
assign O_59 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_59;
assign O_6 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
assign O_60 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_60;
assign O_61 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_61;
assign O_62 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_62;
assign O_63 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_63;
assign O_64 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_64;
assign O_65 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_65;
assign O_66 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_66;
assign O_67 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_67;
assign O_68 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_68;
assign O_69 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_69;
assign O_7 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
assign O_70 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_70;
assign O_71 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_71;
assign O_72 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_72;
assign O_73 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_73;
assign O_74 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_74;
assign O_75 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_75;
assign O_76 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_76;
assign O_77 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_77;
assign O_78 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_78;
assign O_79 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_79;
assign O_8 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
assign O_80 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_80;
assign O_81 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_81;
assign O_82 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_82;
assign O_83 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_83;
assign O_84 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_84;
assign O_85 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_85;
assign O_86 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_86;
assign O_87 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_87;
assign O_88 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_88;
assign O_89 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_89;
assign O_9 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
assign O_90 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_90;
assign O_91 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_91;
assign O_92 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_92;
assign O_93 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_93;
assign O_94 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_94;
assign O_95 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_95;
assign O_96 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_96;
assign O_97 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_97;
assign O_98 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_98;
assign O_99 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_99;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Counter1CER (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/, input RESET/*verilator public*/);
wire [0:0] Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O;
wire [0:0] const_1_1_out;
wire [0:0] coreir_add1_inst0_out;
Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1 Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0(.CE(CE), .CLK(CLK), .I(coreir_add1_inst0_out), .O(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O), .RESET(RESET));
coreir_const #(.value(1'h1), .width(1)) const_1_1(.out(const_1_1_out));
coreir_add #(.width(1)) coreir_add1_inst0(.in0(Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O), .in1(const_1_1_out), .out(coreir_add1_inst0_out));
assign O = Register_has_ce_True_has_reset_True_has_async_reset_False_type_Bits_n_1_inst0_O;
endmodule

module Counter1_Mod2CE (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] Counter1CER_inst0_O;
wire LUT1_2_inst0_O;
wire and_inst0_out;
Counter1CER Counter1CER_inst0(.CE(CE), .CLK(CLK), .O(Counter1CER_inst0_O), .RESET(and_inst0_out));
LUT1_2 LUT1_2_inst0(.I0(Counter1CER_inst0_O[0]), .O(LUT1_2_inst0_O));
corebit_and and_inst0(.in0(LUT1_2_inst0_O), .in1(CE), .out(and_inst0_out));
assign O = Counter1CER_inst0_O;
endmodule

module InitialDelayCounter_1 (input CE/*verilator public*/, input CLK/*verilator public*/, output valid/*verilator public*/);
wire [0:0] Counter1_Mod2CE_inst0_O;
wire and_inst0_out;
wire [0:0] coreir_const11_inst0_out;
wire coreir_eq_1_inst0_out;
wire coreir_ult1_inst0_out;
Counter1_Mod2CE Counter1_Mod2CE_inst0(.CE(and_inst0_out), .CLK(CLK), .O(Counter1_Mod2CE_inst0_O));
corebit_and and_inst0(.in0(CE), .in1(coreir_ult1_inst0_out), .out(and_inst0_out));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
coreir_eq #(.width(1)) coreir_eq_1_inst0(.in0(Counter1_Mod2CE_inst0_O), .in1(coreir_const11_inst0_out), .out(coreir_eq_1_inst0_out));
coreir_ult #(.width(1)) coreir_ult1_inst0(.in0(Counter1_Mod2CE_inst0_O), .in1(coreir_const11_inst0_out), .out(coreir_ult1_inst0_out));
assign valid = coreir_eq_1_inst0_out;
endmodule

module Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire InitialDelayCounter_1_inst0_valid;
wire [7:0] LUT_Array_8_Bit_t_1n_inst0_data;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
InitialDelayCounter_1 InitialDelayCounter_1_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .valid(InitialDelayCounter_1_inst0_valid));
LUT_Array_8_Bit_t_1n LUT_Array_8_Bit_t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data(LUT_Array_8_Bit_t_1n_inst0_data));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(InitialDelayCounter_1_inst0_valid), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O = LUT_Array_8_Bit_t_1n_inst0_data;
assign valid_down = InitialDelayCounter_1_inst0_valid;
endmodule

module Add_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] coreir_add8_inst0_out;
coreir_add #(.width(8)) coreir_add8_inst0(.in0(I__0), .in1(I__1), .out(coreir_add8_inst0_out));
assign O = coreir_add8_inst0_out;
assign valid_down = valid_up;
endmodule

module Module_0 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Add_Atom_inst0_O;
wire Add_Atom_inst0_valid_down;
wire [7:0] Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O;
wire Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire and_inst0_out;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
Add_Atom Add_Atom_inst0(.I__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .I__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .O(Add_Atom_inst0_O), .valid_down(Add_Atom_inst0_valid_down), .valid_up(atomTupleCreator_t0Int_t1Int_inst0_valid_down));
Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .valid_down(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(valid_up), .in1(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I), .I1(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(and_inst0_out));
assign O = Add_Atom_inst0_O;
assign valid_down = Add_Atom_inst0_valid_down;
endmodule

module NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Module_0_inst0_O;
wire Module_0_inst0_valid_down;
wire [7:0] Module_0_inst1_O;
wire Module_0_inst1_valid_down;
wire [7:0] Module_0_inst10_O;
wire Module_0_inst10_valid_down;
wire [7:0] Module_0_inst100_O;
wire Module_0_inst100_valid_down;
wire [7:0] Module_0_inst101_O;
wire Module_0_inst101_valid_down;
wire [7:0] Module_0_inst102_O;
wire Module_0_inst102_valid_down;
wire [7:0] Module_0_inst103_O;
wire Module_0_inst103_valid_down;
wire [7:0] Module_0_inst104_O;
wire Module_0_inst104_valid_down;
wire [7:0] Module_0_inst105_O;
wire Module_0_inst105_valid_down;
wire [7:0] Module_0_inst106_O;
wire Module_0_inst106_valid_down;
wire [7:0] Module_0_inst107_O;
wire Module_0_inst107_valid_down;
wire [7:0] Module_0_inst108_O;
wire Module_0_inst108_valid_down;
wire [7:0] Module_0_inst109_O;
wire Module_0_inst109_valid_down;
wire [7:0] Module_0_inst11_O;
wire Module_0_inst11_valid_down;
wire [7:0] Module_0_inst110_O;
wire Module_0_inst110_valid_down;
wire [7:0] Module_0_inst111_O;
wire Module_0_inst111_valid_down;
wire [7:0] Module_0_inst112_O;
wire Module_0_inst112_valid_down;
wire [7:0] Module_0_inst113_O;
wire Module_0_inst113_valid_down;
wire [7:0] Module_0_inst114_O;
wire Module_0_inst114_valid_down;
wire [7:0] Module_0_inst115_O;
wire Module_0_inst115_valid_down;
wire [7:0] Module_0_inst116_O;
wire Module_0_inst116_valid_down;
wire [7:0] Module_0_inst117_O;
wire Module_0_inst117_valid_down;
wire [7:0] Module_0_inst118_O;
wire Module_0_inst118_valid_down;
wire [7:0] Module_0_inst119_O;
wire Module_0_inst119_valid_down;
wire [7:0] Module_0_inst12_O;
wire Module_0_inst12_valid_down;
wire [7:0] Module_0_inst120_O;
wire Module_0_inst120_valid_down;
wire [7:0] Module_0_inst121_O;
wire Module_0_inst121_valid_down;
wire [7:0] Module_0_inst122_O;
wire Module_0_inst122_valid_down;
wire [7:0] Module_0_inst123_O;
wire Module_0_inst123_valid_down;
wire [7:0] Module_0_inst124_O;
wire Module_0_inst124_valid_down;
wire [7:0] Module_0_inst125_O;
wire Module_0_inst125_valid_down;
wire [7:0] Module_0_inst126_O;
wire Module_0_inst126_valid_down;
wire [7:0] Module_0_inst127_O;
wire Module_0_inst127_valid_down;
wire [7:0] Module_0_inst128_O;
wire Module_0_inst128_valid_down;
wire [7:0] Module_0_inst129_O;
wire Module_0_inst129_valid_down;
wire [7:0] Module_0_inst13_O;
wire Module_0_inst13_valid_down;
wire [7:0] Module_0_inst130_O;
wire Module_0_inst130_valid_down;
wire [7:0] Module_0_inst131_O;
wire Module_0_inst131_valid_down;
wire [7:0] Module_0_inst132_O;
wire Module_0_inst132_valid_down;
wire [7:0] Module_0_inst133_O;
wire Module_0_inst133_valid_down;
wire [7:0] Module_0_inst134_O;
wire Module_0_inst134_valid_down;
wire [7:0] Module_0_inst135_O;
wire Module_0_inst135_valid_down;
wire [7:0] Module_0_inst136_O;
wire Module_0_inst136_valid_down;
wire [7:0] Module_0_inst137_O;
wire Module_0_inst137_valid_down;
wire [7:0] Module_0_inst138_O;
wire Module_0_inst138_valid_down;
wire [7:0] Module_0_inst139_O;
wire Module_0_inst139_valid_down;
wire [7:0] Module_0_inst14_O;
wire Module_0_inst14_valid_down;
wire [7:0] Module_0_inst140_O;
wire Module_0_inst140_valid_down;
wire [7:0] Module_0_inst141_O;
wire Module_0_inst141_valid_down;
wire [7:0] Module_0_inst142_O;
wire Module_0_inst142_valid_down;
wire [7:0] Module_0_inst143_O;
wire Module_0_inst143_valid_down;
wire [7:0] Module_0_inst144_O;
wire Module_0_inst144_valid_down;
wire [7:0] Module_0_inst145_O;
wire Module_0_inst145_valid_down;
wire [7:0] Module_0_inst146_O;
wire Module_0_inst146_valid_down;
wire [7:0] Module_0_inst147_O;
wire Module_0_inst147_valid_down;
wire [7:0] Module_0_inst148_O;
wire Module_0_inst148_valid_down;
wire [7:0] Module_0_inst149_O;
wire Module_0_inst149_valid_down;
wire [7:0] Module_0_inst15_O;
wire Module_0_inst15_valid_down;
wire [7:0] Module_0_inst150_O;
wire Module_0_inst150_valid_down;
wire [7:0] Module_0_inst151_O;
wire Module_0_inst151_valid_down;
wire [7:0] Module_0_inst152_O;
wire Module_0_inst152_valid_down;
wire [7:0] Module_0_inst153_O;
wire Module_0_inst153_valid_down;
wire [7:0] Module_0_inst154_O;
wire Module_0_inst154_valid_down;
wire [7:0] Module_0_inst155_O;
wire Module_0_inst155_valid_down;
wire [7:0] Module_0_inst156_O;
wire Module_0_inst156_valid_down;
wire [7:0] Module_0_inst157_O;
wire Module_0_inst157_valid_down;
wire [7:0] Module_0_inst158_O;
wire Module_0_inst158_valid_down;
wire [7:0] Module_0_inst159_O;
wire Module_0_inst159_valid_down;
wire [7:0] Module_0_inst16_O;
wire Module_0_inst16_valid_down;
wire [7:0] Module_0_inst160_O;
wire Module_0_inst160_valid_down;
wire [7:0] Module_0_inst161_O;
wire Module_0_inst161_valid_down;
wire [7:0] Module_0_inst162_O;
wire Module_0_inst162_valid_down;
wire [7:0] Module_0_inst163_O;
wire Module_0_inst163_valid_down;
wire [7:0] Module_0_inst164_O;
wire Module_0_inst164_valid_down;
wire [7:0] Module_0_inst165_O;
wire Module_0_inst165_valid_down;
wire [7:0] Module_0_inst166_O;
wire Module_0_inst166_valid_down;
wire [7:0] Module_0_inst167_O;
wire Module_0_inst167_valid_down;
wire [7:0] Module_0_inst168_O;
wire Module_0_inst168_valid_down;
wire [7:0] Module_0_inst169_O;
wire Module_0_inst169_valid_down;
wire [7:0] Module_0_inst17_O;
wire Module_0_inst17_valid_down;
wire [7:0] Module_0_inst170_O;
wire Module_0_inst170_valid_down;
wire [7:0] Module_0_inst171_O;
wire Module_0_inst171_valid_down;
wire [7:0] Module_0_inst172_O;
wire Module_0_inst172_valid_down;
wire [7:0] Module_0_inst173_O;
wire Module_0_inst173_valid_down;
wire [7:0] Module_0_inst174_O;
wire Module_0_inst174_valid_down;
wire [7:0] Module_0_inst175_O;
wire Module_0_inst175_valid_down;
wire [7:0] Module_0_inst176_O;
wire Module_0_inst176_valid_down;
wire [7:0] Module_0_inst177_O;
wire Module_0_inst177_valid_down;
wire [7:0] Module_0_inst178_O;
wire Module_0_inst178_valid_down;
wire [7:0] Module_0_inst179_O;
wire Module_0_inst179_valid_down;
wire [7:0] Module_0_inst18_O;
wire Module_0_inst18_valid_down;
wire [7:0] Module_0_inst180_O;
wire Module_0_inst180_valid_down;
wire [7:0] Module_0_inst181_O;
wire Module_0_inst181_valid_down;
wire [7:0] Module_0_inst182_O;
wire Module_0_inst182_valid_down;
wire [7:0] Module_0_inst183_O;
wire Module_0_inst183_valid_down;
wire [7:0] Module_0_inst184_O;
wire Module_0_inst184_valid_down;
wire [7:0] Module_0_inst185_O;
wire Module_0_inst185_valid_down;
wire [7:0] Module_0_inst186_O;
wire Module_0_inst186_valid_down;
wire [7:0] Module_0_inst187_O;
wire Module_0_inst187_valid_down;
wire [7:0] Module_0_inst188_O;
wire Module_0_inst188_valid_down;
wire [7:0] Module_0_inst189_O;
wire Module_0_inst189_valid_down;
wire [7:0] Module_0_inst19_O;
wire Module_0_inst19_valid_down;
wire [7:0] Module_0_inst190_O;
wire Module_0_inst190_valid_down;
wire [7:0] Module_0_inst191_O;
wire Module_0_inst191_valid_down;
wire [7:0] Module_0_inst192_O;
wire Module_0_inst192_valid_down;
wire [7:0] Module_0_inst193_O;
wire Module_0_inst193_valid_down;
wire [7:0] Module_0_inst194_O;
wire Module_0_inst194_valid_down;
wire [7:0] Module_0_inst195_O;
wire Module_0_inst195_valid_down;
wire [7:0] Module_0_inst196_O;
wire Module_0_inst196_valid_down;
wire [7:0] Module_0_inst197_O;
wire Module_0_inst197_valid_down;
wire [7:0] Module_0_inst198_O;
wire Module_0_inst198_valid_down;
wire [7:0] Module_0_inst199_O;
wire Module_0_inst199_valid_down;
wire [7:0] Module_0_inst2_O;
wire Module_0_inst2_valid_down;
wire [7:0] Module_0_inst20_O;
wire Module_0_inst20_valid_down;
wire [7:0] Module_0_inst21_O;
wire Module_0_inst21_valid_down;
wire [7:0] Module_0_inst22_O;
wire Module_0_inst22_valid_down;
wire [7:0] Module_0_inst23_O;
wire Module_0_inst23_valid_down;
wire [7:0] Module_0_inst24_O;
wire Module_0_inst24_valid_down;
wire [7:0] Module_0_inst25_O;
wire Module_0_inst25_valid_down;
wire [7:0] Module_0_inst26_O;
wire Module_0_inst26_valid_down;
wire [7:0] Module_0_inst27_O;
wire Module_0_inst27_valid_down;
wire [7:0] Module_0_inst28_O;
wire Module_0_inst28_valid_down;
wire [7:0] Module_0_inst29_O;
wire Module_0_inst29_valid_down;
wire [7:0] Module_0_inst3_O;
wire Module_0_inst3_valid_down;
wire [7:0] Module_0_inst30_O;
wire Module_0_inst30_valid_down;
wire [7:0] Module_0_inst31_O;
wire Module_0_inst31_valid_down;
wire [7:0] Module_0_inst32_O;
wire Module_0_inst32_valid_down;
wire [7:0] Module_0_inst33_O;
wire Module_0_inst33_valid_down;
wire [7:0] Module_0_inst34_O;
wire Module_0_inst34_valid_down;
wire [7:0] Module_0_inst35_O;
wire Module_0_inst35_valid_down;
wire [7:0] Module_0_inst36_O;
wire Module_0_inst36_valid_down;
wire [7:0] Module_0_inst37_O;
wire Module_0_inst37_valid_down;
wire [7:0] Module_0_inst38_O;
wire Module_0_inst38_valid_down;
wire [7:0] Module_0_inst39_O;
wire Module_0_inst39_valid_down;
wire [7:0] Module_0_inst4_O;
wire Module_0_inst4_valid_down;
wire [7:0] Module_0_inst40_O;
wire Module_0_inst40_valid_down;
wire [7:0] Module_0_inst41_O;
wire Module_0_inst41_valid_down;
wire [7:0] Module_0_inst42_O;
wire Module_0_inst42_valid_down;
wire [7:0] Module_0_inst43_O;
wire Module_0_inst43_valid_down;
wire [7:0] Module_0_inst44_O;
wire Module_0_inst44_valid_down;
wire [7:0] Module_0_inst45_O;
wire Module_0_inst45_valid_down;
wire [7:0] Module_0_inst46_O;
wire Module_0_inst46_valid_down;
wire [7:0] Module_0_inst47_O;
wire Module_0_inst47_valid_down;
wire [7:0] Module_0_inst48_O;
wire Module_0_inst48_valid_down;
wire [7:0] Module_0_inst49_O;
wire Module_0_inst49_valid_down;
wire [7:0] Module_0_inst5_O;
wire Module_0_inst5_valid_down;
wire [7:0] Module_0_inst50_O;
wire Module_0_inst50_valid_down;
wire [7:0] Module_0_inst51_O;
wire Module_0_inst51_valid_down;
wire [7:0] Module_0_inst52_O;
wire Module_0_inst52_valid_down;
wire [7:0] Module_0_inst53_O;
wire Module_0_inst53_valid_down;
wire [7:0] Module_0_inst54_O;
wire Module_0_inst54_valid_down;
wire [7:0] Module_0_inst55_O;
wire Module_0_inst55_valid_down;
wire [7:0] Module_0_inst56_O;
wire Module_0_inst56_valid_down;
wire [7:0] Module_0_inst57_O;
wire Module_0_inst57_valid_down;
wire [7:0] Module_0_inst58_O;
wire Module_0_inst58_valid_down;
wire [7:0] Module_0_inst59_O;
wire Module_0_inst59_valid_down;
wire [7:0] Module_0_inst6_O;
wire Module_0_inst6_valid_down;
wire [7:0] Module_0_inst60_O;
wire Module_0_inst60_valid_down;
wire [7:0] Module_0_inst61_O;
wire Module_0_inst61_valid_down;
wire [7:0] Module_0_inst62_O;
wire Module_0_inst62_valid_down;
wire [7:0] Module_0_inst63_O;
wire Module_0_inst63_valid_down;
wire [7:0] Module_0_inst64_O;
wire Module_0_inst64_valid_down;
wire [7:0] Module_0_inst65_O;
wire Module_0_inst65_valid_down;
wire [7:0] Module_0_inst66_O;
wire Module_0_inst66_valid_down;
wire [7:0] Module_0_inst67_O;
wire Module_0_inst67_valid_down;
wire [7:0] Module_0_inst68_O;
wire Module_0_inst68_valid_down;
wire [7:0] Module_0_inst69_O;
wire Module_0_inst69_valid_down;
wire [7:0] Module_0_inst7_O;
wire Module_0_inst7_valid_down;
wire [7:0] Module_0_inst70_O;
wire Module_0_inst70_valid_down;
wire [7:0] Module_0_inst71_O;
wire Module_0_inst71_valid_down;
wire [7:0] Module_0_inst72_O;
wire Module_0_inst72_valid_down;
wire [7:0] Module_0_inst73_O;
wire Module_0_inst73_valid_down;
wire [7:0] Module_0_inst74_O;
wire Module_0_inst74_valid_down;
wire [7:0] Module_0_inst75_O;
wire Module_0_inst75_valid_down;
wire [7:0] Module_0_inst76_O;
wire Module_0_inst76_valid_down;
wire [7:0] Module_0_inst77_O;
wire Module_0_inst77_valid_down;
wire [7:0] Module_0_inst78_O;
wire Module_0_inst78_valid_down;
wire [7:0] Module_0_inst79_O;
wire Module_0_inst79_valid_down;
wire [7:0] Module_0_inst8_O;
wire Module_0_inst8_valid_down;
wire [7:0] Module_0_inst80_O;
wire Module_0_inst80_valid_down;
wire [7:0] Module_0_inst81_O;
wire Module_0_inst81_valid_down;
wire [7:0] Module_0_inst82_O;
wire Module_0_inst82_valid_down;
wire [7:0] Module_0_inst83_O;
wire Module_0_inst83_valid_down;
wire [7:0] Module_0_inst84_O;
wire Module_0_inst84_valid_down;
wire [7:0] Module_0_inst85_O;
wire Module_0_inst85_valid_down;
wire [7:0] Module_0_inst86_O;
wire Module_0_inst86_valid_down;
wire [7:0] Module_0_inst87_O;
wire Module_0_inst87_valid_down;
wire [7:0] Module_0_inst88_O;
wire Module_0_inst88_valid_down;
wire [7:0] Module_0_inst89_O;
wire Module_0_inst89_valid_down;
wire [7:0] Module_0_inst9_O;
wire Module_0_inst9_valid_down;
wire [7:0] Module_0_inst90_O;
wire Module_0_inst90_valid_down;
wire [7:0] Module_0_inst91_O;
wire Module_0_inst91_valid_down;
wire [7:0] Module_0_inst92_O;
wire Module_0_inst92_valid_down;
wire [7:0] Module_0_inst93_O;
wire Module_0_inst93_valid_down;
wire [7:0] Module_0_inst94_O;
wire Module_0_inst94_valid_down;
wire [7:0] Module_0_inst95_O;
wire Module_0_inst95_valid_down;
wire [7:0] Module_0_inst96_O;
wire Module_0_inst96_valid_down;
wire [7:0] Module_0_inst97_O;
wire Module_0_inst97_valid_down;
wire [7:0] Module_0_inst98_O;
wire Module_0_inst98_valid_down;
wire [7:0] Module_0_inst99_O;
wire Module_0_inst99_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst100_out;
wire and_inst101_out;
wire and_inst102_out;
wire and_inst103_out;
wire and_inst104_out;
wire and_inst105_out;
wire and_inst106_out;
wire and_inst107_out;
wire and_inst108_out;
wire and_inst109_out;
wire and_inst11_out;
wire and_inst110_out;
wire and_inst111_out;
wire and_inst112_out;
wire and_inst113_out;
wire and_inst114_out;
wire and_inst115_out;
wire and_inst116_out;
wire and_inst117_out;
wire and_inst118_out;
wire and_inst119_out;
wire and_inst12_out;
wire and_inst120_out;
wire and_inst121_out;
wire and_inst122_out;
wire and_inst123_out;
wire and_inst124_out;
wire and_inst125_out;
wire and_inst126_out;
wire and_inst127_out;
wire and_inst128_out;
wire and_inst129_out;
wire and_inst13_out;
wire and_inst130_out;
wire and_inst131_out;
wire and_inst132_out;
wire and_inst133_out;
wire and_inst134_out;
wire and_inst135_out;
wire and_inst136_out;
wire and_inst137_out;
wire and_inst138_out;
wire and_inst139_out;
wire and_inst14_out;
wire and_inst140_out;
wire and_inst141_out;
wire and_inst142_out;
wire and_inst143_out;
wire and_inst144_out;
wire and_inst145_out;
wire and_inst146_out;
wire and_inst147_out;
wire and_inst148_out;
wire and_inst149_out;
wire and_inst15_out;
wire and_inst150_out;
wire and_inst151_out;
wire and_inst152_out;
wire and_inst153_out;
wire and_inst154_out;
wire and_inst155_out;
wire and_inst156_out;
wire and_inst157_out;
wire and_inst158_out;
wire and_inst159_out;
wire and_inst16_out;
wire and_inst160_out;
wire and_inst161_out;
wire and_inst162_out;
wire and_inst163_out;
wire and_inst164_out;
wire and_inst165_out;
wire and_inst166_out;
wire and_inst167_out;
wire and_inst168_out;
wire and_inst169_out;
wire and_inst17_out;
wire and_inst170_out;
wire and_inst171_out;
wire and_inst172_out;
wire and_inst173_out;
wire and_inst174_out;
wire and_inst175_out;
wire and_inst176_out;
wire and_inst177_out;
wire and_inst178_out;
wire and_inst179_out;
wire and_inst18_out;
wire and_inst180_out;
wire and_inst181_out;
wire and_inst182_out;
wire and_inst183_out;
wire and_inst184_out;
wire and_inst185_out;
wire and_inst186_out;
wire and_inst187_out;
wire and_inst188_out;
wire and_inst189_out;
wire and_inst19_out;
wire and_inst190_out;
wire and_inst191_out;
wire and_inst192_out;
wire and_inst193_out;
wire and_inst194_out;
wire and_inst195_out;
wire and_inst196_out;
wire and_inst197_out;
wire and_inst198_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst26_out;
wire and_inst27_out;
wire and_inst28_out;
wire and_inst29_out;
wire and_inst3_out;
wire and_inst30_out;
wire and_inst31_out;
wire and_inst32_out;
wire and_inst33_out;
wire and_inst34_out;
wire and_inst35_out;
wire and_inst36_out;
wire and_inst37_out;
wire and_inst38_out;
wire and_inst39_out;
wire and_inst4_out;
wire and_inst40_out;
wire and_inst41_out;
wire and_inst42_out;
wire and_inst43_out;
wire and_inst44_out;
wire and_inst45_out;
wire and_inst46_out;
wire and_inst47_out;
wire and_inst48_out;
wire and_inst49_out;
wire and_inst5_out;
wire and_inst50_out;
wire and_inst51_out;
wire and_inst52_out;
wire and_inst53_out;
wire and_inst54_out;
wire and_inst55_out;
wire and_inst56_out;
wire and_inst57_out;
wire and_inst58_out;
wire and_inst59_out;
wire and_inst6_out;
wire and_inst60_out;
wire and_inst61_out;
wire and_inst62_out;
wire and_inst63_out;
wire and_inst64_out;
wire and_inst65_out;
wire and_inst66_out;
wire and_inst67_out;
wire and_inst68_out;
wire and_inst69_out;
wire and_inst7_out;
wire and_inst70_out;
wire and_inst71_out;
wire and_inst72_out;
wire and_inst73_out;
wire and_inst74_out;
wire and_inst75_out;
wire and_inst76_out;
wire and_inst77_out;
wire and_inst78_out;
wire and_inst79_out;
wire and_inst8_out;
wire and_inst80_out;
wire and_inst81_out;
wire and_inst82_out;
wire and_inst83_out;
wire and_inst84_out;
wire and_inst85_out;
wire and_inst86_out;
wire and_inst87_out;
wire and_inst88_out;
wire and_inst89_out;
wire and_inst9_out;
wire and_inst90_out;
wire and_inst91_out;
wire and_inst92_out;
wire and_inst93_out;
wire and_inst94_out;
wire and_inst95_out;
wire and_inst96_out;
wire and_inst97_out;
wire and_inst98_out;
wire and_inst99_out;
Module_0 Module_0_inst0(.CLK(CLK), .I(I_0), .O(Module_0_inst0_O), .valid_down(Module_0_inst0_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst1(.CLK(CLK), .I(I_1), .O(Module_0_inst1_O), .valid_down(Module_0_inst1_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst10(.CLK(CLK), .I(I_10), .O(Module_0_inst10_O), .valid_down(Module_0_inst10_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst100(.CLK(CLK), .I(I_100), .O(Module_0_inst100_O), .valid_down(Module_0_inst100_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst101(.CLK(CLK), .I(I_101), .O(Module_0_inst101_O), .valid_down(Module_0_inst101_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst102(.CLK(CLK), .I(I_102), .O(Module_0_inst102_O), .valid_down(Module_0_inst102_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst103(.CLK(CLK), .I(I_103), .O(Module_0_inst103_O), .valid_down(Module_0_inst103_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst104(.CLK(CLK), .I(I_104), .O(Module_0_inst104_O), .valid_down(Module_0_inst104_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst105(.CLK(CLK), .I(I_105), .O(Module_0_inst105_O), .valid_down(Module_0_inst105_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst106(.CLK(CLK), .I(I_106), .O(Module_0_inst106_O), .valid_down(Module_0_inst106_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst107(.CLK(CLK), .I(I_107), .O(Module_0_inst107_O), .valid_down(Module_0_inst107_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst108(.CLK(CLK), .I(I_108), .O(Module_0_inst108_O), .valid_down(Module_0_inst108_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst109(.CLK(CLK), .I(I_109), .O(Module_0_inst109_O), .valid_down(Module_0_inst109_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst11(.CLK(CLK), .I(I_11), .O(Module_0_inst11_O), .valid_down(Module_0_inst11_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst110(.CLK(CLK), .I(I_110), .O(Module_0_inst110_O), .valid_down(Module_0_inst110_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst111(.CLK(CLK), .I(I_111), .O(Module_0_inst111_O), .valid_down(Module_0_inst111_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst112(.CLK(CLK), .I(I_112), .O(Module_0_inst112_O), .valid_down(Module_0_inst112_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst113(.CLK(CLK), .I(I_113), .O(Module_0_inst113_O), .valid_down(Module_0_inst113_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst114(.CLK(CLK), .I(I_114), .O(Module_0_inst114_O), .valid_down(Module_0_inst114_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst115(.CLK(CLK), .I(I_115), .O(Module_0_inst115_O), .valid_down(Module_0_inst115_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst116(.CLK(CLK), .I(I_116), .O(Module_0_inst116_O), .valid_down(Module_0_inst116_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst117(.CLK(CLK), .I(I_117), .O(Module_0_inst117_O), .valid_down(Module_0_inst117_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst118(.CLK(CLK), .I(I_118), .O(Module_0_inst118_O), .valid_down(Module_0_inst118_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst119(.CLK(CLK), .I(I_119), .O(Module_0_inst119_O), .valid_down(Module_0_inst119_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst12(.CLK(CLK), .I(I_12), .O(Module_0_inst12_O), .valid_down(Module_0_inst12_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst120(.CLK(CLK), .I(I_120), .O(Module_0_inst120_O), .valid_down(Module_0_inst120_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst121(.CLK(CLK), .I(I_121), .O(Module_0_inst121_O), .valid_down(Module_0_inst121_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst122(.CLK(CLK), .I(I_122), .O(Module_0_inst122_O), .valid_down(Module_0_inst122_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst123(.CLK(CLK), .I(I_123), .O(Module_0_inst123_O), .valid_down(Module_0_inst123_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst124(.CLK(CLK), .I(I_124), .O(Module_0_inst124_O), .valid_down(Module_0_inst124_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst125(.CLK(CLK), .I(I_125), .O(Module_0_inst125_O), .valid_down(Module_0_inst125_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst126(.CLK(CLK), .I(I_126), .O(Module_0_inst126_O), .valid_down(Module_0_inst126_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst127(.CLK(CLK), .I(I_127), .O(Module_0_inst127_O), .valid_down(Module_0_inst127_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst128(.CLK(CLK), .I(I_128), .O(Module_0_inst128_O), .valid_down(Module_0_inst128_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst129(.CLK(CLK), .I(I_129), .O(Module_0_inst129_O), .valid_down(Module_0_inst129_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst13(.CLK(CLK), .I(I_13), .O(Module_0_inst13_O), .valid_down(Module_0_inst13_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst130(.CLK(CLK), .I(I_130), .O(Module_0_inst130_O), .valid_down(Module_0_inst130_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst131(.CLK(CLK), .I(I_131), .O(Module_0_inst131_O), .valid_down(Module_0_inst131_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst132(.CLK(CLK), .I(I_132), .O(Module_0_inst132_O), .valid_down(Module_0_inst132_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst133(.CLK(CLK), .I(I_133), .O(Module_0_inst133_O), .valid_down(Module_0_inst133_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst134(.CLK(CLK), .I(I_134), .O(Module_0_inst134_O), .valid_down(Module_0_inst134_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst135(.CLK(CLK), .I(I_135), .O(Module_0_inst135_O), .valid_down(Module_0_inst135_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst136(.CLK(CLK), .I(I_136), .O(Module_0_inst136_O), .valid_down(Module_0_inst136_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst137(.CLK(CLK), .I(I_137), .O(Module_0_inst137_O), .valid_down(Module_0_inst137_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst138(.CLK(CLK), .I(I_138), .O(Module_0_inst138_O), .valid_down(Module_0_inst138_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst139(.CLK(CLK), .I(I_139), .O(Module_0_inst139_O), .valid_down(Module_0_inst139_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst14(.CLK(CLK), .I(I_14), .O(Module_0_inst14_O), .valid_down(Module_0_inst14_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst140(.CLK(CLK), .I(I_140), .O(Module_0_inst140_O), .valid_down(Module_0_inst140_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst141(.CLK(CLK), .I(I_141), .O(Module_0_inst141_O), .valid_down(Module_0_inst141_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst142(.CLK(CLK), .I(I_142), .O(Module_0_inst142_O), .valid_down(Module_0_inst142_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst143(.CLK(CLK), .I(I_143), .O(Module_0_inst143_O), .valid_down(Module_0_inst143_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst144(.CLK(CLK), .I(I_144), .O(Module_0_inst144_O), .valid_down(Module_0_inst144_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst145(.CLK(CLK), .I(I_145), .O(Module_0_inst145_O), .valid_down(Module_0_inst145_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst146(.CLK(CLK), .I(I_146), .O(Module_0_inst146_O), .valid_down(Module_0_inst146_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst147(.CLK(CLK), .I(I_147), .O(Module_0_inst147_O), .valid_down(Module_0_inst147_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst148(.CLK(CLK), .I(I_148), .O(Module_0_inst148_O), .valid_down(Module_0_inst148_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst149(.CLK(CLK), .I(I_149), .O(Module_0_inst149_O), .valid_down(Module_0_inst149_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst15(.CLK(CLK), .I(I_15), .O(Module_0_inst15_O), .valid_down(Module_0_inst15_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst150(.CLK(CLK), .I(I_150), .O(Module_0_inst150_O), .valid_down(Module_0_inst150_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst151(.CLK(CLK), .I(I_151), .O(Module_0_inst151_O), .valid_down(Module_0_inst151_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst152(.CLK(CLK), .I(I_152), .O(Module_0_inst152_O), .valid_down(Module_0_inst152_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst153(.CLK(CLK), .I(I_153), .O(Module_0_inst153_O), .valid_down(Module_0_inst153_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst154(.CLK(CLK), .I(I_154), .O(Module_0_inst154_O), .valid_down(Module_0_inst154_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst155(.CLK(CLK), .I(I_155), .O(Module_0_inst155_O), .valid_down(Module_0_inst155_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst156(.CLK(CLK), .I(I_156), .O(Module_0_inst156_O), .valid_down(Module_0_inst156_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst157(.CLK(CLK), .I(I_157), .O(Module_0_inst157_O), .valid_down(Module_0_inst157_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst158(.CLK(CLK), .I(I_158), .O(Module_0_inst158_O), .valid_down(Module_0_inst158_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst159(.CLK(CLK), .I(I_159), .O(Module_0_inst159_O), .valid_down(Module_0_inst159_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst16(.CLK(CLK), .I(I_16), .O(Module_0_inst16_O), .valid_down(Module_0_inst16_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst160(.CLK(CLK), .I(I_160), .O(Module_0_inst160_O), .valid_down(Module_0_inst160_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst161(.CLK(CLK), .I(I_161), .O(Module_0_inst161_O), .valid_down(Module_0_inst161_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst162(.CLK(CLK), .I(I_162), .O(Module_0_inst162_O), .valid_down(Module_0_inst162_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst163(.CLK(CLK), .I(I_163), .O(Module_0_inst163_O), .valid_down(Module_0_inst163_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst164(.CLK(CLK), .I(I_164), .O(Module_0_inst164_O), .valid_down(Module_0_inst164_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst165(.CLK(CLK), .I(I_165), .O(Module_0_inst165_O), .valid_down(Module_0_inst165_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst166(.CLK(CLK), .I(I_166), .O(Module_0_inst166_O), .valid_down(Module_0_inst166_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst167(.CLK(CLK), .I(I_167), .O(Module_0_inst167_O), .valid_down(Module_0_inst167_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst168(.CLK(CLK), .I(I_168), .O(Module_0_inst168_O), .valid_down(Module_0_inst168_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst169(.CLK(CLK), .I(I_169), .O(Module_0_inst169_O), .valid_down(Module_0_inst169_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst17(.CLK(CLK), .I(I_17), .O(Module_0_inst17_O), .valid_down(Module_0_inst17_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst170(.CLK(CLK), .I(I_170), .O(Module_0_inst170_O), .valid_down(Module_0_inst170_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst171(.CLK(CLK), .I(I_171), .O(Module_0_inst171_O), .valid_down(Module_0_inst171_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst172(.CLK(CLK), .I(I_172), .O(Module_0_inst172_O), .valid_down(Module_0_inst172_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst173(.CLK(CLK), .I(I_173), .O(Module_0_inst173_O), .valid_down(Module_0_inst173_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst174(.CLK(CLK), .I(I_174), .O(Module_0_inst174_O), .valid_down(Module_0_inst174_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst175(.CLK(CLK), .I(I_175), .O(Module_0_inst175_O), .valid_down(Module_0_inst175_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst176(.CLK(CLK), .I(I_176), .O(Module_0_inst176_O), .valid_down(Module_0_inst176_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst177(.CLK(CLK), .I(I_177), .O(Module_0_inst177_O), .valid_down(Module_0_inst177_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst178(.CLK(CLK), .I(I_178), .O(Module_0_inst178_O), .valid_down(Module_0_inst178_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst179(.CLK(CLK), .I(I_179), .O(Module_0_inst179_O), .valid_down(Module_0_inst179_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst18(.CLK(CLK), .I(I_18), .O(Module_0_inst18_O), .valid_down(Module_0_inst18_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst180(.CLK(CLK), .I(I_180), .O(Module_0_inst180_O), .valid_down(Module_0_inst180_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst181(.CLK(CLK), .I(I_181), .O(Module_0_inst181_O), .valid_down(Module_0_inst181_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst182(.CLK(CLK), .I(I_182), .O(Module_0_inst182_O), .valid_down(Module_0_inst182_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst183(.CLK(CLK), .I(I_183), .O(Module_0_inst183_O), .valid_down(Module_0_inst183_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst184(.CLK(CLK), .I(I_184), .O(Module_0_inst184_O), .valid_down(Module_0_inst184_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst185(.CLK(CLK), .I(I_185), .O(Module_0_inst185_O), .valid_down(Module_0_inst185_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst186(.CLK(CLK), .I(I_186), .O(Module_0_inst186_O), .valid_down(Module_0_inst186_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst187(.CLK(CLK), .I(I_187), .O(Module_0_inst187_O), .valid_down(Module_0_inst187_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst188(.CLK(CLK), .I(I_188), .O(Module_0_inst188_O), .valid_down(Module_0_inst188_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst189(.CLK(CLK), .I(I_189), .O(Module_0_inst189_O), .valid_down(Module_0_inst189_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst19(.CLK(CLK), .I(I_19), .O(Module_0_inst19_O), .valid_down(Module_0_inst19_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst190(.CLK(CLK), .I(I_190), .O(Module_0_inst190_O), .valid_down(Module_0_inst190_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst191(.CLK(CLK), .I(I_191), .O(Module_0_inst191_O), .valid_down(Module_0_inst191_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst192(.CLK(CLK), .I(I_192), .O(Module_0_inst192_O), .valid_down(Module_0_inst192_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst193(.CLK(CLK), .I(I_193), .O(Module_0_inst193_O), .valid_down(Module_0_inst193_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst194(.CLK(CLK), .I(I_194), .O(Module_0_inst194_O), .valid_down(Module_0_inst194_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst195(.CLK(CLK), .I(I_195), .O(Module_0_inst195_O), .valid_down(Module_0_inst195_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst196(.CLK(CLK), .I(I_196), .O(Module_0_inst196_O), .valid_down(Module_0_inst196_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst197(.CLK(CLK), .I(I_197), .O(Module_0_inst197_O), .valid_down(Module_0_inst197_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst198(.CLK(CLK), .I(I_198), .O(Module_0_inst198_O), .valid_down(Module_0_inst198_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst199(.CLK(CLK), .I(I_199), .O(Module_0_inst199_O), .valid_down(Module_0_inst199_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst2(.CLK(CLK), .I(I_2), .O(Module_0_inst2_O), .valid_down(Module_0_inst2_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst20(.CLK(CLK), .I(I_20), .O(Module_0_inst20_O), .valid_down(Module_0_inst20_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst21(.CLK(CLK), .I(I_21), .O(Module_0_inst21_O), .valid_down(Module_0_inst21_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst22(.CLK(CLK), .I(I_22), .O(Module_0_inst22_O), .valid_down(Module_0_inst22_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst23(.CLK(CLK), .I(I_23), .O(Module_0_inst23_O), .valid_down(Module_0_inst23_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst24(.CLK(CLK), .I(I_24), .O(Module_0_inst24_O), .valid_down(Module_0_inst24_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst25(.CLK(CLK), .I(I_25), .O(Module_0_inst25_O), .valid_down(Module_0_inst25_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst26(.CLK(CLK), .I(I_26), .O(Module_0_inst26_O), .valid_down(Module_0_inst26_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst27(.CLK(CLK), .I(I_27), .O(Module_0_inst27_O), .valid_down(Module_0_inst27_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst28(.CLK(CLK), .I(I_28), .O(Module_0_inst28_O), .valid_down(Module_0_inst28_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst29(.CLK(CLK), .I(I_29), .O(Module_0_inst29_O), .valid_down(Module_0_inst29_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst3(.CLK(CLK), .I(I_3), .O(Module_0_inst3_O), .valid_down(Module_0_inst3_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst30(.CLK(CLK), .I(I_30), .O(Module_0_inst30_O), .valid_down(Module_0_inst30_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst31(.CLK(CLK), .I(I_31), .O(Module_0_inst31_O), .valid_down(Module_0_inst31_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst32(.CLK(CLK), .I(I_32), .O(Module_0_inst32_O), .valid_down(Module_0_inst32_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst33(.CLK(CLK), .I(I_33), .O(Module_0_inst33_O), .valid_down(Module_0_inst33_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst34(.CLK(CLK), .I(I_34), .O(Module_0_inst34_O), .valid_down(Module_0_inst34_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst35(.CLK(CLK), .I(I_35), .O(Module_0_inst35_O), .valid_down(Module_0_inst35_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst36(.CLK(CLK), .I(I_36), .O(Module_0_inst36_O), .valid_down(Module_0_inst36_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst37(.CLK(CLK), .I(I_37), .O(Module_0_inst37_O), .valid_down(Module_0_inst37_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst38(.CLK(CLK), .I(I_38), .O(Module_0_inst38_O), .valid_down(Module_0_inst38_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst39(.CLK(CLK), .I(I_39), .O(Module_0_inst39_O), .valid_down(Module_0_inst39_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst4(.CLK(CLK), .I(I_4), .O(Module_0_inst4_O), .valid_down(Module_0_inst4_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst40(.CLK(CLK), .I(I_40), .O(Module_0_inst40_O), .valid_down(Module_0_inst40_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst41(.CLK(CLK), .I(I_41), .O(Module_0_inst41_O), .valid_down(Module_0_inst41_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst42(.CLK(CLK), .I(I_42), .O(Module_0_inst42_O), .valid_down(Module_0_inst42_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst43(.CLK(CLK), .I(I_43), .O(Module_0_inst43_O), .valid_down(Module_0_inst43_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst44(.CLK(CLK), .I(I_44), .O(Module_0_inst44_O), .valid_down(Module_0_inst44_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst45(.CLK(CLK), .I(I_45), .O(Module_0_inst45_O), .valid_down(Module_0_inst45_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst46(.CLK(CLK), .I(I_46), .O(Module_0_inst46_O), .valid_down(Module_0_inst46_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst47(.CLK(CLK), .I(I_47), .O(Module_0_inst47_O), .valid_down(Module_0_inst47_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst48(.CLK(CLK), .I(I_48), .O(Module_0_inst48_O), .valid_down(Module_0_inst48_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst49(.CLK(CLK), .I(I_49), .O(Module_0_inst49_O), .valid_down(Module_0_inst49_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst5(.CLK(CLK), .I(I_5), .O(Module_0_inst5_O), .valid_down(Module_0_inst5_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst50(.CLK(CLK), .I(I_50), .O(Module_0_inst50_O), .valid_down(Module_0_inst50_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst51(.CLK(CLK), .I(I_51), .O(Module_0_inst51_O), .valid_down(Module_0_inst51_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst52(.CLK(CLK), .I(I_52), .O(Module_0_inst52_O), .valid_down(Module_0_inst52_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst53(.CLK(CLK), .I(I_53), .O(Module_0_inst53_O), .valid_down(Module_0_inst53_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst54(.CLK(CLK), .I(I_54), .O(Module_0_inst54_O), .valid_down(Module_0_inst54_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst55(.CLK(CLK), .I(I_55), .O(Module_0_inst55_O), .valid_down(Module_0_inst55_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst56(.CLK(CLK), .I(I_56), .O(Module_0_inst56_O), .valid_down(Module_0_inst56_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst57(.CLK(CLK), .I(I_57), .O(Module_0_inst57_O), .valid_down(Module_0_inst57_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst58(.CLK(CLK), .I(I_58), .O(Module_0_inst58_O), .valid_down(Module_0_inst58_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst59(.CLK(CLK), .I(I_59), .O(Module_0_inst59_O), .valid_down(Module_0_inst59_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst6(.CLK(CLK), .I(I_6), .O(Module_0_inst6_O), .valid_down(Module_0_inst6_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst60(.CLK(CLK), .I(I_60), .O(Module_0_inst60_O), .valid_down(Module_0_inst60_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst61(.CLK(CLK), .I(I_61), .O(Module_0_inst61_O), .valid_down(Module_0_inst61_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst62(.CLK(CLK), .I(I_62), .O(Module_0_inst62_O), .valid_down(Module_0_inst62_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst63(.CLK(CLK), .I(I_63), .O(Module_0_inst63_O), .valid_down(Module_0_inst63_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst64(.CLK(CLK), .I(I_64), .O(Module_0_inst64_O), .valid_down(Module_0_inst64_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst65(.CLK(CLK), .I(I_65), .O(Module_0_inst65_O), .valid_down(Module_0_inst65_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst66(.CLK(CLK), .I(I_66), .O(Module_0_inst66_O), .valid_down(Module_0_inst66_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst67(.CLK(CLK), .I(I_67), .O(Module_0_inst67_O), .valid_down(Module_0_inst67_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst68(.CLK(CLK), .I(I_68), .O(Module_0_inst68_O), .valid_down(Module_0_inst68_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst69(.CLK(CLK), .I(I_69), .O(Module_0_inst69_O), .valid_down(Module_0_inst69_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst7(.CLK(CLK), .I(I_7), .O(Module_0_inst7_O), .valid_down(Module_0_inst7_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst70(.CLK(CLK), .I(I_70), .O(Module_0_inst70_O), .valid_down(Module_0_inst70_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst71(.CLK(CLK), .I(I_71), .O(Module_0_inst71_O), .valid_down(Module_0_inst71_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst72(.CLK(CLK), .I(I_72), .O(Module_0_inst72_O), .valid_down(Module_0_inst72_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst73(.CLK(CLK), .I(I_73), .O(Module_0_inst73_O), .valid_down(Module_0_inst73_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst74(.CLK(CLK), .I(I_74), .O(Module_0_inst74_O), .valid_down(Module_0_inst74_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst75(.CLK(CLK), .I(I_75), .O(Module_0_inst75_O), .valid_down(Module_0_inst75_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst76(.CLK(CLK), .I(I_76), .O(Module_0_inst76_O), .valid_down(Module_0_inst76_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst77(.CLK(CLK), .I(I_77), .O(Module_0_inst77_O), .valid_down(Module_0_inst77_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst78(.CLK(CLK), .I(I_78), .O(Module_0_inst78_O), .valid_down(Module_0_inst78_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst79(.CLK(CLK), .I(I_79), .O(Module_0_inst79_O), .valid_down(Module_0_inst79_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst8(.CLK(CLK), .I(I_8), .O(Module_0_inst8_O), .valid_down(Module_0_inst8_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst80(.CLK(CLK), .I(I_80), .O(Module_0_inst80_O), .valid_down(Module_0_inst80_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst81(.CLK(CLK), .I(I_81), .O(Module_0_inst81_O), .valid_down(Module_0_inst81_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst82(.CLK(CLK), .I(I_82), .O(Module_0_inst82_O), .valid_down(Module_0_inst82_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst83(.CLK(CLK), .I(I_83), .O(Module_0_inst83_O), .valid_down(Module_0_inst83_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst84(.CLK(CLK), .I(I_84), .O(Module_0_inst84_O), .valid_down(Module_0_inst84_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst85(.CLK(CLK), .I(I_85), .O(Module_0_inst85_O), .valid_down(Module_0_inst85_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst86(.CLK(CLK), .I(I_86), .O(Module_0_inst86_O), .valid_down(Module_0_inst86_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst87(.CLK(CLK), .I(I_87), .O(Module_0_inst87_O), .valid_down(Module_0_inst87_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst88(.CLK(CLK), .I(I_88), .O(Module_0_inst88_O), .valid_down(Module_0_inst88_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst89(.CLK(CLK), .I(I_89), .O(Module_0_inst89_O), .valid_down(Module_0_inst89_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst9(.CLK(CLK), .I(I_9), .O(Module_0_inst9_O), .valid_down(Module_0_inst9_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst90(.CLK(CLK), .I(I_90), .O(Module_0_inst90_O), .valid_down(Module_0_inst90_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst91(.CLK(CLK), .I(I_91), .O(Module_0_inst91_O), .valid_down(Module_0_inst91_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst92(.CLK(CLK), .I(I_92), .O(Module_0_inst92_O), .valid_down(Module_0_inst92_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst93(.CLK(CLK), .I(I_93), .O(Module_0_inst93_O), .valid_down(Module_0_inst93_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst94(.CLK(CLK), .I(I_94), .O(Module_0_inst94_O), .valid_down(Module_0_inst94_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst95(.CLK(CLK), .I(I_95), .O(Module_0_inst95_O), .valid_down(Module_0_inst95_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst96(.CLK(CLK), .I(I_96), .O(Module_0_inst96_O), .valid_down(Module_0_inst96_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst97(.CLK(CLK), .I(I_97), .O(Module_0_inst97_O), .valid_down(Module_0_inst97_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst98(.CLK(CLK), .I(I_98), .O(Module_0_inst98_O), .valid_down(Module_0_inst98_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst99(.CLK(CLK), .I(I_99), .O(Module_0_inst99_O), .valid_down(Module_0_inst99_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Module_0_inst0_valid_down), .in1(Module_0_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Module_0_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(Module_0_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst100(.in0(and_inst99_out), .in1(Module_0_inst101_valid_down), .out(and_inst100_out));
corebit_and and_inst101(.in0(and_inst100_out), .in1(Module_0_inst102_valid_down), .out(and_inst101_out));
corebit_and and_inst102(.in0(and_inst101_out), .in1(Module_0_inst103_valid_down), .out(and_inst102_out));
corebit_and and_inst103(.in0(and_inst102_out), .in1(Module_0_inst104_valid_down), .out(and_inst103_out));
corebit_and and_inst104(.in0(and_inst103_out), .in1(Module_0_inst105_valid_down), .out(and_inst104_out));
corebit_and and_inst105(.in0(and_inst104_out), .in1(Module_0_inst106_valid_down), .out(and_inst105_out));
corebit_and and_inst106(.in0(and_inst105_out), .in1(Module_0_inst107_valid_down), .out(and_inst106_out));
corebit_and and_inst107(.in0(and_inst106_out), .in1(Module_0_inst108_valid_down), .out(and_inst107_out));
corebit_and and_inst108(.in0(and_inst107_out), .in1(Module_0_inst109_valid_down), .out(and_inst108_out));
corebit_and and_inst109(.in0(and_inst108_out), .in1(Module_0_inst110_valid_down), .out(and_inst109_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(Module_0_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst110(.in0(and_inst109_out), .in1(Module_0_inst111_valid_down), .out(and_inst110_out));
corebit_and and_inst111(.in0(and_inst110_out), .in1(Module_0_inst112_valid_down), .out(and_inst111_out));
corebit_and and_inst112(.in0(and_inst111_out), .in1(Module_0_inst113_valid_down), .out(and_inst112_out));
corebit_and and_inst113(.in0(and_inst112_out), .in1(Module_0_inst114_valid_down), .out(and_inst113_out));
corebit_and and_inst114(.in0(and_inst113_out), .in1(Module_0_inst115_valid_down), .out(and_inst114_out));
corebit_and and_inst115(.in0(and_inst114_out), .in1(Module_0_inst116_valid_down), .out(and_inst115_out));
corebit_and and_inst116(.in0(and_inst115_out), .in1(Module_0_inst117_valid_down), .out(and_inst116_out));
corebit_and and_inst117(.in0(and_inst116_out), .in1(Module_0_inst118_valid_down), .out(and_inst117_out));
corebit_and and_inst118(.in0(and_inst117_out), .in1(Module_0_inst119_valid_down), .out(and_inst118_out));
corebit_and and_inst119(.in0(and_inst118_out), .in1(Module_0_inst120_valid_down), .out(and_inst119_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(Module_0_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst120(.in0(and_inst119_out), .in1(Module_0_inst121_valid_down), .out(and_inst120_out));
corebit_and and_inst121(.in0(and_inst120_out), .in1(Module_0_inst122_valid_down), .out(and_inst121_out));
corebit_and and_inst122(.in0(and_inst121_out), .in1(Module_0_inst123_valid_down), .out(and_inst122_out));
corebit_and and_inst123(.in0(and_inst122_out), .in1(Module_0_inst124_valid_down), .out(and_inst123_out));
corebit_and and_inst124(.in0(and_inst123_out), .in1(Module_0_inst125_valid_down), .out(and_inst124_out));
corebit_and and_inst125(.in0(and_inst124_out), .in1(Module_0_inst126_valid_down), .out(and_inst125_out));
corebit_and and_inst126(.in0(and_inst125_out), .in1(Module_0_inst127_valid_down), .out(and_inst126_out));
corebit_and and_inst127(.in0(and_inst126_out), .in1(Module_0_inst128_valid_down), .out(and_inst127_out));
corebit_and and_inst128(.in0(and_inst127_out), .in1(Module_0_inst129_valid_down), .out(and_inst128_out));
corebit_and and_inst129(.in0(and_inst128_out), .in1(Module_0_inst130_valid_down), .out(and_inst129_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(Module_0_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst130(.in0(and_inst129_out), .in1(Module_0_inst131_valid_down), .out(and_inst130_out));
corebit_and and_inst131(.in0(and_inst130_out), .in1(Module_0_inst132_valid_down), .out(and_inst131_out));
corebit_and and_inst132(.in0(and_inst131_out), .in1(Module_0_inst133_valid_down), .out(and_inst132_out));
corebit_and and_inst133(.in0(and_inst132_out), .in1(Module_0_inst134_valid_down), .out(and_inst133_out));
corebit_and and_inst134(.in0(and_inst133_out), .in1(Module_0_inst135_valid_down), .out(and_inst134_out));
corebit_and and_inst135(.in0(and_inst134_out), .in1(Module_0_inst136_valid_down), .out(and_inst135_out));
corebit_and and_inst136(.in0(and_inst135_out), .in1(Module_0_inst137_valid_down), .out(and_inst136_out));
corebit_and and_inst137(.in0(and_inst136_out), .in1(Module_0_inst138_valid_down), .out(and_inst137_out));
corebit_and and_inst138(.in0(and_inst137_out), .in1(Module_0_inst139_valid_down), .out(and_inst138_out));
corebit_and and_inst139(.in0(and_inst138_out), .in1(Module_0_inst140_valid_down), .out(and_inst139_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(Module_0_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst140(.in0(and_inst139_out), .in1(Module_0_inst141_valid_down), .out(and_inst140_out));
corebit_and and_inst141(.in0(and_inst140_out), .in1(Module_0_inst142_valid_down), .out(and_inst141_out));
corebit_and and_inst142(.in0(and_inst141_out), .in1(Module_0_inst143_valid_down), .out(and_inst142_out));
corebit_and and_inst143(.in0(and_inst142_out), .in1(Module_0_inst144_valid_down), .out(and_inst143_out));
corebit_and and_inst144(.in0(and_inst143_out), .in1(Module_0_inst145_valid_down), .out(and_inst144_out));
corebit_and and_inst145(.in0(and_inst144_out), .in1(Module_0_inst146_valid_down), .out(and_inst145_out));
corebit_and and_inst146(.in0(and_inst145_out), .in1(Module_0_inst147_valid_down), .out(and_inst146_out));
corebit_and and_inst147(.in0(and_inst146_out), .in1(Module_0_inst148_valid_down), .out(and_inst147_out));
corebit_and and_inst148(.in0(and_inst147_out), .in1(Module_0_inst149_valid_down), .out(and_inst148_out));
corebit_and and_inst149(.in0(and_inst148_out), .in1(Module_0_inst150_valid_down), .out(and_inst149_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(Module_0_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst150(.in0(and_inst149_out), .in1(Module_0_inst151_valid_down), .out(and_inst150_out));
corebit_and and_inst151(.in0(and_inst150_out), .in1(Module_0_inst152_valid_down), .out(and_inst151_out));
corebit_and and_inst152(.in0(and_inst151_out), .in1(Module_0_inst153_valid_down), .out(and_inst152_out));
corebit_and and_inst153(.in0(and_inst152_out), .in1(Module_0_inst154_valid_down), .out(and_inst153_out));
corebit_and and_inst154(.in0(and_inst153_out), .in1(Module_0_inst155_valid_down), .out(and_inst154_out));
corebit_and and_inst155(.in0(and_inst154_out), .in1(Module_0_inst156_valid_down), .out(and_inst155_out));
corebit_and and_inst156(.in0(and_inst155_out), .in1(Module_0_inst157_valid_down), .out(and_inst156_out));
corebit_and and_inst157(.in0(and_inst156_out), .in1(Module_0_inst158_valid_down), .out(and_inst157_out));
corebit_and and_inst158(.in0(and_inst157_out), .in1(Module_0_inst159_valid_down), .out(and_inst158_out));
corebit_and and_inst159(.in0(and_inst158_out), .in1(Module_0_inst160_valid_down), .out(and_inst159_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(Module_0_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst160(.in0(and_inst159_out), .in1(Module_0_inst161_valid_down), .out(and_inst160_out));
corebit_and and_inst161(.in0(and_inst160_out), .in1(Module_0_inst162_valid_down), .out(and_inst161_out));
corebit_and and_inst162(.in0(and_inst161_out), .in1(Module_0_inst163_valid_down), .out(and_inst162_out));
corebit_and and_inst163(.in0(and_inst162_out), .in1(Module_0_inst164_valid_down), .out(and_inst163_out));
corebit_and and_inst164(.in0(and_inst163_out), .in1(Module_0_inst165_valid_down), .out(and_inst164_out));
corebit_and and_inst165(.in0(and_inst164_out), .in1(Module_0_inst166_valid_down), .out(and_inst165_out));
corebit_and and_inst166(.in0(and_inst165_out), .in1(Module_0_inst167_valid_down), .out(and_inst166_out));
corebit_and and_inst167(.in0(and_inst166_out), .in1(Module_0_inst168_valid_down), .out(and_inst167_out));
corebit_and and_inst168(.in0(and_inst167_out), .in1(Module_0_inst169_valid_down), .out(and_inst168_out));
corebit_and and_inst169(.in0(and_inst168_out), .in1(Module_0_inst170_valid_down), .out(and_inst169_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(Module_0_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst170(.in0(and_inst169_out), .in1(Module_0_inst171_valid_down), .out(and_inst170_out));
corebit_and and_inst171(.in0(and_inst170_out), .in1(Module_0_inst172_valid_down), .out(and_inst171_out));
corebit_and and_inst172(.in0(and_inst171_out), .in1(Module_0_inst173_valid_down), .out(and_inst172_out));
corebit_and and_inst173(.in0(and_inst172_out), .in1(Module_0_inst174_valid_down), .out(and_inst173_out));
corebit_and and_inst174(.in0(and_inst173_out), .in1(Module_0_inst175_valid_down), .out(and_inst174_out));
corebit_and and_inst175(.in0(and_inst174_out), .in1(Module_0_inst176_valid_down), .out(and_inst175_out));
corebit_and and_inst176(.in0(and_inst175_out), .in1(Module_0_inst177_valid_down), .out(and_inst176_out));
corebit_and and_inst177(.in0(and_inst176_out), .in1(Module_0_inst178_valid_down), .out(and_inst177_out));
corebit_and and_inst178(.in0(and_inst177_out), .in1(Module_0_inst179_valid_down), .out(and_inst178_out));
corebit_and and_inst179(.in0(and_inst178_out), .in1(Module_0_inst180_valid_down), .out(and_inst179_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(Module_0_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst180(.in0(and_inst179_out), .in1(Module_0_inst181_valid_down), .out(and_inst180_out));
corebit_and and_inst181(.in0(and_inst180_out), .in1(Module_0_inst182_valid_down), .out(and_inst181_out));
corebit_and and_inst182(.in0(and_inst181_out), .in1(Module_0_inst183_valid_down), .out(and_inst182_out));
corebit_and and_inst183(.in0(and_inst182_out), .in1(Module_0_inst184_valid_down), .out(and_inst183_out));
corebit_and and_inst184(.in0(and_inst183_out), .in1(Module_0_inst185_valid_down), .out(and_inst184_out));
corebit_and and_inst185(.in0(and_inst184_out), .in1(Module_0_inst186_valid_down), .out(and_inst185_out));
corebit_and and_inst186(.in0(and_inst185_out), .in1(Module_0_inst187_valid_down), .out(and_inst186_out));
corebit_and and_inst187(.in0(and_inst186_out), .in1(Module_0_inst188_valid_down), .out(and_inst187_out));
corebit_and and_inst188(.in0(and_inst187_out), .in1(Module_0_inst189_valid_down), .out(and_inst188_out));
corebit_and and_inst189(.in0(and_inst188_out), .in1(Module_0_inst190_valid_down), .out(and_inst189_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(Module_0_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst190(.in0(and_inst189_out), .in1(Module_0_inst191_valid_down), .out(and_inst190_out));
corebit_and and_inst191(.in0(and_inst190_out), .in1(Module_0_inst192_valid_down), .out(and_inst191_out));
corebit_and and_inst192(.in0(and_inst191_out), .in1(Module_0_inst193_valid_down), .out(and_inst192_out));
corebit_and and_inst193(.in0(and_inst192_out), .in1(Module_0_inst194_valid_down), .out(and_inst193_out));
corebit_and and_inst194(.in0(and_inst193_out), .in1(Module_0_inst195_valid_down), .out(and_inst194_out));
corebit_and and_inst195(.in0(and_inst194_out), .in1(Module_0_inst196_valid_down), .out(and_inst195_out));
corebit_and and_inst196(.in0(and_inst195_out), .in1(Module_0_inst197_valid_down), .out(and_inst196_out));
corebit_and and_inst197(.in0(and_inst196_out), .in1(Module_0_inst198_valid_down), .out(and_inst197_out));
corebit_and and_inst198(.in0(and_inst197_out), .in1(Module_0_inst199_valid_down), .out(and_inst198_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Module_0_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(Module_0_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(Module_0_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(Module_0_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(Module_0_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(Module_0_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(Module_0_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst26(.in0(and_inst25_out), .in1(Module_0_inst27_valid_down), .out(and_inst26_out));
corebit_and and_inst27(.in0(and_inst26_out), .in1(Module_0_inst28_valid_down), .out(and_inst27_out));
corebit_and and_inst28(.in0(and_inst27_out), .in1(Module_0_inst29_valid_down), .out(and_inst28_out));
corebit_and and_inst29(.in0(and_inst28_out), .in1(Module_0_inst30_valid_down), .out(and_inst29_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Module_0_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst30(.in0(and_inst29_out), .in1(Module_0_inst31_valid_down), .out(and_inst30_out));
corebit_and and_inst31(.in0(and_inst30_out), .in1(Module_0_inst32_valid_down), .out(and_inst31_out));
corebit_and and_inst32(.in0(and_inst31_out), .in1(Module_0_inst33_valid_down), .out(and_inst32_out));
corebit_and and_inst33(.in0(and_inst32_out), .in1(Module_0_inst34_valid_down), .out(and_inst33_out));
corebit_and and_inst34(.in0(and_inst33_out), .in1(Module_0_inst35_valid_down), .out(and_inst34_out));
corebit_and and_inst35(.in0(and_inst34_out), .in1(Module_0_inst36_valid_down), .out(and_inst35_out));
corebit_and and_inst36(.in0(and_inst35_out), .in1(Module_0_inst37_valid_down), .out(and_inst36_out));
corebit_and and_inst37(.in0(and_inst36_out), .in1(Module_0_inst38_valid_down), .out(and_inst37_out));
corebit_and and_inst38(.in0(and_inst37_out), .in1(Module_0_inst39_valid_down), .out(and_inst38_out));
corebit_and and_inst39(.in0(and_inst38_out), .in1(Module_0_inst40_valid_down), .out(and_inst39_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Module_0_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst40(.in0(and_inst39_out), .in1(Module_0_inst41_valid_down), .out(and_inst40_out));
corebit_and and_inst41(.in0(and_inst40_out), .in1(Module_0_inst42_valid_down), .out(and_inst41_out));
corebit_and and_inst42(.in0(and_inst41_out), .in1(Module_0_inst43_valid_down), .out(and_inst42_out));
corebit_and and_inst43(.in0(and_inst42_out), .in1(Module_0_inst44_valid_down), .out(and_inst43_out));
corebit_and and_inst44(.in0(and_inst43_out), .in1(Module_0_inst45_valid_down), .out(and_inst44_out));
corebit_and and_inst45(.in0(and_inst44_out), .in1(Module_0_inst46_valid_down), .out(and_inst45_out));
corebit_and and_inst46(.in0(and_inst45_out), .in1(Module_0_inst47_valid_down), .out(and_inst46_out));
corebit_and and_inst47(.in0(and_inst46_out), .in1(Module_0_inst48_valid_down), .out(and_inst47_out));
corebit_and and_inst48(.in0(and_inst47_out), .in1(Module_0_inst49_valid_down), .out(and_inst48_out));
corebit_and and_inst49(.in0(and_inst48_out), .in1(Module_0_inst50_valid_down), .out(and_inst49_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Module_0_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst50(.in0(and_inst49_out), .in1(Module_0_inst51_valid_down), .out(and_inst50_out));
corebit_and and_inst51(.in0(and_inst50_out), .in1(Module_0_inst52_valid_down), .out(and_inst51_out));
corebit_and and_inst52(.in0(and_inst51_out), .in1(Module_0_inst53_valid_down), .out(and_inst52_out));
corebit_and and_inst53(.in0(and_inst52_out), .in1(Module_0_inst54_valid_down), .out(and_inst53_out));
corebit_and and_inst54(.in0(and_inst53_out), .in1(Module_0_inst55_valid_down), .out(and_inst54_out));
corebit_and and_inst55(.in0(and_inst54_out), .in1(Module_0_inst56_valid_down), .out(and_inst55_out));
corebit_and and_inst56(.in0(and_inst55_out), .in1(Module_0_inst57_valid_down), .out(and_inst56_out));
corebit_and and_inst57(.in0(and_inst56_out), .in1(Module_0_inst58_valid_down), .out(and_inst57_out));
corebit_and and_inst58(.in0(and_inst57_out), .in1(Module_0_inst59_valid_down), .out(and_inst58_out));
corebit_and and_inst59(.in0(and_inst58_out), .in1(Module_0_inst60_valid_down), .out(and_inst59_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Module_0_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst60(.in0(and_inst59_out), .in1(Module_0_inst61_valid_down), .out(and_inst60_out));
corebit_and and_inst61(.in0(and_inst60_out), .in1(Module_0_inst62_valid_down), .out(and_inst61_out));
corebit_and and_inst62(.in0(and_inst61_out), .in1(Module_0_inst63_valid_down), .out(and_inst62_out));
corebit_and and_inst63(.in0(and_inst62_out), .in1(Module_0_inst64_valid_down), .out(and_inst63_out));
corebit_and and_inst64(.in0(and_inst63_out), .in1(Module_0_inst65_valid_down), .out(and_inst64_out));
corebit_and and_inst65(.in0(and_inst64_out), .in1(Module_0_inst66_valid_down), .out(and_inst65_out));
corebit_and and_inst66(.in0(and_inst65_out), .in1(Module_0_inst67_valid_down), .out(and_inst66_out));
corebit_and and_inst67(.in0(and_inst66_out), .in1(Module_0_inst68_valid_down), .out(and_inst67_out));
corebit_and and_inst68(.in0(and_inst67_out), .in1(Module_0_inst69_valid_down), .out(and_inst68_out));
corebit_and and_inst69(.in0(and_inst68_out), .in1(Module_0_inst70_valid_down), .out(and_inst69_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Module_0_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst70(.in0(and_inst69_out), .in1(Module_0_inst71_valid_down), .out(and_inst70_out));
corebit_and and_inst71(.in0(and_inst70_out), .in1(Module_0_inst72_valid_down), .out(and_inst71_out));
corebit_and and_inst72(.in0(and_inst71_out), .in1(Module_0_inst73_valid_down), .out(and_inst72_out));
corebit_and and_inst73(.in0(and_inst72_out), .in1(Module_0_inst74_valid_down), .out(and_inst73_out));
corebit_and and_inst74(.in0(and_inst73_out), .in1(Module_0_inst75_valid_down), .out(and_inst74_out));
corebit_and and_inst75(.in0(and_inst74_out), .in1(Module_0_inst76_valid_down), .out(and_inst75_out));
corebit_and and_inst76(.in0(and_inst75_out), .in1(Module_0_inst77_valid_down), .out(and_inst76_out));
corebit_and and_inst77(.in0(and_inst76_out), .in1(Module_0_inst78_valid_down), .out(and_inst77_out));
corebit_and and_inst78(.in0(and_inst77_out), .in1(Module_0_inst79_valid_down), .out(and_inst78_out));
corebit_and and_inst79(.in0(and_inst78_out), .in1(Module_0_inst80_valid_down), .out(and_inst79_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(Module_0_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst80(.in0(and_inst79_out), .in1(Module_0_inst81_valid_down), .out(and_inst80_out));
corebit_and and_inst81(.in0(and_inst80_out), .in1(Module_0_inst82_valid_down), .out(and_inst81_out));
corebit_and and_inst82(.in0(and_inst81_out), .in1(Module_0_inst83_valid_down), .out(and_inst82_out));
corebit_and and_inst83(.in0(and_inst82_out), .in1(Module_0_inst84_valid_down), .out(and_inst83_out));
corebit_and and_inst84(.in0(and_inst83_out), .in1(Module_0_inst85_valid_down), .out(and_inst84_out));
corebit_and and_inst85(.in0(and_inst84_out), .in1(Module_0_inst86_valid_down), .out(and_inst85_out));
corebit_and and_inst86(.in0(and_inst85_out), .in1(Module_0_inst87_valid_down), .out(and_inst86_out));
corebit_and and_inst87(.in0(and_inst86_out), .in1(Module_0_inst88_valid_down), .out(and_inst87_out));
corebit_and and_inst88(.in0(and_inst87_out), .in1(Module_0_inst89_valid_down), .out(and_inst88_out));
corebit_and and_inst89(.in0(and_inst88_out), .in1(Module_0_inst90_valid_down), .out(and_inst89_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(Module_0_inst10_valid_down), .out(and_inst9_out));
corebit_and and_inst90(.in0(and_inst89_out), .in1(Module_0_inst91_valid_down), .out(and_inst90_out));
corebit_and and_inst91(.in0(and_inst90_out), .in1(Module_0_inst92_valid_down), .out(and_inst91_out));
corebit_and and_inst92(.in0(and_inst91_out), .in1(Module_0_inst93_valid_down), .out(and_inst92_out));
corebit_and and_inst93(.in0(and_inst92_out), .in1(Module_0_inst94_valid_down), .out(and_inst93_out));
corebit_and and_inst94(.in0(and_inst93_out), .in1(Module_0_inst95_valid_down), .out(and_inst94_out));
corebit_and and_inst95(.in0(and_inst94_out), .in1(Module_0_inst96_valid_down), .out(and_inst95_out));
corebit_and and_inst96(.in0(and_inst95_out), .in1(Module_0_inst97_valid_down), .out(and_inst96_out));
corebit_and and_inst97(.in0(and_inst96_out), .in1(Module_0_inst98_valid_down), .out(and_inst97_out));
corebit_and and_inst98(.in0(and_inst97_out), .in1(Module_0_inst99_valid_down), .out(and_inst98_out));
corebit_and and_inst99(.in0(and_inst98_out), .in1(Module_0_inst100_valid_down), .out(and_inst99_out));
assign O_0 = Module_0_inst0_O;
assign O_1 = Module_0_inst1_O;
assign O_10 = Module_0_inst10_O;
assign O_100 = Module_0_inst100_O;
assign O_101 = Module_0_inst101_O;
assign O_102 = Module_0_inst102_O;
assign O_103 = Module_0_inst103_O;
assign O_104 = Module_0_inst104_O;
assign O_105 = Module_0_inst105_O;
assign O_106 = Module_0_inst106_O;
assign O_107 = Module_0_inst107_O;
assign O_108 = Module_0_inst108_O;
assign O_109 = Module_0_inst109_O;
assign O_11 = Module_0_inst11_O;
assign O_110 = Module_0_inst110_O;
assign O_111 = Module_0_inst111_O;
assign O_112 = Module_0_inst112_O;
assign O_113 = Module_0_inst113_O;
assign O_114 = Module_0_inst114_O;
assign O_115 = Module_0_inst115_O;
assign O_116 = Module_0_inst116_O;
assign O_117 = Module_0_inst117_O;
assign O_118 = Module_0_inst118_O;
assign O_119 = Module_0_inst119_O;
assign O_12 = Module_0_inst12_O;
assign O_120 = Module_0_inst120_O;
assign O_121 = Module_0_inst121_O;
assign O_122 = Module_0_inst122_O;
assign O_123 = Module_0_inst123_O;
assign O_124 = Module_0_inst124_O;
assign O_125 = Module_0_inst125_O;
assign O_126 = Module_0_inst126_O;
assign O_127 = Module_0_inst127_O;
assign O_128 = Module_0_inst128_O;
assign O_129 = Module_0_inst129_O;
assign O_13 = Module_0_inst13_O;
assign O_130 = Module_0_inst130_O;
assign O_131 = Module_0_inst131_O;
assign O_132 = Module_0_inst132_O;
assign O_133 = Module_0_inst133_O;
assign O_134 = Module_0_inst134_O;
assign O_135 = Module_0_inst135_O;
assign O_136 = Module_0_inst136_O;
assign O_137 = Module_0_inst137_O;
assign O_138 = Module_0_inst138_O;
assign O_139 = Module_0_inst139_O;
assign O_14 = Module_0_inst14_O;
assign O_140 = Module_0_inst140_O;
assign O_141 = Module_0_inst141_O;
assign O_142 = Module_0_inst142_O;
assign O_143 = Module_0_inst143_O;
assign O_144 = Module_0_inst144_O;
assign O_145 = Module_0_inst145_O;
assign O_146 = Module_0_inst146_O;
assign O_147 = Module_0_inst147_O;
assign O_148 = Module_0_inst148_O;
assign O_149 = Module_0_inst149_O;
assign O_15 = Module_0_inst15_O;
assign O_150 = Module_0_inst150_O;
assign O_151 = Module_0_inst151_O;
assign O_152 = Module_0_inst152_O;
assign O_153 = Module_0_inst153_O;
assign O_154 = Module_0_inst154_O;
assign O_155 = Module_0_inst155_O;
assign O_156 = Module_0_inst156_O;
assign O_157 = Module_0_inst157_O;
assign O_158 = Module_0_inst158_O;
assign O_159 = Module_0_inst159_O;
assign O_16 = Module_0_inst16_O;
assign O_160 = Module_0_inst160_O;
assign O_161 = Module_0_inst161_O;
assign O_162 = Module_0_inst162_O;
assign O_163 = Module_0_inst163_O;
assign O_164 = Module_0_inst164_O;
assign O_165 = Module_0_inst165_O;
assign O_166 = Module_0_inst166_O;
assign O_167 = Module_0_inst167_O;
assign O_168 = Module_0_inst168_O;
assign O_169 = Module_0_inst169_O;
assign O_17 = Module_0_inst17_O;
assign O_170 = Module_0_inst170_O;
assign O_171 = Module_0_inst171_O;
assign O_172 = Module_0_inst172_O;
assign O_173 = Module_0_inst173_O;
assign O_174 = Module_0_inst174_O;
assign O_175 = Module_0_inst175_O;
assign O_176 = Module_0_inst176_O;
assign O_177 = Module_0_inst177_O;
assign O_178 = Module_0_inst178_O;
assign O_179 = Module_0_inst179_O;
assign O_18 = Module_0_inst18_O;
assign O_180 = Module_0_inst180_O;
assign O_181 = Module_0_inst181_O;
assign O_182 = Module_0_inst182_O;
assign O_183 = Module_0_inst183_O;
assign O_184 = Module_0_inst184_O;
assign O_185 = Module_0_inst185_O;
assign O_186 = Module_0_inst186_O;
assign O_187 = Module_0_inst187_O;
assign O_188 = Module_0_inst188_O;
assign O_189 = Module_0_inst189_O;
assign O_19 = Module_0_inst19_O;
assign O_190 = Module_0_inst190_O;
assign O_191 = Module_0_inst191_O;
assign O_192 = Module_0_inst192_O;
assign O_193 = Module_0_inst193_O;
assign O_194 = Module_0_inst194_O;
assign O_195 = Module_0_inst195_O;
assign O_196 = Module_0_inst196_O;
assign O_197 = Module_0_inst197_O;
assign O_198 = Module_0_inst198_O;
assign O_199 = Module_0_inst199_O;
assign O_2 = Module_0_inst2_O;
assign O_20 = Module_0_inst20_O;
assign O_21 = Module_0_inst21_O;
assign O_22 = Module_0_inst22_O;
assign O_23 = Module_0_inst23_O;
assign O_24 = Module_0_inst24_O;
assign O_25 = Module_0_inst25_O;
assign O_26 = Module_0_inst26_O;
assign O_27 = Module_0_inst27_O;
assign O_28 = Module_0_inst28_O;
assign O_29 = Module_0_inst29_O;
assign O_3 = Module_0_inst3_O;
assign O_30 = Module_0_inst30_O;
assign O_31 = Module_0_inst31_O;
assign O_32 = Module_0_inst32_O;
assign O_33 = Module_0_inst33_O;
assign O_34 = Module_0_inst34_O;
assign O_35 = Module_0_inst35_O;
assign O_36 = Module_0_inst36_O;
assign O_37 = Module_0_inst37_O;
assign O_38 = Module_0_inst38_O;
assign O_39 = Module_0_inst39_O;
assign O_4 = Module_0_inst4_O;
assign O_40 = Module_0_inst40_O;
assign O_41 = Module_0_inst41_O;
assign O_42 = Module_0_inst42_O;
assign O_43 = Module_0_inst43_O;
assign O_44 = Module_0_inst44_O;
assign O_45 = Module_0_inst45_O;
assign O_46 = Module_0_inst46_O;
assign O_47 = Module_0_inst47_O;
assign O_48 = Module_0_inst48_O;
assign O_49 = Module_0_inst49_O;
assign O_5 = Module_0_inst5_O;
assign O_50 = Module_0_inst50_O;
assign O_51 = Module_0_inst51_O;
assign O_52 = Module_0_inst52_O;
assign O_53 = Module_0_inst53_O;
assign O_54 = Module_0_inst54_O;
assign O_55 = Module_0_inst55_O;
assign O_56 = Module_0_inst56_O;
assign O_57 = Module_0_inst57_O;
assign O_58 = Module_0_inst58_O;
assign O_59 = Module_0_inst59_O;
assign O_6 = Module_0_inst6_O;
assign O_60 = Module_0_inst60_O;
assign O_61 = Module_0_inst61_O;
assign O_62 = Module_0_inst62_O;
assign O_63 = Module_0_inst63_O;
assign O_64 = Module_0_inst64_O;
assign O_65 = Module_0_inst65_O;
assign O_66 = Module_0_inst66_O;
assign O_67 = Module_0_inst67_O;
assign O_68 = Module_0_inst68_O;
assign O_69 = Module_0_inst69_O;
assign O_7 = Module_0_inst7_O;
assign O_70 = Module_0_inst70_O;
assign O_71 = Module_0_inst71_O;
assign O_72 = Module_0_inst72_O;
assign O_73 = Module_0_inst73_O;
assign O_74 = Module_0_inst74_O;
assign O_75 = Module_0_inst75_O;
assign O_76 = Module_0_inst76_O;
assign O_77 = Module_0_inst77_O;
assign O_78 = Module_0_inst78_O;
assign O_79 = Module_0_inst79_O;
assign O_8 = Module_0_inst8_O;
assign O_80 = Module_0_inst80_O;
assign O_81 = Module_0_inst81_O;
assign O_82 = Module_0_inst82_O;
assign O_83 = Module_0_inst83_O;
assign O_84 = Module_0_inst84_O;
assign O_85 = Module_0_inst85_O;
assign O_86 = Module_0_inst86_O;
assign O_87 = Module_0_inst87_O;
assign O_88 = Module_0_inst88_O;
assign O_89 = Module_0_inst89_O;
assign O_9 = Module_0_inst9_O;
assign O_90 = Module_0_inst90_O;
assign O_91 = Module_0_inst91_O;
assign O_92 = Module_0_inst92_O;
assign O_93 = Module_0_inst93_O;
assign O_94 = Module_0_inst94_O;
assign O_95 = Module_0_inst95_O;
assign O_96 = Module_0_inst96_O;
assign O_97 = Module_0_inst97_O;
assign O_98 = Module_0_inst98_O;
assign O_99 = Module_0_inst99_O;
assign valid_down = and_inst198_out;
endmodule

module top (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_100;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_101;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_102;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_103;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_104;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_105;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_106;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_107;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_108;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_109;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_110;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_111;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_112;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_113;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_114;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_115;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_116;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_117;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_118;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_119;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_120;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_121;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_122;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_123;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_124;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_125;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_126;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_127;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_128;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_129;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_130;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_131;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_132;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_133;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_134;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_135;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_136;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_137;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_138;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_139;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_140;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_141;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_142;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_143;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_144;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_145;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_146;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_147;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_148;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_149;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_150;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_151;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_152;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_153;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_154;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_155;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_156;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_157;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_158;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_159;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_160;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_161;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_162;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_163;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_164;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_165;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_166;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_167;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_168;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_169;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_170;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_171;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_172;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_173;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_174;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_175;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_176;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_177;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_178;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_179;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_180;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_181;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_182;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_183;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_184;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_185;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_186;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_187;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_188;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_189;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_190;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_191;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_192;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_193;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_194;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_195;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_196;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_197;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_198;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_199;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_40;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_41;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_42;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_43;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_44;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_45;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_46;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_47;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_48;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_49;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_50;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_51;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_52;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_53;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_54;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_55;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_56;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_57;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_58;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_59;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_60;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_61;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_62;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_63;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_64;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_65;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_66;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_67;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_68;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_69;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_70;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_71;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_72;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_73;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_74;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_75;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_76;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_77;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_78;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_79;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_80;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_81;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_82;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_83;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_84;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_85;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_86;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_87;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_88;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_89;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_90;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_91;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_92;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_93;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_94;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_95;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_96;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_97;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_98;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_99;
wire NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_100(I_100), .I_101(I_101), .I_102(I_102), .I_103(I_103), .I_104(I_104), .I_105(I_105), .I_106(I_106), .I_107(I_107), .I_108(I_108), .I_109(I_109), .I_11(I_11), .I_110(I_110), .I_111(I_111), .I_112(I_112), .I_113(I_113), .I_114(I_114), .I_115(I_115), .I_116(I_116), .I_117(I_117), .I_118(I_118), .I_119(I_119), .I_12(I_12), .I_120(I_120), .I_121(I_121), .I_122(I_122), .I_123(I_123), .I_124(I_124), .I_125(I_125), .I_126(I_126), .I_127(I_127), .I_128(I_128), .I_129(I_129), .I_13(I_13), .I_130(I_130), .I_131(I_131), .I_132(I_132), .I_133(I_133), .I_134(I_134), .I_135(I_135), .I_136(I_136), .I_137(I_137), .I_138(I_138), .I_139(I_139), .I_14(I_14), .I_140(I_140), .I_141(I_141), .I_142(I_142), .I_143(I_143), .I_144(I_144), .I_145(I_145), .I_146(I_146), .I_147(I_147), .I_148(I_148), .I_149(I_149), .I_15(I_15), .I_150(I_150), .I_151(I_151), .I_152(I_152), .I_153(I_153), .I_154(I_154), .I_155(I_155), .I_156(I_156), .I_157(I_157), .I_158(I_158), .I_159(I_159), .I_16(I_16), .I_160(I_160), .I_161(I_161), .I_162(I_162), .I_163(I_163), .I_164(I_164), .I_165(I_165), .I_166(I_166), .I_167(I_167), .I_168(I_168), .I_169(I_169), .I_17(I_17), .I_170(I_170), .I_171(I_171), .I_172(I_172), .I_173(I_173), .I_174(I_174), .I_175(I_175), .I_176(I_176), .I_177(I_177), .I_178(I_178), .I_179(I_179), .I_18(I_18), .I_180(I_180), .I_181(I_181), .I_182(I_182), .I_183(I_183), .I_184(I_184), .I_185(I_185), .I_186(I_186), .I_187(I_187), .I_188(I_188), .I_189(I_189), .I_19(I_19), .I_190(I_190), .I_191(I_191), .I_192(I_192), .I_193(I_193), .I_194(I_194), .I_195(I_195), .I_196(I_196), .I_197(I_197), .I_198(I_198), .I_199(I_199), .I_2(I_2), .I_20(I_20), .I_21(I_21), .I_22(I_22), .I_23(I_23), .I_24(I_24), .I_25(I_25), .I_26(I_26), .I_27(I_27), .I_28(I_28), .I_29(I_29), .I_3(I_3), .I_30(I_30), .I_31(I_31), .I_32(I_32), .I_33(I_33), .I_34(I_34), .I_35(I_35), .I_36(I_36), .I_37(I_37), .I_38(I_38), .I_39(I_39), .I_4(I_4), .I_40(I_40), .I_41(I_41), .I_42(I_42), .I_43(I_43), .I_44(I_44), .I_45(I_45), .I_46(I_46), .I_47(I_47), .I_48(I_48), .I_49(I_49), .I_5(I_5), .I_50(I_50), .I_51(I_51), .I_52(I_52), .I_53(I_53), .I_54(I_54), .I_55(I_55), .I_56(I_56), .I_57(I_57), .I_58(I_58), .I_59(I_59), .I_6(I_6), .I_60(I_60), .I_61(I_61), .I_62(I_62), .I_63(I_63), .I_64(I_64), .I_65(I_65), .I_66(I_66), .I_67(I_67), .I_68(I_68), .I_69(I_69), .I_7(I_7), .I_70(I_70), .I_71(I_71), .I_72(I_72), .I_73(I_73), .I_74(I_74), .I_75(I_75), .I_76(I_76), .I_77(I_77), .I_78(I_78), .I_79(I_79), .I_8(I_8), .I_80(I_80), .I_81(I_81), .I_82(I_82), .I_83(I_83), .I_84(I_84), .I_85(I_85), .I_86(I_86), .I_87(I_87), .I_88(I_88), .I_89(I_89), .I_9(I_9), .I_90(I_90), .I_91(I_91), .I_92(I_92), .I_93(I_93), .I_94(I_94), .I_95(I_95), .I_96(I_96), .I_97(I_97), .I_98(I_98), .I_99(I_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .I_1(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .I_10(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .I_100(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_100), .I_101(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_101), .I_102(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_102), .I_103(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_103), .I_104(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_104), .I_105(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_105), .I_106(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_106), .I_107(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_107), .I_108(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_108), .I_109(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_109), .I_11(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .I_110(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_110), .I_111(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_111), .I_112(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_112), .I_113(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_113), .I_114(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_114), .I_115(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_115), .I_116(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_116), .I_117(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_117), .I_118(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_118), .I_119(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_119), .I_12(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .I_120(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_120), .I_121(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_121), .I_122(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_122), .I_123(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_123), .I_124(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_124), .I_125(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_125), .I_126(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_126), .I_127(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_127), .I_128(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_128), .I_129(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_129), .I_13(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .I_130(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_130), .I_131(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_131), .I_132(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_132), .I_133(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_133), .I_134(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_134), .I_135(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_135), .I_136(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_136), .I_137(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_137), .I_138(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_138), .I_139(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_139), .I_14(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .I_140(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_140), .I_141(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_141), .I_142(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_142), .I_143(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_143), .I_144(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_144), .I_145(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_145), .I_146(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_146), .I_147(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_147), .I_148(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_148), .I_149(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_149), .I_15(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .I_150(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_150), .I_151(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_151), .I_152(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_152), .I_153(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_153), .I_154(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_154), .I_155(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_155), .I_156(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_156), .I_157(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_157), .I_158(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_158), .I_159(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_159), .I_16(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .I_160(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_160), .I_161(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_161), .I_162(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_162), .I_163(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_163), .I_164(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_164), .I_165(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_165), .I_166(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_166), .I_167(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_167), .I_168(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_168), .I_169(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_169), .I_17(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .I_170(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_170), .I_171(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_171), .I_172(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_172), .I_173(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_173), .I_174(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_174), .I_175(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_175), .I_176(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_176), .I_177(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_177), .I_178(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_178), .I_179(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_179), .I_18(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .I_180(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_180), .I_181(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_181), .I_182(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_182), .I_183(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_183), .I_184(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_184), .I_185(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_185), .I_186(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_186), .I_187(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_187), .I_188(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_188), .I_189(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_189), .I_19(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .I_190(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_190), .I_191(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_191), .I_192(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_192), .I_193(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_193), .I_194(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_194), .I_195(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_195), .I_196(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_196), .I_197(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_197), .I_198(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_198), .I_199(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_199), .I_2(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .I_20(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .I_21(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .I_22(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .I_23(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .I_24(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .I_25(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .I_26(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .I_27(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .I_28(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .I_29(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .I_3(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .I_30(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .I_31(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .I_32(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .I_33(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .I_34(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .I_35(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .I_36(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .I_37(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .I_38(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .I_39(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .I_4(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .I_40(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_40), .I_41(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_41), .I_42(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_42), .I_43(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_43), .I_44(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_44), .I_45(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_45), .I_46(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_46), .I_47(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_47), .I_48(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_48), .I_49(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_49), .I_5(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .I_50(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_50), .I_51(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_51), .I_52(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_52), .I_53(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_53), .I_54(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_54), .I_55(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_55), .I_56(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_56), .I_57(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_57), .I_58(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_58), .I_59(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_59), .I_6(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .I_60(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_60), .I_61(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_61), .I_62(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_62), .I_63(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_63), .I_64(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_64), .I_65(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_65), .I_66(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_66), .I_67(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_67), .I_68(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_68), .I_69(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_69), .I_7(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .I_70(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_70), .I_71(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_71), .I_72(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_72), .I_73(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_73), .I_74(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_74), .I_75(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_75), .I_76(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_76), .I_77(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_77), .I_78(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_78), .I_79(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_79), .I_8(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .I_80(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_80), .I_81(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_81), .I_82(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_82), .I_83(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_83), .I_84(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_84), .I_85(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_85), .I_86(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_86), .I_87(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_87), .I_88(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_88), .I_89(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_89), .I_9(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .I_90(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_90), .I_91(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_91), .I_92(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_92), .I_93(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_93), .I_94(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_94), .I_95(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_95), .I_96(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_96), .I_97(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_97), .I_98(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_98), .I_99(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down));
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .I_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .I_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .I_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_100), .I_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_101), .I_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_102), .I_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_103), .I_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_104), .I_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_105), .I_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_106), .I_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_107), .I_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_108), .I_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_109), .I_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .I_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_110), .I_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_111), .I_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_112), .I_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_113), .I_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_114), .I_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_115), .I_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_116), .I_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_117), .I_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_118), .I_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_119), .I_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .I_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_120), .I_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_121), .I_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_122), .I_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_123), .I_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_124), .I_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_125), .I_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_126), .I_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_127), .I_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_128), .I_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_129), .I_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .I_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_130), .I_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_131), .I_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_132), .I_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_133), .I_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_134), .I_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_135), .I_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_136), .I_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_137), .I_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_138), .I_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_139), .I_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .I_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_140), .I_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_141), .I_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_142), .I_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_143), .I_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_144), .I_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_145), .I_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_146), .I_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_147), .I_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_148), .I_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_149), .I_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .I_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_150), .I_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_151), .I_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_152), .I_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_153), .I_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_154), .I_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_155), .I_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_156), .I_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_157), .I_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_158), .I_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_159), .I_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .I_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_160), .I_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_161), .I_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_162), .I_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_163), .I_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_164), .I_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_165), .I_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_166), .I_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_167), .I_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_168), .I_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_169), .I_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .I_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_170), .I_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_171), .I_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_172), .I_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_173), .I_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_174), .I_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_175), .I_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_176), .I_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_177), .I_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_178), .I_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_179), .I_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .I_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_180), .I_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_181), .I_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_182), .I_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_183), .I_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_184), .I_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_185), .I_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_186), .I_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_187), .I_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_188), .I_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_189), .I_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .I_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_190), .I_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_191), .I_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_192), .I_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_193), .I_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_194), .I_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_195), .I_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_196), .I_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_197), .I_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_198), .I_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_199), .I_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .I_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20), .I_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21), .I_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22), .I_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23), .I_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24), .I_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25), .I_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26), .I_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27), .I_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28), .I_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29), .I_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .I_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30), .I_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31), .I_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32), .I_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33), .I_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34), .I_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35), .I_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36), .I_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37), .I_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38), .I_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39), .I_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .I_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_40), .I_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_41), .I_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_42), .I_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_43), .I_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_44), .I_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_45), .I_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_46), .I_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_47), .I_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_48), .I_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_49), .I_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .I_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_50), .I_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_51), .I_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_52), .I_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_53), .I_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_54), .I_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_55), .I_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_56), .I_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_57), .I_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_58), .I_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_59), .I_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .I_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_60), .I_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_61), .I_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_62), .I_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_63), .I_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_64), .I_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_65), .I_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_66), .I_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_67), .I_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_68), .I_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_69), .I_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .I_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_70), .I_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_71), .I_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_72), .I_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_73), .I_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_74), .I_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_75), .I_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_76), .I_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_77), .I_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_78), .I_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_79), .I_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .I_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_80), .I_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_81), .I_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_82), .I_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_83), .I_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_84), .I_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_85), .I_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_86), .I_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_87), .I_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_88), .I_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_89), .I_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .I_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_90), .I_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_91), .I_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_92), .I_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_93), .I_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_94), .I_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_95), .I_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_96), .I_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_97), .I_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_98), .I_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0(.CLK(CLK), .I_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .I_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_100), .I_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_101), .I_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_102), .I_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_103), .I_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_104), .I_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_105), .I_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_106), .I_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_107), .I_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_108), .I_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_109), .I_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .I_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_110), .I_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_111), .I_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_112), .I_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_113), .I_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_114), .I_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_115), .I_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_116), .I_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_117), .I_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_118), .I_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_119), .I_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .I_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_120), .I_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_121), .I_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_122), .I_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_123), .I_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_124), .I_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_125), .I_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_126), .I_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_127), .I_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_128), .I_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_129), .I_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .I_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_130), .I_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_131), .I_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_132), .I_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_133), .I_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_134), .I_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_135), .I_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_136), .I_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_137), .I_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_138), .I_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_139), .I_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .I_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_140), .I_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_141), .I_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_142), .I_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_143), .I_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_144), .I_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_145), .I_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_146), .I_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_147), .I_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_148), .I_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_149), .I_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .I_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_150), .I_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_151), .I_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_152), .I_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_153), .I_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_154), .I_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_155), .I_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_156), .I_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_157), .I_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_158), .I_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_159), .I_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .I_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_160), .I_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_161), .I_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_162), .I_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_163), .I_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_164), .I_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_165), .I_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_166), .I_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_167), .I_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_168), .I_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_169), .I_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .I_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_170), .I_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_171), .I_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_172), .I_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_173), .I_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_174), .I_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_175), .I_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_176), .I_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_177), .I_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_178), .I_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_179), .I_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .I_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_180), .I_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_181), .I_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_182), .I_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_183), .I_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_184), .I_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_185), .I_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_186), .I_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_187), .I_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_188), .I_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_189), .I_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .I_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_190), .I_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_191), .I_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_192), .I_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_193), .I_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_194), .I_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_195), .I_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_196), .I_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_197), .I_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_198), .I_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_199), .I_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .I_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20), .I_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21), .I_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22), .I_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23), .I_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24), .I_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25), .I_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26), .I_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27), .I_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28), .I_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29), .I_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .I_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30), .I_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31), .I_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32), .I_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33), .I_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34), .I_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35), .I_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36), .I_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37), .I_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38), .I_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39), .I_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .I_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_40), .I_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_41), .I_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_42), .I_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_43), .I_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_44), .I_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_45), .I_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_46), .I_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_47), .I_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_48), .I_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_49), .I_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .I_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_50), .I_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_51), .I_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_52), .I_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_53), .I_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_54), .I_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_55), .I_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_56), .I_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_57), .I_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_58), .I_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_59), .I_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .I_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_60), .I_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_61), .I_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_62), .I_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_63), .I_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_64), .I_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_65), .I_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_66), .I_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_67), .I_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_68), .I_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_69), .I_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .I_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_70), .I_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_71), .I_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_72), .I_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_73), .I_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_74), .I_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_75), .I_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_76), .I_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_77), .I_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_78), .I_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_79), .I_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .I_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_80), .I_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_81), .I_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_82), .I_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_83), .I_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_84), .I_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_85), .I_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_86), .I_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_87), .I_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_88), .I_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_89), .I_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .I_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_90), .I_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_91), .I_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_92), .I_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_93), .I_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_94), .I_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_95), .I_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_96), .I_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_97), .I_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_98), .I_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_99), .O_0(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_10(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .O_100(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_100), .O_101(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_101), .O_102(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_102), .O_103(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_103), .O_104(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_104), .O_105(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_105), .O_106(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_106), .O_107(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_107), .O_108(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_108), .O_109(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_109), .O_11(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .O_110(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_110), .O_111(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_111), .O_112(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_112), .O_113(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_113), .O_114(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_114), .O_115(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_115), .O_116(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_116), .O_117(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_117), .O_118(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_118), .O_119(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_119), .O_12(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .O_120(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_120), .O_121(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_121), .O_122(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_122), .O_123(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_123), .O_124(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_124), .O_125(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_125), .O_126(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_126), .O_127(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_127), .O_128(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_128), .O_129(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_129), .O_13(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .O_130(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_130), .O_131(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_131), .O_132(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_132), .O_133(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_133), .O_134(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_134), .O_135(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_135), .O_136(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_136), .O_137(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_137), .O_138(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_138), .O_139(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_139), .O_14(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .O_140(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_140), .O_141(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_141), .O_142(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_142), .O_143(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_143), .O_144(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_144), .O_145(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_145), .O_146(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_146), .O_147(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_147), .O_148(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_148), .O_149(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_149), .O_15(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .O_150(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_150), .O_151(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_151), .O_152(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_152), .O_153(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_153), .O_154(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_154), .O_155(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_155), .O_156(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_156), .O_157(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_157), .O_158(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_158), .O_159(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_159), .O_16(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .O_160(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_160), .O_161(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_161), .O_162(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_162), .O_163(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_163), .O_164(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_164), .O_165(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_165), .O_166(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_166), .O_167(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_167), .O_168(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_168), .O_169(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_169), .O_17(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .O_170(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_170), .O_171(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_171), .O_172(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_172), .O_173(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_173), .O_174(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_174), .O_175(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_175), .O_176(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_176), .O_177(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_177), .O_178(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_178), .O_179(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_179), .O_18(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .O_180(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_180), .O_181(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_181), .O_182(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_182), .O_183(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_183), .O_184(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_184), .O_185(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_185), .O_186(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_186), .O_187(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_187), .O_188(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_188), .O_189(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_189), .O_19(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .O_190(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_190), .O_191(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_191), .O_192(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_192), .O_193(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_193), .O_194(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_194), .O_195(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_195), .O_196(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_196), .O_197(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_197), .O_198(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_198), .O_199(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_199), .O_2(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .O_20(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .O_21(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .O_22(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .O_23(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .O_24(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .O_25(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .O_26(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .O_27(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .O_28(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .O_29(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .O_3(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .O_30(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .O_31(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .O_32(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .O_33(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .O_34(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .O_35(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .O_36(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .O_37(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .O_38(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .O_39(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .O_4(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .O_40(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_40), .O_41(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_41), .O_42(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_42), .O_43(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_43), .O_44(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_44), .O_45(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_45), .O_46(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_46), .O_47(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_47), .O_48(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_48), .O_49(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_49), .O_5(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .O_50(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_50), .O_51(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_51), .O_52(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_52), .O_53(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_53), .O_54(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_54), .O_55(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_55), .O_56(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_56), .O_57(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_57), .O_58(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_58), .O_59(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_59), .O_6(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .O_60(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_60), .O_61(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_61), .O_62(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_62), .O_63(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_63), .O_64(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_64), .O_65(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_65), .O_66(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_66), .O_67(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_67), .O_68(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_68), .O_69(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_69), .O_7(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .O_70(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_70), .O_71(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_71), .O_72(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_72), .O_73(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_73), .O_74(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_74), .O_75(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_75), .O_76(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_76), .O_77(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_77), .O_78(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_78), .O_79(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_79), .O_8(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .O_80(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_80), .O_81(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_81), .O_82(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_82), .O_83(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_83), .O_84(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_84), .O_85(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_85), .O_86(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_86), .O_87(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_87), .O_88(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_88), .O_89(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_89), .O_9(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .O_90(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_90), .O_91(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_91), .O_92(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_92), .O_93(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_93), .O_94(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_94), .O_95(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_95), .O_96(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_96), .O_97(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_97), .O_98(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_98), .O_99(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_99), .valid_down(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
assign O_0 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
assign O_1 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1;
assign O_10 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10;
assign O_100 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_100;
assign O_101 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_101;
assign O_102 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_102;
assign O_103 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_103;
assign O_104 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_104;
assign O_105 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_105;
assign O_106 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_106;
assign O_107 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_107;
assign O_108 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_108;
assign O_109 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_109;
assign O_11 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11;
assign O_110 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_110;
assign O_111 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_111;
assign O_112 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_112;
assign O_113 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_113;
assign O_114 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_114;
assign O_115 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_115;
assign O_116 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_116;
assign O_117 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_117;
assign O_118 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_118;
assign O_119 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_119;
assign O_12 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12;
assign O_120 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_120;
assign O_121 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_121;
assign O_122 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_122;
assign O_123 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_123;
assign O_124 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_124;
assign O_125 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_125;
assign O_126 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_126;
assign O_127 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_127;
assign O_128 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_128;
assign O_129 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_129;
assign O_13 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13;
assign O_130 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_130;
assign O_131 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_131;
assign O_132 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_132;
assign O_133 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_133;
assign O_134 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_134;
assign O_135 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_135;
assign O_136 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_136;
assign O_137 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_137;
assign O_138 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_138;
assign O_139 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_139;
assign O_14 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14;
assign O_140 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_140;
assign O_141 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_141;
assign O_142 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_142;
assign O_143 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_143;
assign O_144 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_144;
assign O_145 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_145;
assign O_146 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_146;
assign O_147 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_147;
assign O_148 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_148;
assign O_149 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_149;
assign O_15 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15;
assign O_150 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_150;
assign O_151 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_151;
assign O_152 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_152;
assign O_153 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_153;
assign O_154 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_154;
assign O_155 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_155;
assign O_156 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_156;
assign O_157 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_157;
assign O_158 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_158;
assign O_159 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_159;
assign O_16 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16;
assign O_160 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_160;
assign O_161 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_161;
assign O_162 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_162;
assign O_163 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_163;
assign O_164 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_164;
assign O_165 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_165;
assign O_166 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_166;
assign O_167 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_167;
assign O_168 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_168;
assign O_169 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_169;
assign O_17 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17;
assign O_170 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_170;
assign O_171 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_171;
assign O_172 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_172;
assign O_173 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_173;
assign O_174 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_174;
assign O_175 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_175;
assign O_176 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_176;
assign O_177 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_177;
assign O_178 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_178;
assign O_179 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_179;
assign O_18 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18;
assign O_180 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_180;
assign O_181 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_181;
assign O_182 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_182;
assign O_183 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_183;
assign O_184 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_184;
assign O_185 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_185;
assign O_186 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_186;
assign O_187 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_187;
assign O_188 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_188;
assign O_189 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_189;
assign O_19 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19;
assign O_190 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_190;
assign O_191 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_191;
assign O_192 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_192;
assign O_193 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_193;
assign O_194 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_194;
assign O_195 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_195;
assign O_196 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_196;
assign O_197 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_197;
assign O_198 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_198;
assign O_199 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_199;
assign O_2 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2;
assign O_20 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20;
assign O_21 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21;
assign O_22 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22;
assign O_23 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23;
assign O_24 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24;
assign O_25 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25;
assign O_26 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26;
assign O_27 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27;
assign O_28 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28;
assign O_29 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29;
assign O_3 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3;
assign O_30 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30;
assign O_31 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31;
assign O_32 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32;
assign O_33 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33;
assign O_34 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34;
assign O_35 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35;
assign O_36 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36;
assign O_37 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37;
assign O_38 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38;
assign O_39 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39;
assign O_4 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4;
assign O_40 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_40;
assign O_41 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_41;
assign O_42 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_42;
assign O_43 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_43;
assign O_44 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_44;
assign O_45 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_45;
assign O_46 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_46;
assign O_47 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_47;
assign O_48 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_48;
assign O_49 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_49;
assign O_5 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5;
assign O_50 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_50;
assign O_51 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_51;
assign O_52 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_52;
assign O_53 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_53;
assign O_54 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_54;
assign O_55 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_55;
assign O_56 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_56;
assign O_57 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_57;
assign O_58 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_58;
assign O_59 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_59;
assign O_6 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6;
assign O_60 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_60;
assign O_61 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_61;
assign O_62 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_62;
assign O_63 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_63;
assign O_64 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_64;
assign O_65 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_65;
assign O_66 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_66;
assign O_67 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_67;
assign O_68 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_68;
assign O_69 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_69;
assign O_7 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7;
assign O_70 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_70;
assign O_71 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_71;
assign O_72 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_72;
assign O_73 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_73;
assign O_74 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_74;
assign O_75 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_75;
assign O_76 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_76;
assign O_77 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_77;
assign O_78 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_78;
assign O_79 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_79;
assign O_8 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8;
assign O_80 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_80;
assign O_81 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_81;
assign O_82 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_82;
assign O_83 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_83;
assign O_84 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_84;
assign O_85 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_85;
assign O_86 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_86;
assign O_87 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_87;
assign O_88 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_88;
assign O_89 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_89;
assign O_9 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9;
assign O_90 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_90;
assign O_91 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_91;
assign O_92 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_92;
assign O_93 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_93;
assign O_94 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_94;
assign O_95 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_95;
assign O_96 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_96;
assign O_97 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_97;
assign O_98 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_98;
assign O_99 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_99;
assign valid_down = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
endmodule

