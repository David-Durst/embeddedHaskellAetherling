// Latency = 4
module top(
  input CLK/*verilator public*/, 
  input [7:0] I_0_0_0/*verilator public*/, 
  output [7:0] O_0_0_0/*verilator public*/, 
  input [7:0] I_1_0_0/*verilator public*/, 
  output [7:0] O_1_0_0/*verilator public*/, 
  input [7:0] I_2_0_0/*verilator public*/, 
  output [7:0] O_2_0_0/*verilator public*/, 
  input [7:0] I_3_0_0/*verilator public*/, 
  output [7:0] O_3_0_0/*verilator public*/, 
  output valid_down/*verilator public*/, 
  input valid_up/*verilator public*/
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(CLK), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x373_TREADY(dontcare), // @[:@1298.4]
    .io_in_x373_TDATA({I_0_0_0,I_1_0_0,I_2_0_0,I_3_0_0}), // @[:@1298.4]
    .io_in_x373_TID(8'h0),
    .io_in_x373_TDEST(8'h0),
    .io_in_x374_TVALID(valid_down), // @[:@1298.4]
    .io_in_x374_TDATA({O_0_0_0,O_1_0_0,O_2_0_0,O_3_0_0}), // @[:@1298.4]
    .io_in_x374_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x381_ctrchain cchain ( // @[:@2879.2]
    .clock(CLK), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset, // @[:@6.4]
  input         io_wPort_0_en_0 // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 173:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_68; // @[MemPrimitives.scala 177:32:@23.4]
  wire [31:0] _T_69; // @[MemPrimitives.scala 177:12:@24.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 177:32:@23.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : _T_68; // @[MemPrimitives.scala 177:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 178:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@57.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@104.4]
  wire  _T_57; // @[Counter.scala 285:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@118.4]
  FF bases_0 ( // @[Counter.scala 253:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh16); // @[Counter.scala 285:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh16); // @[Counter.scala 325:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@99.4]
  assign bases_0_io_wPort_0_en_0 = 1'h1; // @[Counter.scala 276:29:@100.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 256:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_133 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = io_rst | done_0_io_output; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = synchronize | io_rst; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = done_0_io_output & _T_166; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module x701_outr_UnitPipe_sm( // @[:@2389.2]
  input   clock, // @[:@2390.4]
  input   reset, // @[:@2391.4]
  input   io_enable, // @[:@2392.4]
  output  io_done, // @[:@2392.4]
  input   io_parentAck, // @[:@2392.4]
  input   io_doneIn_0, // @[:@2392.4]
  output  io_enableOut_0, // @[:@2392.4]
  output  io_childAck_0, // @[:@2392.4]
  input   io_ctrCopyDone_0 // @[:@2392.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@2395.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@2395.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@2398.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@2398.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@2415.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@2415.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@2446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@2460.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@2478.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@2515.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@2532.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@2532.4]
  wire  _T_105; // @[Controllers.scala 165:35:@2430.4]
  wire  _T_107; // @[Controllers.scala 165:60:@2431.4]
  wire  _T_108; // @[Controllers.scala 165:58:@2432.4]
  wire  _T_110; // @[Controllers.scala 165:76:@2433.4]
  wire  _T_111; // @[Controllers.scala 165:74:@2434.4]
  wire  _T_115; // @[Controllers.scala 165:109:@2437.4]
  wire  _T_118; // @[Controllers.scala 165:141:@2439.4]
  wire  _T_126; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  wire  _T_130; // @[Controllers.scala 167:54:@2454.4]
  wire  _T_131; // @[Controllers.scala 167:52:@2455.4]
  wire  _T_138; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  wire  _T_156; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  wire  _T_160; // @[Controllers.scala 169:67:@2486.4]
  wire  _T_161; // @[Controllers.scala 169:86:@2487.4]
  wire  _T_174; // @[Controllers.scala 213:68:@2501.4]
  wire  _T_176; // @[Controllers.scala 213:90:@2503.4]
  wire  _T_178; // @[Controllers.scala 213:132:@2505.4]
  reg  _T_186; // @[package.scala 48:56:@2511.4]
  reg [31:0] _RAND_0;
  wire  _T_187; // @[package.scala 100:41:@2513.4]
  reg  _T_200; // @[package.scala 48:56:@2529.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@2395.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@2398.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@2415.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@2446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@2460.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@2478.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@2515.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@2532.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_105 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@2430.4]
  assign _T_107 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@2431.4]
  assign _T_108 = _T_105 & _T_107; // @[Controllers.scala 165:58:@2432.4]
  assign _T_110 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@2433.4]
  assign _T_111 = _T_108 & _T_110; // @[Controllers.scala 165:74:@2434.4]
  assign _T_115 = _T_111 & io_enable; // @[Controllers.scala 165:109:@2437.4]
  assign _T_118 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@2439.4]
  assign _T_126 = RetimeWrapper_io_out; // @[package.scala 96:25:@2451.4 package.scala 96:25:@2452.4]
  assign _T_130 = _T_126 == 1'h0; // @[Controllers.scala 167:54:@2454.4]
  assign _T_131 = io_doneIn_0 | _T_130; // @[Controllers.scala 167:52:@2455.4]
  assign _T_138 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@2465.4 package.scala 96:25:@2466.4]
  assign _T_156 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@2483.4 package.scala 96:25:@2484.4]
  assign _T_160 = _T_156 == 1'h0; // @[Controllers.scala 169:67:@2486.4]
  assign _T_161 = _T_160 & io_enable; // @[Controllers.scala 169:86:@2487.4]
  assign _T_174 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@2501.4]
  assign _T_176 = _T_174 & _T_105; // @[Controllers.scala 213:90:@2503.4]
  assign _T_178 = ~ done_0_io_output; // @[Controllers.scala 213:132:@2505.4]
  assign _T_187 = done_0_io_output & _T_186; // @[package.scala 100:41:@2513.4]
  assign io_done = RetimeWrapper_4_io_out; // @[Controllers.scala 245:13:@2539.4]
  assign io_enableOut_0 = _T_176 & _T_178; // @[Controllers.scala 213:55:@2509.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@2500.4]
  assign active_0_clock = clock; // @[:@2396.4]
  assign active_0_reset = reset; // @[:@2397.4]
  assign active_0_io_input_set = _T_115 & _T_118; // @[Controllers.scala 165:32:@2441.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@2445.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@2403.4]
  assign done_0_clock = clock; // @[:@2399.4]
  assign done_0_reset = reset; // @[:@2400.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_161; // @[Controllers.scala 169:30:@2491.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@2413.4 Controllers.scala 170:32:@2498.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@2404.4]
  assign iterDone_0_clock = clock; // @[:@2416.4]
  assign iterDone_0_reset = reset; // @[:@2417.4]
  assign iterDone_0_io_input_set = _T_131 & io_enable; // @[Controllers.scala 167:34:@2459.4]
  assign iterDone_0_io_input_reset = _T_138 | io_parentAck; // @[Controllers.scala 92:37:@2427.4 Controllers.scala 168:36:@2475.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@2418.4]
  assign RetimeWrapper_clock = clock; // @[:@2447.4]
  assign RetimeWrapper_reset = reset; // @[:@2448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@2450.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@2449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@2461.4]
  assign RetimeWrapper_1_reset = reset; // @[:@2462.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@2464.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@2463.4]
  assign RetimeWrapper_2_clock = clock; // @[:@2479.4]
  assign RetimeWrapper_2_reset = reset; // @[:@2480.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@2482.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@2481.4]
  assign RetimeWrapper_3_clock = clock; // @[:@2516.4]
  assign RetimeWrapper_3_reset = reset; // @[:@2517.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@2519.4]
  assign RetimeWrapper_3_io_in = _T_187 | io_parentAck; // @[package.scala 94:16:@2518.4]
  assign RetimeWrapper_4_clock = clock; // @[:@2533.4]
  assign RetimeWrapper_4_reset = reset; // @[:@2534.4]
  assign RetimeWrapper_4_io_flow = io_enable; // @[package.scala 95:18:@2536.4]
  assign RetimeWrapper_4_io_in = done_0_io_output & _T_200; // @[package.scala 94:16:@2535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_186 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_200 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_186 <= 1'h0;
    end else begin
      _T_186 <= _T_110;
    end
    if (reset) begin
      _T_200 <= 1'h0;
    end else begin
      _T_200 <= _T_110;
    end
  end
endmodule
module SingleCounter_1( // @[:@2659.2]
  input         clock, // @[:@2660.4]
  input         reset, // @[:@2661.4]
  input         io_input_reset, // @[:@2662.4]
  input         io_input_enable, // @[:@2662.4]
  output [31:0] io_output_count_0, // @[:@2662.4]
  output        io_output_oobs_0, // @[:@2662.4]
  output        io_output_done, // @[:@2662.4]
  output        io_output_saturated // @[:@2662.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2675.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2675.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2675.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2691.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2691.4]
  wire  _T_36; // @[Counter.scala 256:45:@2694.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2719.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2720.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2721.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2722.4]
  wire  _T_57; // @[Counter.scala 285:18:@2724.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2732.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2735.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2736.4]
  wire  _T_75; // @[Counter.scala 314:102:@2740.4]
  wire  _T_77; // @[Counter.scala 314:130:@2741.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2675.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2691.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2694.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2719.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2720.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 283:33:@2721.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2722.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2724.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2732.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2735.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 291:74:@2736.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2740.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2741.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2739.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2743.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2745.4]
  assign io_output_saturated = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 332:25:@2748.4]
  assign bases_0_clock = clock; // @[:@2676.4]
  assign bases_0_reset = reset; // @[:@2677.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2738.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2717.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2718.4]
  assign SRFF_clock = clock; // @[:@2692.4]
  assign SRFF_reset = reset; // @[:@2693.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2696.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2698.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2699.4]
endmodule
module SingleCounter_2( // @[:@2788.2]
  input         clock, // @[:@2789.4]
  input         reset, // @[:@2790.4]
  input         io_setup_saturate, // @[:@2791.4]
  input         io_input_reset, // @[:@2791.4]
  input         io_input_enable, // @[:@2791.4]
  output [31:0] io_output_count_0, // @[:@2791.4]
  output        io_output_oobs_0, // @[:@2791.4]
  output        io_output_done // @[:@2791.4]
);
  wire  bases_0_clock; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 253:53:@2804.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 253:53:@2804.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 253:53:@2804.4]
  wire  SRFF_clock; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_set; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 255:22:@2820.4]
  wire  SRFF_io_output; // @[Counter.scala 255:22:@2820.4]
  wire  _T_36; // @[Counter.scala 256:45:@2823.4]
  wire [31:0] _T_48; // @[Counter.scala 279:52:@2848.4]
  wire [32:0] _T_50; // @[Counter.scala 283:33:@2849.4]
  wire [31:0] _T_51; // @[Counter.scala 283:33:@2850.4]
  wire [31:0] _T_52; // @[Counter.scala 283:33:@2851.4]
  wire  _T_57; // @[Counter.scala 285:18:@2853.4]
  wire [31:0] _T_68; // @[Counter.scala 291:115:@2861.4]
  wire [31:0] _T_70; // @[Counter.scala 291:85:@2863.4]
  wire [31:0] _T_71; // @[Counter.scala 291:152:@2864.4]
  wire [31:0] _T_72; // @[Counter.scala 291:74:@2865.4]
  wire  _T_75; // @[Counter.scala 314:102:@2869.4]
  wire  _T_77; // @[Counter.scala 314:130:@2870.4]
  FF bases_0 ( // @[Counter.scala 253:53:@2804.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 255:22:@2820.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 256:45:@2823.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 279:52:@2848.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2849.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh4); // @[Counter.scala 283:33:@2850.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 283:33:@2851.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh4); // @[Counter.scala 285:18:@2853.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 291:115:@2861.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 32'h0; // @[Counter.scala 291:85:@2863.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 291:152:@2864.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 291:74:@2865.4]
  assign _T_75 = $signed(_T_48) < $signed(32'sh0); // @[Counter.scala 314:102:@2869.4]
  assign _T_77 = $signed(_T_48) >= $signed(32'sh4); // @[Counter.scala 314:130:@2870.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 296:28:@2868.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 314:60:@2872.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 325:20:@2874.4]
  assign bases_0_clock = clock; // @[:@2805.4]
  assign bases_0_reset = reset; // @[:@2806.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 291:31:@2867.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 273:27:@2846.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 276:29:@2847.4]
  assign SRFF_clock = clock; // @[:@2821.4]
  assign SRFF_reset = reset; // @[:@2822.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 256:23:@2825.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 257:25:@2827.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 258:30:@2828.4]
endmodule
module x381_ctrchain( // @[:@2879.2]
  input         clock, // @[:@2880.4]
  input         reset, // @[:@2881.4]
  input         io_input_reset, // @[:@2882.4]
  input         io_input_enable, // @[:@2882.4]
  output [31:0] io_output_counts_1, // @[:@2882.4]
  output [31:0] io_output_counts_0, // @[:@2882.4]
  output        io_output_oobs_0, // @[:@2882.4]
  output        io_output_oobs_1, // @[:@2882.4]
  output        io_output_done // @[:@2882.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 505:46:@2884.4]
  wire [31:0] ctrs_0_io_output_count_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 505:46:@2884.4]
  wire  ctrs_1_clock; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 505:46:@2887.4]
  wire [31:0] ctrs_1_io_output_count_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 505:46:@2887.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 505:46:@2887.4]
  wire  isDone; // @[Counter.scala 533:51:@2904.4]
  reg  wasDone; // @[Counter.scala 534:24:@2905.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 538:69:@2913.4]
  wire  _T_66; // @[Counter.scala 538:80:@2914.4]
  reg  doneLatch; // @[Counter.scala 542:26:@2919.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 543:48:@2920.4]
  wire  _T_74; // @[Counter.scala 543:19:@2921.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 505:46:@2884.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 505:46:@2887.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 533:51:@2904.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 538:69:@2913.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 538:80:@2914.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 543:48:@2920.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 543:19:@2921.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 549:32:@2926.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 549:32:@2923.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2925.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 550:30:@2928.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 538:18:@2916.4]
  assign ctrs_0_clock = clock; // @[:@2885.4]
  assign ctrs_0_reset = reset; // @[:@2886.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2893.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 518:29:@2900.4]
  assign ctrs_1_clock = clock; // @[:@2888.4]
  assign ctrs_1_reset = reset; // @[:@2889.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 524:31:@2903.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 512:24:@2897.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 516:33:@2898.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_12( // @[:@2968.2]
  input   clock, // @[:@2969.4]
  input   reset, // @[:@2970.4]
  input   io_flow, // @[:@2971.4]
  input   io_in, // @[:@2971.4]
  output  io_out // @[:@2971.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@2973.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(41)) sr ( // @[RetimeShiftRegister.scala 15:20:@2973.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@2986.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@2985.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@2984.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@2983.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@2982.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@2980.4]
endmodule
module RetimeWrapper_16( // @[:@3096.2]
  input   clock, // @[:@3097.4]
  input   reset, // @[:@3098.4]
  input   io_flow, // @[:@3099.4]
  input   io_in, // @[:@3099.4]
  output  io_out // @[:@3099.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3101.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@3101.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3114.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3113.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3112.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3111.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3110.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3108.4]
endmodule
module x700_inr_Foreach_SAMPLER_BOX_sm( // @[:@3116.2]
  input   clock, // @[:@3117.4]
  input   reset, // @[:@3118.4]
  input   io_enable, // @[:@3119.4]
  output  io_done, // @[:@3119.4]
  output  io_doneLatch, // @[:@3119.4]
  input   io_ctrDone, // @[:@3119.4]
  output  io_datapathEn, // @[:@3119.4]
  output  io_ctrInc, // @[:@3119.4]
  output  io_ctrRst, // @[:@3119.4]
  input   io_parentAck, // @[:@3119.4]
  input   io_backpressure, // @[:@3119.4]
  input   io_break // @[:@3119.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3121.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3121.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3121.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3124.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3124.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3124.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3180.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3192.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3200.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3216.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3216.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3129.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3130.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3131.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3132.4]
  wire  _T_100; // @[package.scala 100:49:@3149.4]
  reg  _T_103; // @[package.scala 48:56:@3150.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  wire  _T_110; // @[package.scala 100:49:@3165.4]
  reg  _T_113; // @[package.scala 48:56:@3166.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3168.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3173.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3174.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3177.4]
  wire  _T_124; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  wire  _T_126; // @[package.scala 100:49:@3187.4]
  reg  _T_129; // @[package.scala 48:56:@3188.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3210.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3212.4]
  reg  _T_153; // @[package.scala 48:56:@3213.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3223.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3224.4]
  SRFF active ( // @[Controllers.scala 261:22:@3121.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3124.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_12 RetimeWrapper ( // @[package.scala 93:22:@3158.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_12 RetimeWrapper_1 ( // @[package.scala 93:22:@3180.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3192.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3200.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_16 RetimeWrapper_4 ( // @[package.scala 93:22:@3216.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3129.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3130.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3131.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3132.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3149.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3163.4 package.scala 96:25:@3164.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3165.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3168.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3173.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3174.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3177.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3185.4 package.scala 96:25:@3186.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3187.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3212.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3221.4 package.scala 96:25:@3222.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3223.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3224.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3191.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3226.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3176.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3179.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3171.4]
  assign active_clock = clock; // @[:@3122.4]
  assign active_reset = reset; // @[:@3123.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3134.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3138.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3139.4]
  assign done_clock = clock; // @[:@3125.4]
  assign done_reset = reset; // @[:@3126.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3154.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3147.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3148.4]
  assign RetimeWrapper_clock = clock; // @[:@3159.4]
  assign RetimeWrapper_reset = reset; // @[:@3160.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3162.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3161.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3181.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3182.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3184.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3183.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3193.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3194.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3196.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3195.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3201.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3202.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3204.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3203.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3217.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3218.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3220.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3332.2]
  input  [31:0] io_a, // @[:@3335.4]
  output [31:0] io_b // @[:@3335.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3345.4]
endmodule
module _( // @[:@3347.2]
  input  [31:0] io_b, // @[:@3350.4]
  output [31:0] io_result // @[:@3350.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3355.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3355.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3355.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3368.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3363.4]
endmodule
module RetimeWrapper_21( // @[:@3452.2]
  input        clock, // @[:@3453.4]
  input        reset, // @[:@3454.4]
  input        io_flow, // @[:@3455.4]
  input  [7:0] io_in, // @[:@3455.4]
  output [7:0] io_out // @[:@3455.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3457.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3457.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3470.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3469.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@3468.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3467.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3466.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3464.4]
endmodule
module Mem1D_4( // @[:@3472.2]
  input        clock, // @[:@3473.4]
  input        reset, // @[:@3474.4]
  input        io_r_ofs_0, // @[:@3475.4]
  input        io_r_backpressure, // @[:@3475.4]
  input        io_w_ofs_0, // @[:@3475.4]
  input  [7:0] io_w_data_0, // @[:@3475.4]
  input        io_w_en_0, // @[:@3475.4]
  output [7:0] io_output // @[:@3475.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3485.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3494.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@3494.4]
  wire [7:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@3494.4]
  reg [7:0] _T_127; // @[MemPrimitives.scala 560:26:@3479.4]
  reg [31:0] _RAND_0;
  wire  _T_130; // @[MemPrimitives.scala 561:61:@3481.4]
  wire  _T_131; // @[MemPrimitives.scala 561:44:@3482.4]
  wire [7:0] _T_132; // @[MemPrimitives.scala 561:19:@3483.4]
  wire  _T_135; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  wire  _T_137; // @[Mux.scala 46:19:@3492.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@3485.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3494.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_130 = io_w_ofs_0 == 1'h0; // @[MemPrimitives.scala 561:61:@3481.4]
  assign _T_131 = io_w_en_0 & _T_130; // @[MemPrimitives.scala 561:44:@3482.4]
  assign _T_132 = _T_131 ? io_w_data_0 : _T_127; // @[MemPrimitives.scala 561:19:@3483.4]
  assign _T_135 = RetimeWrapper_io_out; // @[package.scala 96:25:@3490.4 package.scala 96:25:@3491.4]
  assign _T_137 = 1'h0 == _T_135; // @[Mux.scala 46:19:@3492.4]
  assign io_output = RetimeWrapper_1_io_out; // @[MemPrimitives.scala 565:17:@3501.4]
  assign RetimeWrapper_clock = clock; // @[:@3486.4]
  assign RetimeWrapper_reset = reset; // @[:@3487.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@3489.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@3488.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3495.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3496.4]
  assign RetimeWrapper_1_io_flow = io_r_backpressure; // @[package.scala 95:18:@3498.4]
  assign RetimeWrapper_1_io_in = _T_137 ? _T_127 : 8'h0; // @[package.scala 94:16:@3497.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_127 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_127 <= 8'h0;
    end else begin
      if (_T_131) begin
        _T_127 <= io_w_data_0;
      end
    end
  end
endmodule
module StickySelects( // @[:@4928.2]
  input   clock, // @[:@4929.4]
  input   reset, // @[:@4930.4]
  input   io_ins_0, // @[:@4931.4]
  input   io_ins_1, // @[:@4931.4]
  input   io_ins_2, // @[:@4931.4]
  output  io_outs_0, // @[:@4931.4]
  output  io_outs_1, // @[:@4931.4]
  output  io_outs_2 // @[:@4931.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4933.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4934.4]
  wire  _T_22; // @[StickySelects.scala 24:52:@4935.4]
  wire  _T_23; // @[StickySelects.scala 24:21:@4936.4]
  reg  _T_26; // @[StickySelects.scala 21:22:@4938.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[StickySelects.scala 22:54:@4939.4]
  wire  _T_29; // @[StickySelects.scala 24:52:@4940.4]
  wire  _T_30; // @[StickySelects.scala 24:21:@4941.4]
  reg  _T_33; // @[StickySelects.scala 21:22:@4943.4]
  reg [31:0] _RAND_2;
  wire  _T_34; // @[StickySelects.scala 22:54:@4944.4]
  wire  _T_36; // @[StickySelects.scala 24:52:@4945.4]
  wire  _T_37; // @[StickySelects.scala 24:21:@4946.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4934.4]
  assign _T_22 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4935.4]
  assign _T_23 = _T_20 ? 1'h0 : _T_22; // @[StickySelects.scala 24:21:@4936.4]
  assign _T_27 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4939.4]
  assign _T_29 = io_ins_1 | _T_26; // @[StickySelects.scala 24:52:@4940.4]
  assign _T_30 = _T_27 ? 1'h0 : _T_29; // @[StickySelects.scala 24:21:@4941.4]
  assign _T_34 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4944.4]
  assign _T_36 = io_ins_2 | _T_33; // @[StickySelects.scala 24:52:@4945.4]
  assign _T_37 = _T_34 ? 1'h0 : _T_36; // @[StickySelects.scala 24:21:@4946.4]
  assign io_outs_0 = _T_20 ? 1'h0 : _T_22; // @[StickySelects.scala 28:52:@4948.4]
  assign io_outs_1 = _T_27 ? 1'h0 : _T_29; // @[StickySelects.scala 28:52:@4949.4]
  assign io_outs_2 = _T_34 ? 1'h0 : _T_36; // @[StickySelects.scala 28:52:@4950.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_33 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_20) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_22;
      end
    end
    if (reset) begin
      _T_26 <= 1'h0;
    end else begin
      if (_T_27) begin
        _T_26 <= 1'h0;
      end else begin
        _T_26 <= _T_29;
      end
    end
    if (reset) begin
      _T_33 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_33 <= 1'h0;
      end else begin
        _T_33 <= _T_36;
      end
    end
  end
endmodule
module StickySelects_2( // @[:@4976.2]
  input   clock, // @[:@4977.4]
  input   reset, // @[:@4978.4]
  input   io_ins_0, // @[:@4979.4]
  input   io_ins_1, // @[:@4979.4]
  input   io_ins_2, // @[:@4979.4]
  input   io_ins_3, // @[:@4979.4]
  input   io_ins_4, // @[:@4979.4]
  input   io_ins_5, // @[:@4979.4]
  output  io_outs_0, // @[:@4979.4]
  output  io_outs_1, // @[:@4979.4]
  output  io_outs_2, // @[:@4979.4]
  output  io_outs_3, // @[:@4979.4]
  output  io_outs_4, // @[:@4979.4]
  output  io_outs_5 // @[:@4979.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@4981.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@4982.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@4983.4]
  wire  _T_22; // @[StickySelects.scala 22:54:@4984.4]
  wire  _T_23; // @[StickySelects.scala 22:54:@4985.4]
  wire  _T_25; // @[StickySelects.scala 24:52:@4986.4]
  wire  _T_26; // @[StickySelects.scala 24:21:@4987.4]
  reg  _T_29; // @[StickySelects.scala 21:22:@4989.4]
  reg [31:0] _RAND_1;
  wire  _T_30; // @[StickySelects.scala 22:54:@4990.4]
  wire  _T_31; // @[StickySelects.scala 22:54:@4991.4]
  wire  _T_32; // @[StickySelects.scala 22:54:@4992.4]
  wire  _T_33; // @[StickySelects.scala 22:54:@4993.4]
  wire  _T_35; // @[StickySelects.scala 24:52:@4994.4]
  wire  _T_36; // @[StickySelects.scala 24:21:@4995.4]
  reg  _T_39; // @[StickySelects.scala 21:22:@4997.4]
  reg [31:0] _RAND_2;
  wire  _T_40; // @[StickySelects.scala 22:54:@4998.4]
  wire  _T_41; // @[StickySelects.scala 22:54:@4999.4]
  wire  _T_42; // @[StickySelects.scala 22:54:@5000.4]
  wire  _T_43; // @[StickySelects.scala 22:54:@5001.4]
  wire  _T_45; // @[StickySelects.scala 24:52:@5002.4]
  wire  _T_46; // @[StickySelects.scala 24:21:@5003.4]
  reg  _T_49; // @[StickySelects.scala 21:22:@5005.4]
  reg [31:0] _RAND_3;
  wire  _T_51; // @[StickySelects.scala 22:54:@5007.4]
  wire  _T_52; // @[StickySelects.scala 22:54:@5008.4]
  wire  _T_53; // @[StickySelects.scala 22:54:@5009.4]
  wire  _T_55; // @[StickySelects.scala 24:52:@5010.4]
  wire  _T_56; // @[StickySelects.scala 24:21:@5011.4]
  reg  _T_59; // @[StickySelects.scala 21:22:@5013.4]
  reg [31:0] _RAND_4;
  wire  _T_62; // @[StickySelects.scala 22:54:@5016.4]
  wire  _T_63; // @[StickySelects.scala 22:54:@5017.4]
  wire  _T_65; // @[StickySelects.scala 24:52:@5018.4]
  wire  _T_66; // @[StickySelects.scala 24:21:@5019.4]
  reg  _T_69; // @[StickySelects.scala 21:22:@5021.4]
  reg [31:0] _RAND_5;
  wire  _T_73; // @[StickySelects.scala 22:54:@5025.4]
  wire  _T_75; // @[StickySelects.scala 24:52:@5026.4]
  wire  _T_76; // @[StickySelects.scala 24:21:@5027.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@4982.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@4983.4]
  assign _T_22 = _T_21 | io_ins_4; // @[StickySelects.scala 22:54:@4984.4]
  assign _T_23 = _T_22 | io_ins_5; // @[StickySelects.scala 22:54:@4985.4]
  assign _T_25 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@4986.4]
  assign _T_26 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 24:21:@4987.4]
  assign _T_30 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@4990.4]
  assign _T_31 = _T_30 | io_ins_3; // @[StickySelects.scala 22:54:@4991.4]
  assign _T_32 = _T_31 | io_ins_4; // @[StickySelects.scala 22:54:@4992.4]
  assign _T_33 = _T_32 | io_ins_5; // @[StickySelects.scala 22:54:@4993.4]
  assign _T_35 = io_ins_1 | _T_29; // @[StickySelects.scala 24:52:@4994.4]
  assign _T_36 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 24:21:@4995.4]
  assign _T_40 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@4998.4]
  assign _T_41 = _T_40 | io_ins_3; // @[StickySelects.scala 22:54:@4999.4]
  assign _T_42 = _T_41 | io_ins_4; // @[StickySelects.scala 22:54:@5000.4]
  assign _T_43 = _T_42 | io_ins_5; // @[StickySelects.scala 22:54:@5001.4]
  assign _T_45 = io_ins_2 | _T_39; // @[StickySelects.scala 24:52:@5002.4]
  assign _T_46 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 24:21:@5003.4]
  assign _T_51 = _T_40 | io_ins_2; // @[StickySelects.scala 22:54:@5007.4]
  assign _T_52 = _T_51 | io_ins_4; // @[StickySelects.scala 22:54:@5008.4]
  assign _T_53 = _T_52 | io_ins_5; // @[StickySelects.scala 22:54:@5009.4]
  assign _T_55 = io_ins_3 | _T_49; // @[StickySelects.scala 24:52:@5010.4]
  assign _T_56 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 24:21:@5011.4]
  assign _T_62 = _T_51 | io_ins_3; // @[StickySelects.scala 22:54:@5016.4]
  assign _T_63 = _T_62 | io_ins_5; // @[StickySelects.scala 22:54:@5017.4]
  assign _T_65 = io_ins_4 | _T_59; // @[StickySelects.scala 24:52:@5018.4]
  assign _T_66 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 24:21:@5019.4]
  assign _T_73 = _T_62 | io_ins_4; // @[StickySelects.scala 22:54:@5025.4]
  assign _T_75 = io_ins_5 | _T_69; // @[StickySelects.scala 24:52:@5026.4]
  assign _T_76 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 24:21:@5027.4]
  assign io_outs_0 = _T_23 ? 1'h0 : _T_25; // @[StickySelects.scala 28:52:@5029.4]
  assign io_outs_1 = _T_33 ? 1'h0 : _T_35; // @[StickySelects.scala 28:52:@5030.4]
  assign io_outs_2 = _T_43 ? 1'h0 : _T_45; // @[StickySelects.scala 28:52:@5031.4]
  assign io_outs_3 = _T_53 ? 1'h0 : _T_55; // @[StickySelects.scala 28:52:@5032.4]
  assign io_outs_4 = _T_63 ? 1'h0 : _T_65; // @[StickySelects.scala 28:52:@5033.4]
  assign io_outs_5 = _T_73 ? 1'h0 : _T_75; // @[StickySelects.scala 28:52:@5034.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_29 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_39 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_49 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_59 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_69 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_23) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_25;
      end
    end
    if (reset) begin
      _T_29 <= 1'h0;
    end else begin
      if (_T_33) begin
        _T_29 <= 1'h0;
      end else begin
        _T_29 <= _T_35;
      end
    end
    if (reset) begin
      _T_39 <= 1'h0;
    end else begin
      if (_T_43) begin
        _T_39 <= 1'h0;
      end else begin
        _T_39 <= _T_45;
      end
    end
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      if (_T_53) begin
        _T_49 <= 1'h0;
      end else begin
        _T_49 <= _T_55;
      end
    end
    if (reset) begin
      _T_59 <= 1'h0;
    end else begin
      if (_T_63) begin
        _T_59 <= 1'h0;
      end else begin
        _T_59 <= _T_65;
      end
    end
    if (reset) begin
      _T_69 <= 1'h0;
    end else begin
      if (_T_73) begin
        _T_69 <= 1'h0;
      end else begin
        _T_69 <= _T_75;
      end
    end
  end
endmodule
module RetimeWrapper_52( // @[:@5612.2]
  input   clock, // @[:@5613.4]
  input   reset, // @[:@5614.4]
  input   io_flow, // @[:@5615.4]
  input   io_in, // @[:@5615.4]
  output  io_out // @[:@5615.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@5617.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@5617.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@5630.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@5629.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@5628.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@5627.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@5626.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@5624.4]
endmodule
module x386_lb_0( // @[:@7904.2]
  input        clock, // @[:@7905.4]
  input        reset, // @[:@7906.4]
  input  [2:0] io_rPort_17_banks_0, // @[:@7907.4]
  input        io_rPort_17_ofs_0, // @[:@7907.4]
  input        io_rPort_17_en_0, // @[:@7907.4]
  input        io_rPort_17_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_17_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_16_banks_0, // @[:@7907.4]
  input        io_rPort_16_ofs_0, // @[:@7907.4]
  input        io_rPort_16_en_0, // @[:@7907.4]
  input        io_rPort_16_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_16_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_15_banks_0, // @[:@7907.4]
  input        io_rPort_15_ofs_0, // @[:@7907.4]
  input        io_rPort_15_en_0, // @[:@7907.4]
  input        io_rPort_15_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_15_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_14_banks_0, // @[:@7907.4]
  input        io_rPort_14_ofs_0, // @[:@7907.4]
  input        io_rPort_14_en_0, // @[:@7907.4]
  input        io_rPort_14_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_14_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_13_banks_0, // @[:@7907.4]
  input        io_rPort_13_ofs_0, // @[:@7907.4]
  input        io_rPort_13_en_0, // @[:@7907.4]
  input        io_rPort_13_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_13_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_12_banks_0, // @[:@7907.4]
  input        io_rPort_12_ofs_0, // @[:@7907.4]
  input        io_rPort_12_en_0, // @[:@7907.4]
  input        io_rPort_12_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_12_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@7907.4]
  input        io_rPort_11_ofs_0, // @[:@7907.4]
  input        io_rPort_11_en_0, // @[:@7907.4]
  input        io_rPort_11_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_11_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@7907.4]
  input        io_rPort_10_ofs_0, // @[:@7907.4]
  input        io_rPort_10_en_0, // @[:@7907.4]
  input        io_rPort_10_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_10_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@7907.4]
  input        io_rPort_9_ofs_0, // @[:@7907.4]
  input        io_rPort_9_en_0, // @[:@7907.4]
  input        io_rPort_9_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_9_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@7907.4]
  input        io_rPort_8_ofs_0, // @[:@7907.4]
  input        io_rPort_8_en_0, // @[:@7907.4]
  input        io_rPort_8_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_8_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@7907.4]
  input        io_rPort_7_ofs_0, // @[:@7907.4]
  input        io_rPort_7_en_0, // @[:@7907.4]
  input        io_rPort_7_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_7_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@7907.4]
  input        io_rPort_6_ofs_0, // @[:@7907.4]
  input        io_rPort_6_en_0, // @[:@7907.4]
  input        io_rPort_6_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_6_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@7907.4]
  input        io_rPort_5_ofs_0, // @[:@7907.4]
  input        io_rPort_5_en_0, // @[:@7907.4]
  input        io_rPort_5_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_5_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@7907.4]
  input        io_rPort_4_ofs_0, // @[:@7907.4]
  input        io_rPort_4_en_0, // @[:@7907.4]
  input        io_rPort_4_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_4_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@7907.4]
  input        io_rPort_3_ofs_0, // @[:@7907.4]
  input        io_rPort_3_en_0, // @[:@7907.4]
  input        io_rPort_3_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_3_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@7907.4]
  input        io_rPort_2_ofs_0, // @[:@7907.4]
  input        io_rPort_2_en_0, // @[:@7907.4]
  input        io_rPort_2_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_2_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@7907.4]
  input        io_rPort_1_ofs_0, // @[:@7907.4]
  input        io_rPort_1_en_0, // @[:@7907.4]
  input        io_rPort_1_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_1_output_0, // @[:@7907.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@7907.4]
  input        io_rPort_0_ofs_0, // @[:@7907.4]
  input        io_rPort_0_en_0, // @[:@7907.4]
  input        io_rPort_0_backpressure, // @[:@7907.4]
  output [7:0] io_rPort_0_output_0, // @[:@7907.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@7907.4]
  input        io_wPort_3_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_3_data_0, // @[:@7907.4]
  input        io_wPort_3_en_0, // @[:@7907.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@7907.4]
  input        io_wPort_2_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_2_data_0, // @[:@7907.4]
  input        io_wPort_2_en_0, // @[:@7907.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@7907.4]
  input        io_wPort_1_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_1_data_0, // @[:@7907.4]
  input        io_wPort_1_en_0, // @[:@7907.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@7907.4]
  input        io_wPort_0_ofs_0, // @[:@7907.4]
  input  [7:0] io_wPort_0_data_0, // @[:@7907.4]
  input        io_wPort_0_en_0 // @[:@7907.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@8050.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@8050.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@8066.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@8066.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@8082.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@8082.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@8098.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@8098.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@8114.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@8114.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@8130.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@8130.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@8146.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@8146.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@8162.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@8162.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@8178.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@8178.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@8194.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@8194.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@8210.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@8210.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@8226.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@8226.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@8242.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@8242.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@8258.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@8258.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@8274.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@8274.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@8290.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@8290.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@8491.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@8523.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@8564.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@8620.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@8667.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@8699.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@8740.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@8796.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@8843.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@8875.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@8916.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@8972.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@9019.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@9051.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@9092.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@9148.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@9199.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@9207.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@9215.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@9223.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@9247.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@9255.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@9263.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@9271.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@9295.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@9303.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@9311.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@9319.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@9343.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@9351.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@9359.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@9367.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@9391.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@9399.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@9407.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@9415.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@9439.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@9447.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@9455.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@9463.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@9487.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@9495.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@9503.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@9511.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@9535.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@9543.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@9551.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@9559.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@9583.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@9591.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@9599.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@9607.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@9631.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@9639.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@9647.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@9655.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@9679.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@9687.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@9695.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@9703.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@9727.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@9735.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@9743.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@9751.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@9775.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@9783.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@9791.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@9799.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@9823.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@9831.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@9839.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@9847.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@9871.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@9879.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@9887.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@9895.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@9919.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@9927.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@9935.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@9943.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@9967.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@9975.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@9983.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@9991.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@10015.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@10023.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@10031.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@10039.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@10039.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@8306.4]
  wire  _T_703; // @[MemPrimitives.scala 83:102:@8308.4]
  wire [9:0] _T_705; // @[Cat.scala 30:58:@8310.4]
  wire  _T_710; // @[MemPrimitives.scala 82:210:@8317.4]
  wire  _T_713; // @[MemPrimitives.scala 83:102:@8319.4]
  wire [9:0] _T_715; // @[Cat.scala 30:58:@8321.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@8328.4]
  wire  _T_723; // @[MemPrimitives.scala 83:102:@8330.4]
  wire [9:0] _T_725; // @[Cat.scala 30:58:@8332.4]
  wire  _T_730; // @[MemPrimitives.scala 82:210:@8339.4]
  wire  _T_733; // @[MemPrimitives.scala 83:102:@8341.4]
  wire [9:0] _T_735; // @[Cat.scala 30:58:@8343.4]
  wire  _T_740; // @[MemPrimitives.scala 82:210:@8350.4]
  wire  _T_743; // @[MemPrimitives.scala 83:102:@8352.4]
  wire [9:0] _T_745; // @[Cat.scala 30:58:@8354.4]
  wire  _T_750; // @[MemPrimitives.scala 82:210:@8361.4]
  wire  _T_753; // @[MemPrimitives.scala 83:102:@8363.4]
  wire [9:0] _T_755; // @[Cat.scala 30:58:@8365.4]
  wire  _T_760; // @[MemPrimitives.scala 82:210:@8372.4]
  wire  _T_763; // @[MemPrimitives.scala 83:102:@8374.4]
  wire [9:0] _T_765; // @[Cat.scala 30:58:@8376.4]
  wire  _T_770; // @[MemPrimitives.scala 82:210:@8383.4]
  wire  _T_773; // @[MemPrimitives.scala 83:102:@8385.4]
  wire [9:0] _T_775; // @[Cat.scala 30:58:@8387.4]
  wire  _T_780; // @[MemPrimitives.scala 82:210:@8394.4]
  wire  _T_783; // @[MemPrimitives.scala 83:102:@8396.4]
  wire [9:0] _T_785; // @[Cat.scala 30:58:@8398.4]
  wire  _T_790; // @[MemPrimitives.scala 82:210:@8405.4]
  wire  _T_793; // @[MemPrimitives.scala 83:102:@8407.4]
  wire [9:0] _T_795; // @[Cat.scala 30:58:@8409.4]
  wire  _T_800; // @[MemPrimitives.scala 82:210:@8416.4]
  wire  _T_803; // @[MemPrimitives.scala 83:102:@8418.4]
  wire [9:0] _T_805; // @[Cat.scala 30:58:@8420.4]
  wire  _T_810; // @[MemPrimitives.scala 82:210:@8427.4]
  wire  _T_813; // @[MemPrimitives.scala 83:102:@8429.4]
  wire [9:0] _T_815; // @[Cat.scala 30:58:@8431.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@8438.4]
  wire  _T_823; // @[MemPrimitives.scala 83:102:@8440.4]
  wire [9:0] _T_825; // @[Cat.scala 30:58:@8442.4]
  wire  _T_830; // @[MemPrimitives.scala 82:210:@8449.4]
  wire  _T_833; // @[MemPrimitives.scala 83:102:@8451.4]
  wire [9:0] _T_835; // @[Cat.scala 30:58:@8453.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@8460.4]
  wire  _T_843; // @[MemPrimitives.scala 83:102:@8462.4]
  wire [9:0] _T_845; // @[Cat.scala 30:58:@8464.4]
  wire  _T_850; // @[MemPrimitives.scala 82:210:@8471.4]
  wire  _T_853; // @[MemPrimitives.scala 83:102:@8473.4]
  wire [9:0] _T_855; // @[Cat.scala 30:58:@8475.4]
  wire  _T_860; // @[MemPrimitives.scala 110:210:@8482.4]
  wire  _T_865; // @[MemPrimitives.scala 110:210:@8485.4]
  wire  _T_870; // @[MemPrimitives.scala 110:210:@8488.4]
  wire  _T_874; // @[MemPrimitives.scala 123:41:@8497.4]
  wire  _T_875; // @[MemPrimitives.scala 123:41:@8498.4]
  wire  _T_876; // @[MemPrimitives.scala 123:41:@8499.4]
  wire [2:0] _T_878; // @[Cat.scala 30:58:@8501.4]
  wire [2:0] _T_880; // @[Cat.scala 30:58:@8503.4]
  wire [2:0] _T_882; // @[Cat.scala 30:58:@8505.4]
  wire [2:0] _T_883; // @[Mux.scala 31:69:@8506.4]
  wire [2:0] _T_884; // @[Mux.scala 31:69:@8507.4]
  wire  _T_889; // @[MemPrimitives.scala 110:210:@8514.4]
  wire  _T_894; // @[MemPrimitives.scala 110:210:@8517.4]
  wire  _T_899; // @[MemPrimitives.scala 110:210:@8520.4]
  wire  _T_903; // @[MemPrimitives.scala 123:41:@8529.4]
  wire  _T_904; // @[MemPrimitives.scala 123:41:@8530.4]
  wire  _T_905; // @[MemPrimitives.scala 123:41:@8531.4]
  wire [2:0] _T_907; // @[Cat.scala 30:58:@8533.4]
  wire [2:0] _T_909; // @[Cat.scala 30:58:@8535.4]
  wire [2:0] _T_911; // @[Cat.scala 30:58:@8537.4]
  wire [2:0] _T_912; // @[Mux.scala 31:69:@8538.4]
  wire [2:0] _T_913; // @[Mux.scala 31:69:@8539.4]
  wire  _T_918; // @[MemPrimitives.scala 110:210:@8546.4]
  wire  _T_923; // @[MemPrimitives.scala 110:210:@8549.4]
  wire  _T_928; // @[MemPrimitives.scala 110:210:@8552.4]
  wire  _T_933; // @[MemPrimitives.scala 110:210:@8555.4]
  wire  _T_938; // @[MemPrimitives.scala 110:210:@8558.4]
  wire  _T_943; // @[MemPrimitives.scala 110:210:@8561.4]
  wire  _T_947; // @[MemPrimitives.scala 123:41:@8573.4]
  wire  _T_948; // @[MemPrimitives.scala 123:41:@8574.4]
  wire  _T_949; // @[MemPrimitives.scala 123:41:@8575.4]
  wire  _T_950; // @[MemPrimitives.scala 123:41:@8576.4]
  wire  _T_951; // @[MemPrimitives.scala 123:41:@8577.4]
  wire  _T_952; // @[MemPrimitives.scala 123:41:@8578.4]
  wire [2:0] _T_954; // @[Cat.scala 30:58:@8580.4]
  wire [2:0] _T_956; // @[Cat.scala 30:58:@8582.4]
  wire [2:0] _T_958; // @[Cat.scala 30:58:@8584.4]
  wire [2:0] _T_960; // @[Cat.scala 30:58:@8586.4]
  wire [2:0] _T_962; // @[Cat.scala 30:58:@8588.4]
  wire [2:0] _T_964; // @[Cat.scala 30:58:@8590.4]
  wire [2:0] _T_965; // @[Mux.scala 31:69:@8591.4]
  wire [2:0] _T_966; // @[Mux.scala 31:69:@8592.4]
  wire [2:0] _T_967; // @[Mux.scala 31:69:@8593.4]
  wire [2:0] _T_968; // @[Mux.scala 31:69:@8594.4]
  wire [2:0] _T_969; // @[Mux.scala 31:69:@8595.4]
  wire  _T_974; // @[MemPrimitives.scala 110:210:@8602.4]
  wire  _T_979; // @[MemPrimitives.scala 110:210:@8605.4]
  wire  _T_984; // @[MemPrimitives.scala 110:210:@8608.4]
  wire  _T_989; // @[MemPrimitives.scala 110:210:@8611.4]
  wire  _T_994; // @[MemPrimitives.scala 110:210:@8614.4]
  wire  _T_999; // @[MemPrimitives.scala 110:210:@8617.4]
  wire  _T_1003; // @[MemPrimitives.scala 123:41:@8629.4]
  wire  _T_1004; // @[MemPrimitives.scala 123:41:@8630.4]
  wire  _T_1005; // @[MemPrimitives.scala 123:41:@8631.4]
  wire  _T_1006; // @[MemPrimitives.scala 123:41:@8632.4]
  wire  _T_1007; // @[MemPrimitives.scala 123:41:@8633.4]
  wire  _T_1008; // @[MemPrimitives.scala 123:41:@8634.4]
  wire [2:0] _T_1010; // @[Cat.scala 30:58:@8636.4]
  wire [2:0] _T_1012; // @[Cat.scala 30:58:@8638.4]
  wire [2:0] _T_1014; // @[Cat.scala 30:58:@8640.4]
  wire [2:0] _T_1016; // @[Cat.scala 30:58:@8642.4]
  wire [2:0] _T_1018; // @[Cat.scala 30:58:@8644.4]
  wire [2:0] _T_1020; // @[Cat.scala 30:58:@8646.4]
  wire [2:0] _T_1021; // @[Mux.scala 31:69:@8647.4]
  wire [2:0] _T_1022; // @[Mux.scala 31:69:@8648.4]
  wire [2:0] _T_1023; // @[Mux.scala 31:69:@8649.4]
  wire [2:0] _T_1024; // @[Mux.scala 31:69:@8650.4]
  wire [2:0] _T_1025; // @[Mux.scala 31:69:@8651.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@8658.4]
  wire  _T_1035; // @[MemPrimitives.scala 110:210:@8661.4]
  wire  _T_1040; // @[MemPrimitives.scala 110:210:@8664.4]
  wire  _T_1044; // @[MemPrimitives.scala 123:41:@8673.4]
  wire  _T_1045; // @[MemPrimitives.scala 123:41:@8674.4]
  wire  _T_1046; // @[MemPrimitives.scala 123:41:@8675.4]
  wire [2:0] _T_1048; // @[Cat.scala 30:58:@8677.4]
  wire [2:0] _T_1050; // @[Cat.scala 30:58:@8679.4]
  wire [2:0] _T_1052; // @[Cat.scala 30:58:@8681.4]
  wire [2:0] _T_1053; // @[Mux.scala 31:69:@8682.4]
  wire [2:0] _T_1054; // @[Mux.scala 31:69:@8683.4]
  wire  _T_1059; // @[MemPrimitives.scala 110:210:@8690.4]
  wire  _T_1064; // @[MemPrimitives.scala 110:210:@8693.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:210:@8696.4]
  wire  _T_1073; // @[MemPrimitives.scala 123:41:@8705.4]
  wire  _T_1074; // @[MemPrimitives.scala 123:41:@8706.4]
  wire  _T_1075; // @[MemPrimitives.scala 123:41:@8707.4]
  wire [2:0] _T_1077; // @[Cat.scala 30:58:@8709.4]
  wire [2:0] _T_1079; // @[Cat.scala 30:58:@8711.4]
  wire [2:0] _T_1081; // @[Cat.scala 30:58:@8713.4]
  wire [2:0] _T_1082; // @[Mux.scala 31:69:@8714.4]
  wire [2:0] _T_1083; // @[Mux.scala 31:69:@8715.4]
  wire  _T_1088; // @[MemPrimitives.scala 110:210:@8722.4]
  wire  _T_1093; // @[MemPrimitives.scala 110:210:@8725.4]
  wire  _T_1098; // @[MemPrimitives.scala 110:210:@8728.4]
  wire  _T_1103; // @[MemPrimitives.scala 110:210:@8731.4]
  wire  _T_1108; // @[MemPrimitives.scala 110:210:@8734.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:210:@8737.4]
  wire  _T_1117; // @[MemPrimitives.scala 123:41:@8749.4]
  wire  _T_1118; // @[MemPrimitives.scala 123:41:@8750.4]
  wire  _T_1119; // @[MemPrimitives.scala 123:41:@8751.4]
  wire  _T_1120; // @[MemPrimitives.scala 123:41:@8752.4]
  wire  _T_1121; // @[MemPrimitives.scala 123:41:@8753.4]
  wire  _T_1122; // @[MemPrimitives.scala 123:41:@8754.4]
  wire [2:0] _T_1124; // @[Cat.scala 30:58:@8756.4]
  wire [2:0] _T_1126; // @[Cat.scala 30:58:@8758.4]
  wire [2:0] _T_1128; // @[Cat.scala 30:58:@8760.4]
  wire [2:0] _T_1130; // @[Cat.scala 30:58:@8762.4]
  wire [2:0] _T_1132; // @[Cat.scala 30:58:@8764.4]
  wire [2:0] _T_1134; // @[Cat.scala 30:58:@8766.4]
  wire [2:0] _T_1135; // @[Mux.scala 31:69:@8767.4]
  wire [2:0] _T_1136; // @[Mux.scala 31:69:@8768.4]
  wire [2:0] _T_1137; // @[Mux.scala 31:69:@8769.4]
  wire [2:0] _T_1138; // @[Mux.scala 31:69:@8770.4]
  wire [2:0] _T_1139; // @[Mux.scala 31:69:@8771.4]
  wire  _T_1144; // @[MemPrimitives.scala 110:210:@8778.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:210:@8781.4]
  wire  _T_1154; // @[MemPrimitives.scala 110:210:@8784.4]
  wire  _T_1159; // @[MemPrimitives.scala 110:210:@8787.4]
  wire  _T_1164; // @[MemPrimitives.scala 110:210:@8790.4]
  wire  _T_1169; // @[MemPrimitives.scala 110:210:@8793.4]
  wire  _T_1173; // @[MemPrimitives.scala 123:41:@8805.4]
  wire  _T_1174; // @[MemPrimitives.scala 123:41:@8806.4]
  wire  _T_1175; // @[MemPrimitives.scala 123:41:@8807.4]
  wire  _T_1176; // @[MemPrimitives.scala 123:41:@8808.4]
  wire  _T_1177; // @[MemPrimitives.scala 123:41:@8809.4]
  wire  _T_1178; // @[MemPrimitives.scala 123:41:@8810.4]
  wire [2:0] _T_1180; // @[Cat.scala 30:58:@8812.4]
  wire [2:0] _T_1182; // @[Cat.scala 30:58:@8814.4]
  wire [2:0] _T_1184; // @[Cat.scala 30:58:@8816.4]
  wire [2:0] _T_1186; // @[Cat.scala 30:58:@8818.4]
  wire [2:0] _T_1188; // @[Cat.scala 30:58:@8820.4]
  wire [2:0] _T_1190; // @[Cat.scala 30:58:@8822.4]
  wire [2:0] _T_1191; // @[Mux.scala 31:69:@8823.4]
  wire [2:0] _T_1192; // @[Mux.scala 31:69:@8824.4]
  wire [2:0] _T_1193; // @[Mux.scala 31:69:@8825.4]
  wire [2:0] _T_1194; // @[Mux.scala 31:69:@8826.4]
  wire [2:0] _T_1195; // @[Mux.scala 31:69:@8827.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@8834.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:210:@8837.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@8840.4]
  wire  _T_1214; // @[MemPrimitives.scala 123:41:@8849.4]
  wire  _T_1215; // @[MemPrimitives.scala 123:41:@8850.4]
  wire  _T_1216; // @[MemPrimitives.scala 123:41:@8851.4]
  wire [2:0] _T_1218; // @[Cat.scala 30:58:@8853.4]
  wire [2:0] _T_1220; // @[Cat.scala 30:58:@8855.4]
  wire [2:0] _T_1222; // @[Cat.scala 30:58:@8857.4]
  wire [2:0] _T_1223; // @[Mux.scala 31:69:@8858.4]
  wire [2:0] _T_1224; // @[Mux.scala 31:69:@8859.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:210:@8866.4]
  wire  _T_1234; // @[MemPrimitives.scala 110:210:@8869.4]
  wire  _T_1239; // @[MemPrimitives.scala 110:210:@8872.4]
  wire  _T_1243; // @[MemPrimitives.scala 123:41:@8881.4]
  wire  _T_1244; // @[MemPrimitives.scala 123:41:@8882.4]
  wire  _T_1245; // @[MemPrimitives.scala 123:41:@8883.4]
  wire [2:0] _T_1247; // @[Cat.scala 30:58:@8885.4]
  wire [2:0] _T_1249; // @[Cat.scala 30:58:@8887.4]
  wire [2:0] _T_1251; // @[Cat.scala 30:58:@8889.4]
  wire [2:0] _T_1252; // @[Mux.scala 31:69:@8890.4]
  wire [2:0] _T_1253; // @[Mux.scala 31:69:@8891.4]
  wire  _T_1258; // @[MemPrimitives.scala 110:210:@8898.4]
  wire  _T_1263; // @[MemPrimitives.scala 110:210:@8901.4]
  wire  _T_1268; // @[MemPrimitives.scala 110:210:@8904.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:210:@8907.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@8910.4]
  wire  _T_1283; // @[MemPrimitives.scala 110:210:@8913.4]
  wire  _T_1287; // @[MemPrimitives.scala 123:41:@8925.4]
  wire  _T_1288; // @[MemPrimitives.scala 123:41:@8926.4]
  wire  _T_1289; // @[MemPrimitives.scala 123:41:@8927.4]
  wire  _T_1290; // @[MemPrimitives.scala 123:41:@8928.4]
  wire  _T_1291; // @[MemPrimitives.scala 123:41:@8929.4]
  wire  _T_1292; // @[MemPrimitives.scala 123:41:@8930.4]
  wire [2:0] _T_1294; // @[Cat.scala 30:58:@8932.4]
  wire [2:0] _T_1296; // @[Cat.scala 30:58:@8934.4]
  wire [2:0] _T_1298; // @[Cat.scala 30:58:@8936.4]
  wire [2:0] _T_1300; // @[Cat.scala 30:58:@8938.4]
  wire [2:0] _T_1302; // @[Cat.scala 30:58:@8940.4]
  wire [2:0] _T_1304; // @[Cat.scala 30:58:@8942.4]
  wire [2:0] _T_1305; // @[Mux.scala 31:69:@8943.4]
  wire [2:0] _T_1306; // @[Mux.scala 31:69:@8944.4]
  wire [2:0] _T_1307; // @[Mux.scala 31:69:@8945.4]
  wire [2:0] _T_1308; // @[Mux.scala 31:69:@8946.4]
  wire [2:0] _T_1309; // @[Mux.scala 31:69:@8947.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@8954.4]
  wire  _T_1319; // @[MemPrimitives.scala 110:210:@8957.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@8960.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:210:@8963.4]
  wire  _T_1334; // @[MemPrimitives.scala 110:210:@8966.4]
  wire  _T_1339; // @[MemPrimitives.scala 110:210:@8969.4]
  wire  _T_1343; // @[MemPrimitives.scala 123:41:@8981.4]
  wire  _T_1344; // @[MemPrimitives.scala 123:41:@8982.4]
  wire  _T_1345; // @[MemPrimitives.scala 123:41:@8983.4]
  wire  _T_1346; // @[MemPrimitives.scala 123:41:@8984.4]
  wire  _T_1347; // @[MemPrimitives.scala 123:41:@8985.4]
  wire  _T_1348; // @[MemPrimitives.scala 123:41:@8986.4]
  wire [2:0] _T_1350; // @[Cat.scala 30:58:@8988.4]
  wire [2:0] _T_1352; // @[Cat.scala 30:58:@8990.4]
  wire [2:0] _T_1354; // @[Cat.scala 30:58:@8992.4]
  wire [2:0] _T_1356; // @[Cat.scala 30:58:@8994.4]
  wire [2:0] _T_1358; // @[Cat.scala 30:58:@8996.4]
  wire [2:0] _T_1360; // @[Cat.scala 30:58:@8998.4]
  wire [2:0] _T_1361; // @[Mux.scala 31:69:@8999.4]
  wire [2:0] _T_1362; // @[Mux.scala 31:69:@9000.4]
  wire [2:0] _T_1363; // @[Mux.scala 31:69:@9001.4]
  wire [2:0] _T_1364; // @[Mux.scala 31:69:@9002.4]
  wire [2:0] _T_1365; // @[Mux.scala 31:69:@9003.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@9010.4]
  wire  _T_1375; // @[MemPrimitives.scala 110:210:@9013.4]
  wire  _T_1380; // @[MemPrimitives.scala 110:210:@9016.4]
  wire  _T_1384; // @[MemPrimitives.scala 123:41:@9025.4]
  wire  _T_1385; // @[MemPrimitives.scala 123:41:@9026.4]
  wire  _T_1386; // @[MemPrimitives.scala 123:41:@9027.4]
  wire [2:0] _T_1388; // @[Cat.scala 30:58:@9029.4]
  wire [2:0] _T_1390; // @[Cat.scala 30:58:@9031.4]
  wire [2:0] _T_1392; // @[Cat.scala 30:58:@9033.4]
  wire [2:0] _T_1393; // @[Mux.scala 31:69:@9034.4]
  wire [2:0] _T_1394; // @[Mux.scala 31:69:@9035.4]
  wire  _T_1399; // @[MemPrimitives.scala 110:210:@9042.4]
  wire  _T_1404; // @[MemPrimitives.scala 110:210:@9045.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:210:@9048.4]
  wire  _T_1413; // @[MemPrimitives.scala 123:41:@9057.4]
  wire  _T_1414; // @[MemPrimitives.scala 123:41:@9058.4]
  wire  _T_1415; // @[MemPrimitives.scala 123:41:@9059.4]
  wire [2:0] _T_1417; // @[Cat.scala 30:58:@9061.4]
  wire [2:0] _T_1419; // @[Cat.scala 30:58:@9063.4]
  wire [2:0] _T_1421; // @[Cat.scala 30:58:@9065.4]
  wire [2:0] _T_1422; // @[Mux.scala 31:69:@9066.4]
  wire [2:0] _T_1423; // @[Mux.scala 31:69:@9067.4]
  wire  _T_1428; // @[MemPrimitives.scala 110:210:@9074.4]
  wire  _T_1433; // @[MemPrimitives.scala 110:210:@9077.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@9080.4]
  wire  _T_1443; // @[MemPrimitives.scala 110:210:@9083.4]
  wire  _T_1448; // @[MemPrimitives.scala 110:210:@9086.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:210:@9089.4]
  wire  _T_1457; // @[MemPrimitives.scala 123:41:@9101.4]
  wire  _T_1458; // @[MemPrimitives.scala 123:41:@9102.4]
  wire  _T_1459; // @[MemPrimitives.scala 123:41:@9103.4]
  wire  _T_1460; // @[MemPrimitives.scala 123:41:@9104.4]
  wire  _T_1461; // @[MemPrimitives.scala 123:41:@9105.4]
  wire  _T_1462; // @[MemPrimitives.scala 123:41:@9106.4]
  wire [2:0] _T_1464; // @[Cat.scala 30:58:@9108.4]
  wire [2:0] _T_1466; // @[Cat.scala 30:58:@9110.4]
  wire [2:0] _T_1468; // @[Cat.scala 30:58:@9112.4]
  wire [2:0] _T_1470; // @[Cat.scala 30:58:@9114.4]
  wire [2:0] _T_1472; // @[Cat.scala 30:58:@9116.4]
  wire [2:0] _T_1474; // @[Cat.scala 30:58:@9118.4]
  wire [2:0] _T_1475; // @[Mux.scala 31:69:@9119.4]
  wire [2:0] _T_1476; // @[Mux.scala 31:69:@9120.4]
  wire [2:0] _T_1477; // @[Mux.scala 31:69:@9121.4]
  wire [2:0] _T_1478; // @[Mux.scala 31:69:@9122.4]
  wire [2:0] _T_1479; // @[Mux.scala 31:69:@9123.4]
  wire  _T_1484; // @[MemPrimitives.scala 110:210:@9130.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:210:@9133.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@9136.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:210:@9139.4]
  wire  _T_1504; // @[MemPrimitives.scala 110:210:@9142.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:210:@9145.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@9157.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@9158.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@9159.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@9160.4]
  wire  _T_1517; // @[MemPrimitives.scala 123:41:@9161.4]
  wire  _T_1518; // @[MemPrimitives.scala 123:41:@9162.4]
  wire [2:0] _T_1520; // @[Cat.scala 30:58:@9164.4]
  wire [2:0] _T_1522; // @[Cat.scala 30:58:@9166.4]
  wire [2:0] _T_1524; // @[Cat.scala 30:58:@9168.4]
  wire [2:0] _T_1526; // @[Cat.scala 30:58:@9170.4]
  wire [2:0] _T_1528; // @[Cat.scala 30:58:@9172.4]
  wire [2:0] _T_1530; // @[Cat.scala 30:58:@9174.4]
  wire [2:0] _T_1531; // @[Mux.scala 31:69:@9175.4]
  wire [2:0] _T_1532; // @[Mux.scala 31:69:@9176.4]
  wire [2:0] _T_1533; // @[Mux.scala 31:69:@9177.4]
  wire [2:0] _T_1534; // @[Mux.scala 31:69:@9178.4]
  wire [2:0] _T_1535; // @[Mux.scala 31:69:@9179.4]
  wire  _T_1567; // @[package.scala 96:25:@9220.4 package.scala 96:25:@9221.4]
  wire [7:0] _T_1571; // @[Mux.scala 31:69:@9230.4]
  wire  _T_1564; // @[package.scala 96:25:@9212.4 package.scala 96:25:@9213.4]
  wire [7:0] _T_1572; // @[Mux.scala 31:69:@9231.4]
  wire  _T_1561; // @[package.scala 96:25:@9204.4 package.scala 96:25:@9205.4]
  wire  _T_1602; // @[package.scala 96:25:@9268.4 package.scala 96:25:@9269.4]
  wire [7:0] _T_1606; // @[Mux.scala 31:69:@9278.4]
  wire  _T_1599; // @[package.scala 96:25:@9260.4 package.scala 96:25:@9261.4]
  wire [7:0] _T_1607; // @[Mux.scala 31:69:@9279.4]
  wire  _T_1596; // @[package.scala 96:25:@9252.4 package.scala 96:25:@9253.4]
  wire  _T_1637; // @[package.scala 96:25:@9316.4 package.scala 96:25:@9317.4]
  wire [7:0] _T_1641; // @[Mux.scala 31:69:@9326.4]
  wire  _T_1634; // @[package.scala 96:25:@9308.4 package.scala 96:25:@9309.4]
  wire [7:0] _T_1642; // @[Mux.scala 31:69:@9327.4]
  wire  _T_1631; // @[package.scala 96:25:@9300.4 package.scala 96:25:@9301.4]
  wire  _T_1672; // @[package.scala 96:25:@9364.4 package.scala 96:25:@9365.4]
  wire [7:0] _T_1676; // @[Mux.scala 31:69:@9374.4]
  wire  _T_1669; // @[package.scala 96:25:@9356.4 package.scala 96:25:@9357.4]
  wire [7:0] _T_1677; // @[Mux.scala 31:69:@9375.4]
  wire  _T_1666; // @[package.scala 96:25:@9348.4 package.scala 96:25:@9349.4]
  wire  _T_1707; // @[package.scala 96:25:@9412.4 package.scala 96:25:@9413.4]
  wire [7:0] _T_1711; // @[Mux.scala 31:69:@9422.4]
  wire  _T_1704; // @[package.scala 96:25:@9404.4 package.scala 96:25:@9405.4]
  wire [7:0] _T_1712; // @[Mux.scala 31:69:@9423.4]
  wire  _T_1701; // @[package.scala 96:25:@9396.4 package.scala 96:25:@9397.4]
  wire  _T_1742; // @[package.scala 96:25:@9460.4 package.scala 96:25:@9461.4]
  wire [7:0] _T_1746; // @[Mux.scala 31:69:@9470.4]
  wire  _T_1739; // @[package.scala 96:25:@9452.4 package.scala 96:25:@9453.4]
  wire [7:0] _T_1747; // @[Mux.scala 31:69:@9471.4]
  wire  _T_1736; // @[package.scala 96:25:@9444.4 package.scala 96:25:@9445.4]
  wire  _T_1777; // @[package.scala 96:25:@9508.4 package.scala 96:25:@9509.4]
  wire [7:0] _T_1781; // @[Mux.scala 31:69:@9518.4]
  wire  _T_1774; // @[package.scala 96:25:@9500.4 package.scala 96:25:@9501.4]
  wire [7:0] _T_1782; // @[Mux.scala 31:69:@9519.4]
  wire  _T_1771; // @[package.scala 96:25:@9492.4 package.scala 96:25:@9493.4]
  wire  _T_1812; // @[package.scala 96:25:@9556.4 package.scala 96:25:@9557.4]
  wire [7:0] _T_1816; // @[Mux.scala 31:69:@9566.4]
  wire  _T_1809; // @[package.scala 96:25:@9548.4 package.scala 96:25:@9549.4]
  wire [7:0] _T_1817; // @[Mux.scala 31:69:@9567.4]
  wire  _T_1806; // @[package.scala 96:25:@9540.4 package.scala 96:25:@9541.4]
  wire  _T_1847; // @[package.scala 96:25:@9604.4 package.scala 96:25:@9605.4]
  wire [7:0] _T_1851; // @[Mux.scala 31:69:@9614.4]
  wire  _T_1844; // @[package.scala 96:25:@9596.4 package.scala 96:25:@9597.4]
  wire [7:0] _T_1852; // @[Mux.scala 31:69:@9615.4]
  wire  _T_1841; // @[package.scala 96:25:@9588.4 package.scala 96:25:@9589.4]
  wire  _T_1882; // @[package.scala 96:25:@9652.4 package.scala 96:25:@9653.4]
  wire [7:0] _T_1886; // @[Mux.scala 31:69:@9662.4]
  wire  _T_1879; // @[package.scala 96:25:@9644.4 package.scala 96:25:@9645.4]
  wire [7:0] _T_1887; // @[Mux.scala 31:69:@9663.4]
  wire  _T_1876; // @[package.scala 96:25:@9636.4 package.scala 96:25:@9637.4]
  wire  _T_1917; // @[package.scala 96:25:@9700.4 package.scala 96:25:@9701.4]
  wire [7:0] _T_1921; // @[Mux.scala 31:69:@9710.4]
  wire  _T_1914; // @[package.scala 96:25:@9692.4 package.scala 96:25:@9693.4]
  wire [7:0] _T_1922; // @[Mux.scala 31:69:@9711.4]
  wire  _T_1911; // @[package.scala 96:25:@9684.4 package.scala 96:25:@9685.4]
  wire  _T_1952; // @[package.scala 96:25:@9748.4 package.scala 96:25:@9749.4]
  wire [7:0] _T_1956; // @[Mux.scala 31:69:@9758.4]
  wire  _T_1949; // @[package.scala 96:25:@9740.4 package.scala 96:25:@9741.4]
  wire [7:0] _T_1957; // @[Mux.scala 31:69:@9759.4]
  wire  _T_1946; // @[package.scala 96:25:@9732.4 package.scala 96:25:@9733.4]
  wire  _T_1987; // @[package.scala 96:25:@9796.4 package.scala 96:25:@9797.4]
  wire [7:0] _T_1991; // @[Mux.scala 31:69:@9806.4]
  wire  _T_1984; // @[package.scala 96:25:@9788.4 package.scala 96:25:@9789.4]
  wire [7:0] _T_1992; // @[Mux.scala 31:69:@9807.4]
  wire  _T_1981; // @[package.scala 96:25:@9780.4 package.scala 96:25:@9781.4]
  wire  _T_2022; // @[package.scala 96:25:@9844.4 package.scala 96:25:@9845.4]
  wire [7:0] _T_2026; // @[Mux.scala 31:69:@9854.4]
  wire  _T_2019; // @[package.scala 96:25:@9836.4 package.scala 96:25:@9837.4]
  wire [7:0] _T_2027; // @[Mux.scala 31:69:@9855.4]
  wire  _T_2016; // @[package.scala 96:25:@9828.4 package.scala 96:25:@9829.4]
  wire  _T_2057; // @[package.scala 96:25:@9892.4 package.scala 96:25:@9893.4]
  wire [7:0] _T_2061; // @[Mux.scala 31:69:@9902.4]
  wire  _T_2054; // @[package.scala 96:25:@9884.4 package.scala 96:25:@9885.4]
  wire [7:0] _T_2062; // @[Mux.scala 31:69:@9903.4]
  wire  _T_2051; // @[package.scala 96:25:@9876.4 package.scala 96:25:@9877.4]
  wire  _T_2092; // @[package.scala 96:25:@9940.4 package.scala 96:25:@9941.4]
  wire [7:0] _T_2096; // @[Mux.scala 31:69:@9950.4]
  wire  _T_2089; // @[package.scala 96:25:@9932.4 package.scala 96:25:@9933.4]
  wire [7:0] _T_2097; // @[Mux.scala 31:69:@9951.4]
  wire  _T_2086; // @[package.scala 96:25:@9924.4 package.scala 96:25:@9925.4]
  wire  _T_2127; // @[package.scala 96:25:@9988.4 package.scala 96:25:@9989.4]
  wire [7:0] _T_2131; // @[Mux.scala 31:69:@9998.4]
  wire  _T_2124; // @[package.scala 96:25:@9980.4 package.scala 96:25:@9981.4]
  wire [7:0] _T_2132; // @[Mux.scala 31:69:@9999.4]
  wire  _T_2121; // @[package.scala 96:25:@9972.4 package.scala 96:25:@9973.4]
  wire  _T_2162; // @[package.scala 96:25:@10036.4 package.scala 96:25:@10037.4]
  wire [7:0] _T_2166; // @[Mux.scala 31:69:@10046.4]
  wire  _T_2159; // @[package.scala 96:25:@10028.4 package.scala 96:25:@10029.4]
  wire [7:0] _T_2167; // @[Mux.scala 31:69:@10047.4]
  wire  _T_2156; // @[package.scala 96:25:@10020.4 package.scala 96:25:@10021.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@8050.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@8066.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@8082.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@8098.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@8114.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@8130.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@8146.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@8162.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@8178.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@8194.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@8210.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@8226.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@8242.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@8258.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@8274.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@8290.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@8491.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2)
  );
  StickySelects StickySelects_1 ( // @[MemPrimitives.scala 121:29:@8523.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2)
  );
  StickySelects_2 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@8564.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_2 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@8620.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects StickySelects_4 ( // @[MemPrimitives.scala 121:29:@8667.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2)
  );
  StickySelects StickySelects_5 ( // @[MemPrimitives.scala 121:29:@8699.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2)
  );
  StickySelects_2 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@8740.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_2 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@8796.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects StickySelects_8 ( // @[MemPrimitives.scala 121:29:@8843.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2)
  );
  StickySelects StickySelects_9 ( // @[MemPrimitives.scala 121:29:@8875.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2)
  );
  StickySelects_2 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@8916.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_2 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@8972.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects StickySelects_12 ( // @[MemPrimitives.scala 121:29:@9019.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2)
  );
  StickySelects StickySelects_13 ( // @[MemPrimitives.scala 121:29:@9051.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2)
  );
  StickySelects_2 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@9092.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_2 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@9148.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@9199.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@9207.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@9215.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@9223.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@9247.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@9255.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@9263.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@9271.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@9295.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@9303.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@9311.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@9319.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@9343.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@9351.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@9359.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@9367.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@9391.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@9399.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@9407.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@9415.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@9439.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@9447.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@9455.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@9463.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@9487.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@9495.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@9503.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@9511.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@9535.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@9543.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@9551.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@9559.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@9583.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@9591.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@9599.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@9607.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@9631.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@9639.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@9647.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@9655.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_40 ( // @[package.scala 93:22:@9679.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_41 ( // @[package.scala 93:22:@9687.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_42 ( // @[package.scala 93:22:@9695.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_43 ( // @[package.scala 93:22:@9703.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_44 ( // @[package.scala 93:22:@9727.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_45 ( // @[package.scala 93:22:@9735.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_46 ( // @[package.scala 93:22:@9743.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_47 ( // @[package.scala 93:22:@9751.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_48 ( // @[package.scala 93:22:@9775.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_49 ( // @[package.scala 93:22:@9783.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_50 ( // @[package.scala 93:22:@9791.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_51 ( // @[package.scala 93:22:@9799.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_52 ( // @[package.scala 93:22:@9823.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_53 ( // @[package.scala 93:22:@9831.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_54 ( // @[package.scala 93:22:@9839.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_55 ( // @[package.scala 93:22:@9847.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_56 ( // @[package.scala 93:22:@9871.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_57 ( // @[package.scala 93:22:@9879.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_58 ( // @[package.scala 93:22:@9887.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_59 ( // @[package.scala 93:22:@9895.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_60 ( // @[package.scala 93:22:@9919.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_61 ( // @[package.scala 93:22:@9927.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_62 ( // @[package.scala 93:22:@9935.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_63 ( // @[package.scala 93:22:@9943.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_64 ( // @[package.scala 93:22:@9967.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_65 ( // @[package.scala 93:22:@9975.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_66 ( // @[package.scala 93:22:@9983.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_67 ( // @[package.scala 93:22:@9991.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_68 ( // @[package.scala 93:22:@10015.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_69 ( // @[package.scala 93:22:@10023.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_70 ( // @[package.scala 93:22:@10031.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_71 ( // @[package.scala 93:22:@10039.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8306.4]
  assign _T_703 = io_wPort_0_en_0 & _T_700; // @[MemPrimitives.scala 83:102:@8308.4]
  assign _T_705 = {_T_703,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8310.4]
  assign _T_710 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8317.4]
  assign _T_713 = io_wPort_1_en_0 & _T_710; // @[MemPrimitives.scala 83:102:@8319.4]
  assign _T_715 = {_T_713,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8321.4]
  assign _T_720 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8328.4]
  assign _T_723 = io_wPort_2_en_0 & _T_720; // @[MemPrimitives.scala 83:102:@8330.4]
  assign _T_725 = {_T_723,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8332.4]
  assign _T_730 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@8339.4]
  assign _T_733 = io_wPort_3_en_0 & _T_730; // @[MemPrimitives.scala 83:102:@8341.4]
  assign _T_735 = {_T_733,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8343.4]
  assign _T_740 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8350.4]
  assign _T_743 = io_wPort_0_en_0 & _T_740; // @[MemPrimitives.scala 83:102:@8352.4]
  assign _T_745 = {_T_743,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8354.4]
  assign _T_750 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8361.4]
  assign _T_753 = io_wPort_1_en_0 & _T_750; // @[MemPrimitives.scala 83:102:@8363.4]
  assign _T_755 = {_T_753,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8365.4]
  assign _T_760 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8372.4]
  assign _T_763 = io_wPort_2_en_0 & _T_760; // @[MemPrimitives.scala 83:102:@8374.4]
  assign _T_765 = {_T_763,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8376.4]
  assign _T_770 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@8383.4]
  assign _T_773 = io_wPort_3_en_0 & _T_770; // @[MemPrimitives.scala 83:102:@8385.4]
  assign _T_775 = {_T_773,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8387.4]
  assign _T_780 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8394.4]
  assign _T_783 = io_wPort_0_en_0 & _T_780; // @[MemPrimitives.scala 83:102:@8396.4]
  assign _T_785 = {_T_783,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8398.4]
  assign _T_790 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8405.4]
  assign _T_793 = io_wPort_1_en_0 & _T_790; // @[MemPrimitives.scala 83:102:@8407.4]
  assign _T_795 = {_T_793,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8409.4]
  assign _T_800 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8416.4]
  assign _T_803 = io_wPort_2_en_0 & _T_800; // @[MemPrimitives.scala 83:102:@8418.4]
  assign _T_805 = {_T_803,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8420.4]
  assign _T_810 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@8427.4]
  assign _T_813 = io_wPort_3_en_0 & _T_810; // @[MemPrimitives.scala 83:102:@8429.4]
  assign _T_815 = {_T_813,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8431.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8438.4]
  assign _T_823 = io_wPort_0_en_0 & _T_820; // @[MemPrimitives.scala 83:102:@8440.4]
  assign _T_825 = {_T_823,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@8442.4]
  assign _T_830 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8449.4]
  assign _T_833 = io_wPort_1_en_0 & _T_830; // @[MemPrimitives.scala 83:102:@8451.4]
  assign _T_835 = {_T_833,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@8453.4]
  assign _T_840 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8460.4]
  assign _T_843 = io_wPort_2_en_0 & _T_840; // @[MemPrimitives.scala 83:102:@8462.4]
  assign _T_845 = {_T_843,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@8464.4]
  assign _T_850 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@8471.4]
  assign _T_853 = io_wPort_3_en_0 & _T_850; // @[MemPrimitives.scala 83:102:@8473.4]
  assign _T_855 = {_T_853,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@8475.4]
  assign _T_860 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8482.4]
  assign _T_865 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8485.4]
  assign _T_870 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8488.4]
  assign _T_874 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@8497.4]
  assign _T_875 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@8498.4]
  assign _T_876 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@8499.4]
  assign _T_878 = {_T_874,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@8501.4]
  assign _T_880 = {_T_875,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@8503.4]
  assign _T_882 = {_T_876,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@8505.4]
  assign _T_883 = _T_875 ? _T_880 : _T_882; // @[Mux.scala 31:69:@8506.4]
  assign _T_884 = _T_874 ? _T_878 : _T_883; // @[Mux.scala 31:69:@8507.4]
  assign _T_889 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8514.4]
  assign _T_894 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8517.4]
  assign _T_899 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8520.4]
  assign _T_903 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@8529.4]
  assign _T_904 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@8530.4]
  assign _T_905 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@8531.4]
  assign _T_907 = {_T_903,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@8533.4]
  assign _T_909 = {_T_904,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@8535.4]
  assign _T_911 = {_T_905,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@8537.4]
  assign _T_912 = _T_904 ? _T_909 : _T_911; // @[Mux.scala 31:69:@8538.4]
  assign _T_913 = _T_903 ? _T_907 : _T_912; // @[Mux.scala 31:69:@8539.4]
  assign _T_918 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8546.4]
  assign _T_923 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8549.4]
  assign _T_928 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8552.4]
  assign _T_933 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8555.4]
  assign _T_938 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8558.4]
  assign _T_943 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8561.4]
  assign _T_947 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@8573.4]
  assign _T_948 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@8574.4]
  assign _T_949 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@8575.4]
  assign _T_950 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@8576.4]
  assign _T_951 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@8577.4]
  assign _T_952 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@8578.4]
  assign _T_954 = {_T_947,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@8580.4]
  assign _T_956 = {_T_948,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@8582.4]
  assign _T_958 = {_T_949,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@8584.4]
  assign _T_960 = {_T_950,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@8586.4]
  assign _T_962 = {_T_951,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@8588.4]
  assign _T_964 = {_T_952,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@8590.4]
  assign _T_965 = _T_951 ? _T_962 : _T_964; // @[Mux.scala 31:69:@8591.4]
  assign _T_966 = _T_950 ? _T_960 : _T_965; // @[Mux.scala 31:69:@8592.4]
  assign _T_967 = _T_949 ? _T_958 : _T_966; // @[Mux.scala 31:69:@8593.4]
  assign _T_968 = _T_948 ? _T_956 : _T_967; // @[Mux.scala 31:69:@8594.4]
  assign _T_969 = _T_947 ? _T_954 : _T_968; // @[Mux.scala 31:69:@8595.4]
  assign _T_974 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8602.4]
  assign _T_979 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8605.4]
  assign _T_984 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8608.4]
  assign _T_989 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8611.4]
  assign _T_994 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8614.4]
  assign _T_999 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@8617.4]
  assign _T_1003 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@8629.4]
  assign _T_1004 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@8630.4]
  assign _T_1005 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@8631.4]
  assign _T_1006 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@8632.4]
  assign _T_1007 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@8633.4]
  assign _T_1008 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@8634.4]
  assign _T_1010 = {_T_1003,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@8636.4]
  assign _T_1012 = {_T_1004,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@8638.4]
  assign _T_1014 = {_T_1005,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@8640.4]
  assign _T_1016 = {_T_1006,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@8642.4]
  assign _T_1018 = {_T_1007,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@8644.4]
  assign _T_1020 = {_T_1008,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@8646.4]
  assign _T_1021 = _T_1007 ? _T_1018 : _T_1020; // @[Mux.scala 31:69:@8647.4]
  assign _T_1022 = _T_1006 ? _T_1016 : _T_1021; // @[Mux.scala 31:69:@8648.4]
  assign _T_1023 = _T_1005 ? _T_1014 : _T_1022; // @[Mux.scala 31:69:@8649.4]
  assign _T_1024 = _T_1004 ? _T_1012 : _T_1023; // @[Mux.scala 31:69:@8650.4]
  assign _T_1025 = _T_1003 ? _T_1010 : _T_1024; // @[Mux.scala 31:69:@8651.4]
  assign _T_1030 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8658.4]
  assign _T_1035 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8661.4]
  assign _T_1040 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8664.4]
  assign _T_1044 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@8673.4]
  assign _T_1045 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@8674.4]
  assign _T_1046 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@8675.4]
  assign _T_1048 = {_T_1044,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@8677.4]
  assign _T_1050 = {_T_1045,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@8679.4]
  assign _T_1052 = {_T_1046,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@8681.4]
  assign _T_1053 = _T_1045 ? _T_1050 : _T_1052; // @[Mux.scala 31:69:@8682.4]
  assign _T_1054 = _T_1044 ? _T_1048 : _T_1053; // @[Mux.scala 31:69:@8683.4]
  assign _T_1059 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8690.4]
  assign _T_1064 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8693.4]
  assign _T_1069 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8696.4]
  assign _T_1073 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@8705.4]
  assign _T_1074 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@8706.4]
  assign _T_1075 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@8707.4]
  assign _T_1077 = {_T_1073,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@8709.4]
  assign _T_1079 = {_T_1074,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@8711.4]
  assign _T_1081 = {_T_1075,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@8713.4]
  assign _T_1082 = _T_1074 ? _T_1079 : _T_1081; // @[Mux.scala 31:69:@8714.4]
  assign _T_1083 = _T_1073 ? _T_1077 : _T_1082; // @[Mux.scala 31:69:@8715.4]
  assign _T_1088 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8722.4]
  assign _T_1093 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8725.4]
  assign _T_1098 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8728.4]
  assign _T_1103 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8731.4]
  assign _T_1108 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8734.4]
  assign _T_1113 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8737.4]
  assign _T_1117 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@8749.4]
  assign _T_1118 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@8750.4]
  assign _T_1119 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@8751.4]
  assign _T_1120 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@8752.4]
  assign _T_1121 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@8753.4]
  assign _T_1122 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@8754.4]
  assign _T_1124 = {_T_1117,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@8756.4]
  assign _T_1126 = {_T_1118,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@8758.4]
  assign _T_1128 = {_T_1119,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@8760.4]
  assign _T_1130 = {_T_1120,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@8762.4]
  assign _T_1132 = {_T_1121,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@8764.4]
  assign _T_1134 = {_T_1122,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@8766.4]
  assign _T_1135 = _T_1121 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@8767.4]
  assign _T_1136 = _T_1120 ? _T_1130 : _T_1135; // @[Mux.scala 31:69:@8768.4]
  assign _T_1137 = _T_1119 ? _T_1128 : _T_1136; // @[Mux.scala 31:69:@8769.4]
  assign _T_1138 = _T_1118 ? _T_1126 : _T_1137; // @[Mux.scala 31:69:@8770.4]
  assign _T_1139 = _T_1117 ? _T_1124 : _T_1138; // @[Mux.scala 31:69:@8771.4]
  assign _T_1144 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8778.4]
  assign _T_1149 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8781.4]
  assign _T_1154 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8784.4]
  assign _T_1159 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8787.4]
  assign _T_1164 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8790.4]
  assign _T_1169 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@8793.4]
  assign _T_1173 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@8805.4]
  assign _T_1174 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@8806.4]
  assign _T_1175 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@8807.4]
  assign _T_1176 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@8808.4]
  assign _T_1177 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@8809.4]
  assign _T_1178 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@8810.4]
  assign _T_1180 = {_T_1173,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@8812.4]
  assign _T_1182 = {_T_1174,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@8814.4]
  assign _T_1184 = {_T_1175,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@8816.4]
  assign _T_1186 = {_T_1176,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@8818.4]
  assign _T_1188 = {_T_1177,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@8820.4]
  assign _T_1190 = {_T_1178,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@8822.4]
  assign _T_1191 = _T_1177 ? _T_1188 : _T_1190; // @[Mux.scala 31:69:@8823.4]
  assign _T_1192 = _T_1176 ? _T_1186 : _T_1191; // @[Mux.scala 31:69:@8824.4]
  assign _T_1193 = _T_1175 ? _T_1184 : _T_1192; // @[Mux.scala 31:69:@8825.4]
  assign _T_1194 = _T_1174 ? _T_1182 : _T_1193; // @[Mux.scala 31:69:@8826.4]
  assign _T_1195 = _T_1173 ? _T_1180 : _T_1194; // @[Mux.scala 31:69:@8827.4]
  assign _T_1200 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8834.4]
  assign _T_1205 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8837.4]
  assign _T_1210 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8840.4]
  assign _T_1214 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@8849.4]
  assign _T_1215 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@8850.4]
  assign _T_1216 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@8851.4]
  assign _T_1218 = {_T_1214,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@8853.4]
  assign _T_1220 = {_T_1215,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@8855.4]
  assign _T_1222 = {_T_1216,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@8857.4]
  assign _T_1223 = _T_1215 ? _T_1220 : _T_1222; // @[Mux.scala 31:69:@8858.4]
  assign _T_1224 = _T_1214 ? _T_1218 : _T_1223; // @[Mux.scala 31:69:@8859.4]
  assign _T_1229 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8866.4]
  assign _T_1234 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8869.4]
  assign _T_1239 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8872.4]
  assign _T_1243 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@8881.4]
  assign _T_1244 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@8882.4]
  assign _T_1245 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@8883.4]
  assign _T_1247 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@8885.4]
  assign _T_1249 = {_T_1244,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@8887.4]
  assign _T_1251 = {_T_1245,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@8889.4]
  assign _T_1252 = _T_1244 ? _T_1249 : _T_1251; // @[Mux.scala 31:69:@8890.4]
  assign _T_1253 = _T_1243 ? _T_1247 : _T_1252; // @[Mux.scala 31:69:@8891.4]
  assign _T_1258 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8898.4]
  assign _T_1263 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8901.4]
  assign _T_1268 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8904.4]
  assign _T_1273 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8907.4]
  assign _T_1278 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8910.4]
  assign _T_1283 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8913.4]
  assign _T_1287 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@8925.4]
  assign _T_1288 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@8926.4]
  assign _T_1289 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@8927.4]
  assign _T_1290 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@8928.4]
  assign _T_1291 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@8929.4]
  assign _T_1292 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@8930.4]
  assign _T_1294 = {_T_1287,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@8932.4]
  assign _T_1296 = {_T_1288,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@8934.4]
  assign _T_1298 = {_T_1289,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@8936.4]
  assign _T_1300 = {_T_1290,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@8938.4]
  assign _T_1302 = {_T_1291,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@8940.4]
  assign _T_1304 = {_T_1292,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@8942.4]
  assign _T_1305 = _T_1291 ? _T_1302 : _T_1304; // @[Mux.scala 31:69:@8943.4]
  assign _T_1306 = _T_1290 ? _T_1300 : _T_1305; // @[Mux.scala 31:69:@8944.4]
  assign _T_1307 = _T_1289 ? _T_1298 : _T_1306; // @[Mux.scala 31:69:@8945.4]
  assign _T_1308 = _T_1288 ? _T_1296 : _T_1307; // @[Mux.scala 31:69:@8946.4]
  assign _T_1309 = _T_1287 ? _T_1294 : _T_1308; // @[Mux.scala 31:69:@8947.4]
  assign _T_1314 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8954.4]
  assign _T_1319 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8957.4]
  assign _T_1324 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8960.4]
  assign _T_1329 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8963.4]
  assign _T_1334 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8966.4]
  assign _T_1339 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@8969.4]
  assign _T_1343 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@8981.4]
  assign _T_1344 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@8982.4]
  assign _T_1345 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@8983.4]
  assign _T_1346 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@8984.4]
  assign _T_1347 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@8985.4]
  assign _T_1348 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@8986.4]
  assign _T_1350 = {_T_1343,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@8988.4]
  assign _T_1352 = {_T_1344,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@8990.4]
  assign _T_1354 = {_T_1345,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@8992.4]
  assign _T_1356 = {_T_1346,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@8994.4]
  assign _T_1358 = {_T_1347,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@8996.4]
  assign _T_1360 = {_T_1348,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@8998.4]
  assign _T_1361 = _T_1347 ? _T_1358 : _T_1360; // @[Mux.scala 31:69:@8999.4]
  assign _T_1362 = _T_1346 ? _T_1356 : _T_1361; // @[Mux.scala 31:69:@9000.4]
  assign _T_1363 = _T_1345 ? _T_1354 : _T_1362; // @[Mux.scala 31:69:@9001.4]
  assign _T_1364 = _T_1344 ? _T_1352 : _T_1363; // @[Mux.scala 31:69:@9002.4]
  assign _T_1365 = _T_1343 ? _T_1350 : _T_1364; // @[Mux.scala 31:69:@9003.4]
  assign _T_1370 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9010.4]
  assign _T_1375 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9013.4]
  assign _T_1380 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9016.4]
  assign _T_1384 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@9025.4]
  assign _T_1385 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@9026.4]
  assign _T_1386 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@9027.4]
  assign _T_1388 = {_T_1384,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@9029.4]
  assign _T_1390 = {_T_1385,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@9031.4]
  assign _T_1392 = {_T_1386,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@9033.4]
  assign _T_1393 = _T_1385 ? _T_1390 : _T_1392; // @[Mux.scala 31:69:@9034.4]
  assign _T_1394 = _T_1384 ? _T_1388 : _T_1393; // @[Mux.scala 31:69:@9035.4]
  assign _T_1399 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9042.4]
  assign _T_1404 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9045.4]
  assign _T_1409 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9048.4]
  assign _T_1413 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@9057.4]
  assign _T_1414 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@9058.4]
  assign _T_1415 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@9059.4]
  assign _T_1417 = {_T_1413,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@9061.4]
  assign _T_1419 = {_T_1414,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@9063.4]
  assign _T_1421 = {_T_1415,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@9065.4]
  assign _T_1422 = _T_1414 ? _T_1419 : _T_1421; // @[Mux.scala 31:69:@9066.4]
  assign _T_1423 = _T_1413 ? _T_1417 : _T_1422; // @[Mux.scala 31:69:@9067.4]
  assign _T_1428 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9074.4]
  assign _T_1433 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9077.4]
  assign _T_1438 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9080.4]
  assign _T_1443 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9083.4]
  assign _T_1448 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9086.4]
  assign _T_1453 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9089.4]
  assign _T_1457 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@9101.4]
  assign _T_1458 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@9102.4]
  assign _T_1459 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@9103.4]
  assign _T_1460 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@9104.4]
  assign _T_1461 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@9105.4]
  assign _T_1462 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@9106.4]
  assign _T_1464 = {_T_1457,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@9108.4]
  assign _T_1466 = {_T_1458,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@9110.4]
  assign _T_1468 = {_T_1459,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@9112.4]
  assign _T_1470 = {_T_1460,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@9114.4]
  assign _T_1472 = {_T_1461,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@9116.4]
  assign _T_1474 = {_T_1462,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@9118.4]
  assign _T_1475 = _T_1461 ? _T_1472 : _T_1474; // @[Mux.scala 31:69:@9119.4]
  assign _T_1476 = _T_1460 ? _T_1470 : _T_1475; // @[Mux.scala 31:69:@9120.4]
  assign _T_1477 = _T_1459 ? _T_1468 : _T_1476; // @[Mux.scala 31:69:@9121.4]
  assign _T_1478 = _T_1458 ? _T_1466 : _T_1477; // @[Mux.scala 31:69:@9122.4]
  assign _T_1479 = _T_1457 ? _T_1464 : _T_1478; // @[Mux.scala 31:69:@9123.4]
  assign _T_1484 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9130.4]
  assign _T_1489 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9133.4]
  assign _T_1494 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9136.4]
  assign _T_1499 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9139.4]
  assign _T_1504 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9142.4]
  assign _T_1509 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@9145.4]
  assign _T_1513 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@9157.4]
  assign _T_1514 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@9158.4]
  assign _T_1515 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@9159.4]
  assign _T_1516 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@9160.4]
  assign _T_1517 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@9161.4]
  assign _T_1518 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@9162.4]
  assign _T_1520 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@9164.4]
  assign _T_1522 = {_T_1514,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@9166.4]
  assign _T_1524 = {_T_1515,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@9168.4]
  assign _T_1526 = {_T_1516,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@9170.4]
  assign _T_1528 = {_T_1517,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@9172.4]
  assign _T_1530 = {_T_1518,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@9174.4]
  assign _T_1531 = _T_1517 ? _T_1528 : _T_1530; // @[Mux.scala 31:69:@9175.4]
  assign _T_1532 = _T_1516 ? _T_1526 : _T_1531; // @[Mux.scala 31:69:@9176.4]
  assign _T_1533 = _T_1515 ? _T_1524 : _T_1532; // @[Mux.scala 31:69:@9177.4]
  assign _T_1534 = _T_1514 ? _T_1522 : _T_1533; // @[Mux.scala 31:69:@9178.4]
  assign _T_1535 = _T_1513 ? _T_1520 : _T_1534; // @[Mux.scala 31:69:@9179.4]
  assign _T_1567 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@9220.4 package.scala 96:25:@9221.4]
  assign _T_1571 = _T_1567 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9230.4]
  assign _T_1564 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@9212.4 package.scala 96:25:@9213.4]
  assign _T_1572 = _T_1564 ? Mem1D_7_io_output : _T_1571; // @[Mux.scala 31:69:@9231.4]
  assign _T_1561 = RetimeWrapper_io_out; // @[package.scala 96:25:@9204.4 package.scala 96:25:@9205.4]
  assign _T_1602 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@9268.4 package.scala 96:25:@9269.4]
  assign _T_1606 = _T_1602 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9278.4]
  assign _T_1599 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@9260.4 package.scala 96:25:@9261.4]
  assign _T_1607 = _T_1599 ? Mem1D_6_io_output : _T_1606; // @[Mux.scala 31:69:@9279.4]
  assign _T_1596 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@9252.4 package.scala 96:25:@9253.4]
  assign _T_1637 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@9316.4 package.scala 96:25:@9317.4]
  assign _T_1641 = _T_1637 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9326.4]
  assign _T_1634 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@9308.4 package.scala 96:25:@9309.4]
  assign _T_1642 = _T_1634 ? Mem1D_6_io_output : _T_1641; // @[Mux.scala 31:69:@9327.4]
  assign _T_1631 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@9300.4 package.scala 96:25:@9301.4]
  assign _T_1672 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@9364.4 package.scala 96:25:@9365.4]
  assign _T_1676 = _T_1672 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9374.4]
  assign _T_1669 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@9356.4 package.scala 96:25:@9357.4]
  assign _T_1677 = _T_1669 ? Mem1D_7_io_output : _T_1676; // @[Mux.scala 31:69:@9375.4]
  assign _T_1666 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@9348.4 package.scala 96:25:@9349.4]
  assign _T_1707 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@9412.4 package.scala 96:25:@9413.4]
  assign _T_1711 = _T_1707 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9422.4]
  assign _T_1704 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@9404.4 package.scala 96:25:@9405.4]
  assign _T_1712 = _T_1704 ? Mem1D_7_io_output : _T_1711; // @[Mux.scala 31:69:@9423.4]
  assign _T_1701 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@9396.4 package.scala 96:25:@9397.4]
  assign _T_1742 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@9460.4 package.scala 96:25:@9461.4]
  assign _T_1746 = _T_1742 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9470.4]
  assign _T_1739 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@9452.4 package.scala 96:25:@9453.4]
  assign _T_1747 = _T_1739 ? Mem1D_6_io_output : _T_1746; // @[Mux.scala 31:69:@9471.4]
  assign _T_1736 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@9444.4 package.scala 96:25:@9445.4]
  assign _T_1777 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@9508.4 package.scala 96:25:@9509.4]
  assign _T_1781 = _T_1777 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@9518.4]
  assign _T_1774 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@9500.4 package.scala 96:25:@9501.4]
  assign _T_1782 = _T_1774 ? Mem1D_5_io_output : _T_1781; // @[Mux.scala 31:69:@9519.4]
  assign _T_1771 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@9492.4 package.scala 96:25:@9493.4]
  assign _T_1812 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@9556.4 package.scala 96:25:@9557.4]
  assign _T_1816 = _T_1812 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9566.4]
  assign _T_1809 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@9548.4 package.scala 96:25:@9549.4]
  assign _T_1817 = _T_1809 ? Mem1D_6_io_output : _T_1816; // @[Mux.scala 31:69:@9567.4]
  assign _T_1806 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@9540.4 package.scala 96:25:@9541.4]
  assign _T_1847 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@9604.4 package.scala 96:25:@9605.4]
  assign _T_1851 = _T_1847 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@9614.4]
  assign _T_1844 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@9596.4 package.scala 96:25:@9597.4]
  assign _T_1852 = _T_1844 ? Mem1D_6_io_output : _T_1851; // @[Mux.scala 31:69:@9615.4]
  assign _T_1841 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@9588.4 package.scala 96:25:@9589.4]
  assign _T_1882 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@9652.4 package.scala 96:25:@9653.4]
  assign _T_1886 = _T_1882 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9662.4]
  assign _T_1879 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@9644.4 package.scala 96:25:@9645.4]
  assign _T_1887 = _T_1879 ? Mem1D_7_io_output : _T_1886; // @[Mux.scala 31:69:@9663.4]
  assign _T_1876 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@9636.4 package.scala 96:25:@9637.4]
  assign _T_1917 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@9700.4 package.scala 96:25:@9701.4]
  assign _T_1921 = _T_1917 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@9710.4]
  assign _T_1914 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@9692.4 package.scala 96:25:@9693.4]
  assign _T_1922 = _T_1914 ? Mem1D_5_io_output : _T_1921; // @[Mux.scala 31:69:@9711.4]
  assign _T_1911 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@9684.4 package.scala 96:25:@9685.4]
  assign _T_1952 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@9748.4 package.scala 96:25:@9749.4]
  assign _T_1956 = _T_1952 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@9758.4]
  assign _T_1949 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@9740.4 package.scala 96:25:@9741.4]
  assign _T_1957 = _T_1949 ? Mem1D_5_io_output : _T_1956; // @[Mux.scala 31:69:@9759.4]
  assign _T_1946 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@9732.4 package.scala 96:25:@9733.4]
  assign _T_1987 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@9796.4 package.scala 96:25:@9797.4]
  assign _T_1991 = _T_1987 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@9806.4]
  assign _T_1984 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@9788.4 package.scala 96:25:@9789.4]
  assign _T_1992 = _T_1984 ? Mem1D_4_io_output : _T_1991; // @[Mux.scala 31:69:@9807.4]
  assign _T_1981 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@9780.4 package.scala 96:25:@9781.4]
  assign _T_2022 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@9844.4 package.scala 96:25:@9845.4]
  assign _T_2026 = _T_2022 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@9854.4]
  assign _T_2019 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@9836.4 package.scala 96:25:@9837.4]
  assign _T_2027 = _T_2019 ? Mem1D_4_io_output : _T_2026; // @[Mux.scala 31:69:@9855.4]
  assign _T_2016 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@9828.4 package.scala 96:25:@9829.4]
  assign _T_2057 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@9892.4 package.scala 96:25:@9893.4]
  assign _T_2061 = _T_2057 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9902.4]
  assign _T_2054 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@9884.4 package.scala 96:25:@9885.4]
  assign _T_2062 = _T_2054 ? Mem1D_7_io_output : _T_2061; // @[Mux.scala 31:69:@9903.4]
  assign _T_2051 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@9876.4 package.scala 96:25:@9877.4]
  assign _T_2092 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@9940.4 package.scala 96:25:@9941.4]
  assign _T_2096 = _T_2092 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@9950.4]
  assign _T_2089 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@9932.4 package.scala 96:25:@9933.4]
  assign _T_2097 = _T_2089 ? Mem1D_7_io_output : _T_2096; // @[Mux.scala 31:69:@9951.4]
  assign _T_2086 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@9924.4 package.scala 96:25:@9925.4]
  assign _T_2127 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@9988.4 package.scala 96:25:@9989.4]
  assign _T_2131 = _T_2127 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@9998.4]
  assign _T_2124 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@9980.4 package.scala 96:25:@9981.4]
  assign _T_2132 = _T_2124 ? Mem1D_4_io_output : _T_2131; // @[Mux.scala 31:69:@9999.4]
  assign _T_2121 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@9972.4 package.scala 96:25:@9973.4]
  assign _T_2162 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@10036.4 package.scala 96:25:@10037.4]
  assign _T_2166 = _T_2162 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@10046.4]
  assign _T_2159 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@10028.4 package.scala 96:25:@10029.4]
  assign _T_2167 = _T_2159 ? Mem1D_6_io_output : _T_2166; // @[Mux.scala 31:69:@10047.4]
  assign _T_2156 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@10020.4 package.scala 96:25:@10021.4]
  assign io_rPort_17_output_0 = _T_2156 ? Mem1D_2_io_output : _T_2167; // @[MemPrimitives.scala 148:13:@10049.4]
  assign io_rPort_16_output_0 = _T_2121 ? Mem1D_io_output : _T_2132; // @[MemPrimitives.scala 148:13:@10001.4]
  assign io_rPort_15_output_0 = _T_2086 ? Mem1D_3_io_output : _T_2097; // @[MemPrimitives.scala 148:13:@9953.4]
  assign io_rPort_14_output_0 = _T_2051 ? Mem1D_3_io_output : _T_2062; // @[MemPrimitives.scala 148:13:@9905.4]
  assign io_rPort_13_output_0 = _T_2016 ? Mem1D_io_output : _T_2027; // @[MemPrimitives.scala 148:13:@9857.4]
  assign io_rPort_12_output_0 = _T_1981 ? Mem1D_io_output : _T_1992; // @[MemPrimitives.scala 148:13:@9809.4]
  assign io_rPort_11_output_0 = _T_1946 ? Mem1D_1_io_output : _T_1957; // @[MemPrimitives.scala 148:13:@9761.4]
  assign io_rPort_10_output_0 = _T_1911 ? Mem1D_1_io_output : _T_1922; // @[MemPrimitives.scala 148:13:@9713.4]
  assign io_rPort_9_output_0 = _T_1876 ? Mem1D_3_io_output : _T_1887; // @[MemPrimitives.scala 148:13:@9665.4]
  assign io_rPort_8_output_0 = _T_1841 ? Mem1D_2_io_output : _T_1852; // @[MemPrimitives.scala 148:13:@9617.4]
  assign io_rPort_7_output_0 = _T_1806 ? Mem1D_2_io_output : _T_1817; // @[MemPrimitives.scala 148:13:@9569.4]
  assign io_rPort_6_output_0 = _T_1771 ? Mem1D_1_io_output : _T_1782; // @[MemPrimitives.scala 148:13:@9521.4]
  assign io_rPort_5_output_0 = _T_1736 ? Mem1D_2_io_output : _T_1747; // @[MemPrimitives.scala 148:13:@9473.4]
  assign io_rPort_4_output_0 = _T_1701 ? Mem1D_3_io_output : _T_1712; // @[MemPrimitives.scala 148:13:@9425.4]
  assign io_rPort_3_output_0 = _T_1666 ? Mem1D_3_io_output : _T_1677; // @[MemPrimitives.scala 148:13:@9377.4]
  assign io_rPort_2_output_0 = _T_1631 ? Mem1D_2_io_output : _T_1642; // @[MemPrimitives.scala 148:13:@9329.4]
  assign io_rPort_1_output_0 = _T_1596 ? Mem1D_2_io_output : _T_1607; // @[MemPrimitives.scala 148:13:@9281.4]
  assign io_rPort_0_output_0 = _T_1561 ? Mem1D_3_io_output : _T_1572; // @[MemPrimitives.scala 148:13:@9233.4]
  assign Mem1D_clock = clock; // @[:@8051.4]
  assign Mem1D_reset = reset; // @[:@8052.4]
  assign Mem1D_io_r_ofs_0 = _T_884[0]; // @[MemPrimitives.scala 127:28:@8511.4]
  assign Mem1D_io_r_backpressure = _T_884[1]; // @[MemPrimitives.scala 128:32:@8512.4]
  assign Mem1D_io_w_ofs_0 = _T_705[0]; // @[MemPrimitives.scala 94:28:@8314.4]
  assign Mem1D_io_w_data_0 = _T_705[8:1]; // @[MemPrimitives.scala 95:29:@8315.4]
  assign Mem1D_io_w_en_0 = _T_705[9]; // @[MemPrimitives.scala 96:27:@8316.4]
  assign Mem1D_1_clock = clock; // @[:@8067.4]
  assign Mem1D_1_reset = reset; // @[:@8068.4]
  assign Mem1D_1_io_r_ofs_0 = _T_913[0]; // @[MemPrimitives.scala 127:28:@8543.4]
  assign Mem1D_1_io_r_backpressure = _T_913[1]; // @[MemPrimitives.scala 128:32:@8544.4]
  assign Mem1D_1_io_w_ofs_0 = _T_715[0]; // @[MemPrimitives.scala 94:28:@8325.4]
  assign Mem1D_1_io_w_data_0 = _T_715[8:1]; // @[MemPrimitives.scala 95:29:@8326.4]
  assign Mem1D_1_io_w_en_0 = _T_715[9]; // @[MemPrimitives.scala 96:27:@8327.4]
  assign Mem1D_2_clock = clock; // @[:@8083.4]
  assign Mem1D_2_reset = reset; // @[:@8084.4]
  assign Mem1D_2_io_r_ofs_0 = _T_969[0]; // @[MemPrimitives.scala 127:28:@8599.4]
  assign Mem1D_2_io_r_backpressure = _T_969[1]; // @[MemPrimitives.scala 128:32:@8600.4]
  assign Mem1D_2_io_w_ofs_0 = _T_725[0]; // @[MemPrimitives.scala 94:28:@8336.4]
  assign Mem1D_2_io_w_data_0 = _T_725[8:1]; // @[MemPrimitives.scala 95:29:@8337.4]
  assign Mem1D_2_io_w_en_0 = _T_725[9]; // @[MemPrimitives.scala 96:27:@8338.4]
  assign Mem1D_3_clock = clock; // @[:@8099.4]
  assign Mem1D_3_reset = reset; // @[:@8100.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1025[0]; // @[MemPrimitives.scala 127:28:@8655.4]
  assign Mem1D_3_io_r_backpressure = _T_1025[1]; // @[MemPrimitives.scala 128:32:@8656.4]
  assign Mem1D_3_io_w_ofs_0 = _T_735[0]; // @[MemPrimitives.scala 94:28:@8347.4]
  assign Mem1D_3_io_w_data_0 = _T_735[8:1]; // @[MemPrimitives.scala 95:29:@8348.4]
  assign Mem1D_3_io_w_en_0 = _T_735[9]; // @[MemPrimitives.scala 96:27:@8349.4]
  assign Mem1D_4_clock = clock; // @[:@8115.4]
  assign Mem1D_4_reset = reset; // @[:@8116.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1054[0]; // @[MemPrimitives.scala 127:28:@8687.4]
  assign Mem1D_4_io_r_backpressure = _T_1054[1]; // @[MemPrimitives.scala 128:32:@8688.4]
  assign Mem1D_4_io_w_ofs_0 = _T_745[0]; // @[MemPrimitives.scala 94:28:@8358.4]
  assign Mem1D_4_io_w_data_0 = _T_745[8:1]; // @[MemPrimitives.scala 95:29:@8359.4]
  assign Mem1D_4_io_w_en_0 = _T_745[9]; // @[MemPrimitives.scala 96:27:@8360.4]
  assign Mem1D_5_clock = clock; // @[:@8131.4]
  assign Mem1D_5_reset = reset; // @[:@8132.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1083[0]; // @[MemPrimitives.scala 127:28:@8719.4]
  assign Mem1D_5_io_r_backpressure = _T_1083[1]; // @[MemPrimitives.scala 128:32:@8720.4]
  assign Mem1D_5_io_w_ofs_0 = _T_755[0]; // @[MemPrimitives.scala 94:28:@8369.4]
  assign Mem1D_5_io_w_data_0 = _T_755[8:1]; // @[MemPrimitives.scala 95:29:@8370.4]
  assign Mem1D_5_io_w_en_0 = _T_755[9]; // @[MemPrimitives.scala 96:27:@8371.4]
  assign Mem1D_6_clock = clock; // @[:@8147.4]
  assign Mem1D_6_reset = reset; // @[:@8148.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1139[0]; // @[MemPrimitives.scala 127:28:@8775.4]
  assign Mem1D_6_io_r_backpressure = _T_1139[1]; // @[MemPrimitives.scala 128:32:@8776.4]
  assign Mem1D_6_io_w_ofs_0 = _T_765[0]; // @[MemPrimitives.scala 94:28:@8380.4]
  assign Mem1D_6_io_w_data_0 = _T_765[8:1]; // @[MemPrimitives.scala 95:29:@8381.4]
  assign Mem1D_6_io_w_en_0 = _T_765[9]; // @[MemPrimitives.scala 96:27:@8382.4]
  assign Mem1D_7_clock = clock; // @[:@8163.4]
  assign Mem1D_7_reset = reset; // @[:@8164.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1195[0]; // @[MemPrimitives.scala 127:28:@8831.4]
  assign Mem1D_7_io_r_backpressure = _T_1195[1]; // @[MemPrimitives.scala 128:32:@8832.4]
  assign Mem1D_7_io_w_ofs_0 = _T_775[0]; // @[MemPrimitives.scala 94:28:@8391.4]
  assign Mem1D_7_io_w_data_0 = _T_775[8:1]; // @[MemPrimitives.scala 95:29:@8392.4]
  assign Mem1D_7_io_w_en_0 = _T_775[9]; // @[MemPrimitives.scala 96:27:@8393.4]
  assign Mem1D_8_clock = clock; // @[:@8179.4]
  assign Mem1D_8_reset = reset; // @[:@8180.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1224[0]; // @[MemPrimitives.scala 127:28:@8863.4]
  assign Mem1D_8_io_r_backpressure = _T_1224[1]; // @[MemPrimitives.scala 128:32:@8864.4]
  assign Mem1D_8_io_w_ofs_0 = _T_785[0]; // @[MemPrimitives.scala 94:28:@8402.4]
  assign Mem1D_8_io_w_data_0 = _T_785[8:1]; // @[MemPrimitives.scala 95:29:@8403.4]
  assign Mem1D_8_io_w_en_0 = _T_785[9]; // @[MemPrimitives.scala 96:27:@8404.4]
  assign Mem1D_9_clock = clock; // @[:@8195.4]
  assign Mem1D_9_reset = reset; // @[:@8196.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1253[0]; // @[MemPrimitives.scala 127:28:@8895.4]
  assign Mem1D_9_io_r_backpressure = _T_1253[1]; // @[MemPrimitives.scala 128:32:@8896.4]
  assign Mem1D_9_io_w_ofs_0 = _T_795[0]; // @[MemPrimitives.scala 94:28:@8413.4]
  assign Mem1D_9_io_w_data_0 = _T_795[8:1]; // @[MemPrimitives.scala 95:29:@8414.4]
  assign Mem1D_9_io_w_en_0 = _T_795[9]; // @[MemPrimitives.scala 96:27:@8415.4]
  assign Mem1D_10_clock = clock; // @[:@8211.4]
  assign Mem1D_10_reset = reset; // @[:@8212.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1309[0]; // @[MemPrimitives.scala 127:28:@8951.4]
  assign Mem1D_10_io_r_backpressure = _T_1309[1]; // @[MemPrimitives.scala 128:32:@8952.4]
  assign Mem1D_10_io_w_ofs_0 = _T_805[0]; // @[MemPrimitives.scala 94:28:@8424.4]
  assign Mem1D_10_io_w_data_0 = _T_805[8:1]; // @[MemPrimitives.scala 95:29:@8425.4]
  assign Mem1D_10_io_w_en_0 = _T_805[9]; // @[MemPrimitives.scala 96:27:@8426.4]
  assign Mem1D_11_clock = clock; // @[:@8227.4]
  assign Mem1D_11_reset = reset; // @[:@8228.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1365[0]; // @[MemPrimitives.scala 127:28:@9007.4]
  assign Mem1D_11_io_r_backpressure = _T_1365[1]; // @[MemPrimitives.scala 128:32:@9008.4]
  assign Mem1D_11_io_w_ofs_0 = _T_815[0]; // @[MemPrimitives.scala 94:28:@8435.4]
  assign Mem1D_11_io_w_data_0 = _T_815[8:1]; // @[MemPrimitives.scala 95:29:@8436.4]
  assign Mem1D_11_io_w_en_0 = _T_815[9]; // @[MemPrimitives.scala 96:27:@8437.4]
  assign Mem1D_12_clock = clock; // @[:@8243.4]
  assign Mem1D_12_reset = reset; // @[:@8244.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1394[0]; // @[MemPrimitives.scala 127:28:@9039.4]
  assign Mem1D_12_io_r_backpressure = _T_1394[1]; // @[MemPrimitives.scala 128:32:@9040.4]
  assign Mem1D_12_io_w_ofs_0 = _T_825[0]; // @[MemPrimitives.scala 94:28:@8446.4]
  assign Mem1D_12_io_w_data_0 = _T_825[8:1]; // @[MemPrimitives.scala 95:29:@8447.4]
  assign Mem1D_12_io_w_en_0 = _T_825[9]; // @[MemPrimitives.scala 96:27:@8448.4]
  assign Mem1D_13_clock = clock; // @[:@8259.4]
  assign Mem1D_13_reset = reset; // @[:@8260.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1423[0]; // @[MemPrimitives.scala 127:28:@9071.4]
  assign Mem1D_13_io_r_backpressure = _T_1423[1]; // @[MemPrimitives.scala 128:32:@9072.4]
  assign Mem1D_13_io_w_ofs_0 = _T_835[0]; // @[MemPrimitives.scala 94:28:@8457.4]
  assign Mem1D_13_io_w_data_0 = _T_835[8:1]; // @[MemPrimitives.scala 95:29:@8458.4]
  assign Mem1D_13_io_w_en_0 = _T_835[9]; // @[MemPrimitives.scala 96:27:@8459.4]
  assign Mem1D_14_clock = clock; // @[:@8275.4]
  assign Mem1D_14_reset = reset; // @[:@8276.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1479[0]; // @[MemPrimitives.scala 127:28:@9127.4]
  assign Mem1D_14_io_r_backpressure = _T_1479[1]; // @[MemPrimitives.scala 128:32:@9128.4]
  assign Mem1D_14_io_w_ofs_0 = _T_845[0]; // @[MemPrimitives.scala 94:28:@8468.4]
  assign Mem1D_14_io_w_data_0 = _T_845[8:1]; // @[MemPrimitives.scala 95:29:@8469.4]
  assign Mem1D_14_io_w_en_0 = _T_845[9]; // @[MemPrimitives.scala 96:27:@8470.4]
  assign Mem1D_15_clock = clock; // @[:@8291.4]
  assign Mem1D_15_reset = reset; // @[:@8292.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1535[0]; // @[MemPrimitives.scala 127:28:@9183.4]
  assign Mem1D_15_io_r_backpressure = _T_1535[1]; // @[MemPrimitives.scala 128:32:@9184.4]
  assign Mem1D_15_io_w_ofs_0 = _T_855[0]; // @[MemPrimitives.scala 94:28:@8479.4]
  assign Mem1D_15_io_w_data_0 = _T_855[8:1]; // @[MemPrimitives.scala 95:29:@8480.4]
  assign Mem1D_15_io_w_en_0 = _T_855[9]; // @[MemPrimitives.scala 96:27:@8481.4]
  assign StickySelects_clock = clock; // @[:@8492.4]
  assign StickySelects_reset = reset; // @[:@8493.4]
  assign StickySelects_io_ins_0 = io_rPort_12_en_0 & _T_860; // @[MemPrimitives.scala 122:60:@8494.4]
  assign StickySelects_io_ins_1 = io_rPort_13_en_0 & _T_865; // @[MemPrimitives.scala 122:60:@8495.4]
  assign StickySelects_io_ins_2 = io_rPort_16_en_0 & _T_870; // @[MemPrimitives.scala 122:60:@8496.4]
  assign StickySelects_1_clock = clock; // @[:@8524.4]
  assign StickySelects_1_reset = reset; // @[:@8525.4]
  assign StickySelects_1_io_ins_0 = io_rPort_6_en_0 & _T_889; // @[MemPrimitives.scala 122:60:@8526.4]
  assign StickySelects_1_io_ins_1 = io_rPort_10_en_0 & _T_894; // @[MemPrimitives.scala 122:60:@8527.4]
  assign StickySelects_1_io_ins_2 = io_rPort_11_en_0 & _T_899; // @[MemPrimitives.scala 122:60:@8528.4]
  assign StickySelects_2_clock = clock; // @[:@8565.4]
  assign StickySelects_2_reset = reset; // @[:@8566.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_918; // @[MemPrimitives.scala 122:60:@8567.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 122:60:@8568.4]
  assign StickySelects_2_io_ins_2 = io_rPort_5_en_0 & _T_928; // @[MemPrimitives.scala 122:60:@8569.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_933; // @[MemPrimitives.scala 122:60:@8570.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_938; // @[MemPrimitives.scala 122:60:@8571.4]
  assign StickySelects_2_io_ins_5 = io_rPort_17_en_0 & _T_943; // @[MemPrimitives.scala 122:60:@8572.4]
  assign StickySelects_3_clock = clock; // @[:@8621.4]
  assign StickySelects_3_reset = reset; // @[:@8622.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_974; // @[MemPrimitives.scala 122:60:@8623.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_979; // @[MemPrimitives.scala 122:60:@8624.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_984; // @[MemPrimitives.scala 122:60:@8625.4]
  assign StickySelects_3_io_ins_3 = io_rPort_9_en_0 & _T_989; // @[MemPrimitives.scala 122:60:@8626.4]
  assign StickySelects_3_io_ins_4 = io_rPort_14_en_0 & _T_994; // @[MemPrimitives.scala 122:60:@8627.4]
  assign StickySelects_3_io_ins_5 = io_rPort_15_en_0 & _T_999; // @[MemPrimitives.scala 122:60:@8628.4]
  assign StickySelects_4_clock = clock; // @[:@8668.4]
  assign StickySelects_4_reset = reset; // @[:@8669.4]
  assign StickySelects_4_io_ins_0 = io_rPort_12_en_0 & _T_1030; // @[MemPrimitives.scala 122:60:@8670.4]
  assign StickySelects_4_io_ins_1 = io_rPort_13_en_0 & _T_1035; // @[MemPrimitives.scala 122:60:@8671.4]
  assign StickySelects_4_io_ins_2 = io_rPort_16_en_0 & _T_1040; // @[MemPrimitives.scala 122:60:@8672.4]
  assign StickySelects_5_clock = clock; // @[:@8700.4]
  assign StickySelects_5_reset = reset; // @[:@8701.4]
  assign StickySelects_5_io_ins_0 = io_rPort_6_en_0 & _T_1059; // @[MemPrimitives.scala 122:60:@8702.4]
  assign StickySelects_5_io_ins_1 = io_rPort_10_en_0 & _T_1064; // @[MemPrimitives.scala 122:60:@8703.4]
  assign StickySelects_5_io_ins_2 = io_rPort_11_en_0 & _T_1069; // @[MemPrimitives.scala 122:60:@8704.4]
  assign StickySelects_6_clock = clock; // @[:@8741.4]
  assign StickySelects_6_reset = reset; // @[:@8742.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_1088; // @[MemPrimitives.scala 122:60:@8743.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_1093; // @[MemPrimitives.scala 122:60:@8744.4]
  assign StickySelects_6_io_ins_2 = io_rPort_5_en_0 & _T_1098; // @[MemPrimitives.scala 122:60:@8745.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1103; // @[MemPrimitives.scala 122:60:@8746.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1108; // @[MemPrimitives.scala 122:60:@8747.4]
  assign StickySelects_6_io_ins_5 = io_rPort_17_en_0 & _T_1113; // @[MemPrimitives.scala 122:60:@8748.4]
  assign StickySelects_7_clock = clock; // @[:@8797.4]
  assign StickySelects_7_reset = reset; // @[:@8798.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1144; // @[MemPrimitives.scala 122:60:@8799.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_1149; // @[MemPrimitives.scala 122:60:@8800.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_1154; // @[MemPrimitives.scala 122:60:@8801.4]
  assign StickySelects_7_io_ins_3 = io_rPort_9_en_0 & _T_1159; // @[MemPrimitives.scala 122:60:@8802.4]
  assign StickySelects_7_io_ins_4 = io_rPort_14_en_0 & _T_1164; // @[MemPrimitives.scala 122:60:@8803.4]
  assign StickySelects_7_io_ins_5 = io_rPort_15_en_0 & _T_1169; // @[MemPrimitives.scala 122:60:@8804.4]
  assign StickySelects_8_clock = clock; // @[:@8844.4]
  assign StickySelects_8_reset = reset; // @[:@8845.4]
  assign StickySelects_8_io_ins_0 = io_rPort_12_en_0 & _T_1200; // @[MemPrimitives.scala 122:60:@8846.4]
  assign StickySelects_8_io_ins_1 = io_rPort_13_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@8847.4]
  assign StickySelects_8_io_ins_2 = io_rPort_16_en_0 & _T_1210; // @[MemPrimitives.scala 122:60:@8848.4]
  assign StickySelects_9_clock = clock; // @[:@8876.4]
  assign StickySelects_9_reset = reset; // @[:@8877.4]
  assign StickySelects_9_io_ins_0 = io_rPort_6_en_0 & _T_1229; // @[MemPrimitives.scala 122:60:@8878.4]
  assign StickySelects_9_io_ins_1 = io_rPort_10_en_0 & _T_1234; // @[MemPrimitives.scala 122:60:@8879.4]
  assign StickySelects_9_io_ins_2 = io_rPort_11_en_0 & _T_1239; // @[MemPrimitives.scala 122:60:@8880.4]
  assign StickySelects_10_clock = clock; // @[:@8917.4]
  assign StickySelects_10_reset = reset; // @[:@8918.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_1258; // @[MemPrimitives.scala 122:60:@8919.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_1263; // @[MemPrimitives.scala 122:60:@8920.4]
  assign StickySelects_10_io_ins_2 = io_rPort_5_en_0 & _T_1268; // @[MemPrimitives.scala 122:60:@8921.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@8922.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_1278; // @[MemPrimitives.scala 122:60:@8923.4]
  assign StickySelects_10_io_ins_5 = io_rPort_17_en_0 & _T_1283; // @[MemPrimitives.scala 122:60:@8924.4]
  assign StickySelects_11_clock = clock; // @[:@8973.4]
  assign StickySelects_11_reset = reset; // @[:@8974.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1314; // @[MemPrimitives.scala 122:60:@8975.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_1319; // @[MemPrimitives.scala 122:60:@8976.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_1324; // @[MemPrimitives.scala 122:60:@8977.4]
  assign StickySelects_11_io_ins_3 = io_rPort_9_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@8978.4]
  assign StickySelects_11_io_ins_4 = io_rPort_14_en_0 & _T_1334; // @[MemPrimitives.scala 122:60:@8979.4]
  assign StickySelects_11_io_ins_5 = io_rPort_15_en_0 & _T_1339; // @[MemPrimitives.scala 122:60:@8980.4]
  assign StickySelects_12_clock = clock; // @[:@9020.4]
  assign StickySelects_12_reset = reset; // @[:@9021.4]
  assign StickySelects_12_io_ins_0 = io_rPort_12_en_0 & _T_1370; // @[MemPrimitives.scala 122:60:@9022.4]
  assign StickySelects_12_io_ins_1 = io_rPort_13_en_0 & _T_1375; // @[MemPrimitives.scala 122:60:@9023.4]
  assign StickySelects_12_io_ins_2 = io_rPort_16_en_0 & _T_1380; // @[MemPrimitives.scala 122:60:@9024.4]
  assign StickySelects_13_clock = clock; // @[:@9052.4]
  assign StickySelects_13_reset = reset; // @[:@9053.4]
  assign StickySelects_13_io_ins_0 = io_rPort_6_en_0 & _T_1399; // @[MemPrimitives.scala 122:60:@9054.4]
  assign StickySelects_13_io_ins_1 = io_rPort_10_en_0 & _T_1404; // @[MemPrimitives.scala 122:60:@9055.4]
  assign StickySelects_13_io_ins_2 = io_rPort_11_en_0 & _T_1409; // @[MemPrimitives.scala 122:60:@9056.4]
  assign StickySelects_14_clock = clock; // @[:@9093.4]
  assign StickySelects_14_reset = reset; // @[:@9094.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_1428; // @[MemPrimitives.scala 122:60:@9095.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_1433; // @[MemPrimitives.scala 122:60:@9096.4]
  assign StickySelects_14_io_ins_2 = io_rPort_5_en_0 & _T_1438; // @[MemPrimitives.scala 122:60:@9097.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_1443; // @[MemPrimitives.scala 122:60:@9098.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_1448; // @[MemPrimitives.scala 122:60:@9099.4]
  assign StickySelects_14_io_ins_5 = io_rPort_17_en_0 & _T_1453; // @[MemPrimitives.scala 122:60:@9100.4]
  assign StickySelects_15_clock = clock; // @[:@9149.4]
  assign StickySelects_15_reset = reset; // @[:@9150.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1484; // @[MemPrimitives.scala 122:60:@9151.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_1489; // @[MemPrimitives.scala 122:60:@9152.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_1494; // @[MemPrimitives.scala 122:60:@9153.4]
  assign StickySelects_15_io_ins_3 = io_rPort_9_en_0 & _T_1499; // @[MemPrimitives.scala 122:60:@9154.4]
  assign StickySelects_15_io_ins_4 = io_rPort_14_en_0 & _T_1504; // @[MemPrimitives.scala 122:60:@9155.4]
  assign StickySelects_15_io_ins_5 = io_rPort_15_en_0 & _T_1509; // @[MemPrimitives.scala 122:60:@9156.4]
  assign RetimeWrapper_clock = clock; // @[:@9200.4]
  assign RetimeWrapper_reset = reset; // @[:@9201.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9203.4]
  assign RetimeWrapper_io_in = _T_974 & io_rPort_0_en_0; // @[package.scala 94:16:@9202.4]
  assign RetimeWrapper_1_clock = clock; // @[:@9208.4]
  assign RetimeWrapper_1_reset = reset; // @[:@9209.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9211.4]
  assign RetimeWrapper_1_io_in = _T_1144 & io_rPort_0_en_0; // @[package.scala 94:16:@9210.4]
  assign RetimeWrapper_2_clock = clock; // @[:@9216.4]
  assign RetimeWrapper_2_reset = reset; // @[:@9217.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9219.4]
  assign RetimeWrapper_2_io_in = _T_1314 & io_rPort_0_en_0; // @[package.scala 94:16:@9218.4]
  assign RetimeWrapper_3_clock = clock; // @[:@9224.4]
  assign RetimeWrapper_3_reset = reset; // @[:@9225.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@9227.4]
  assign RetimeWrapper_3_io_in = _T_1484 & io_rPort_0_en_0; // @[package.scala 94:16:@9226.4]
  assign RetimeWrapper_4_clock = clock; // @[:@9248.4]
  assign RetimeWrapper_4_reset = reset; // @[:@9249.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9251.4]
  assign RetimeWrapper_4_io_in = _T_918 & io_rPort_1_en_0; // @[package.scala 94:16:@9250.4]
  assign RetimeWrapper_5_clock = clock; // @[:@9256.4]
  assign RetimeWrapper_5_reset = reset; // @[:@9257.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9259.4]
  assign RetimeWrapper_5_io_in = _T_1088 & io_rPort_1_en_0; // @[package.scala 94:16:@9258.4]
  assign RetimeWrapper_6_clock = clock; // @[:@9264.4]
  assign RetimeWrapper_6_reset = reset; // @[:@9265.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9267.4]
  assign RetimeWrapper_6_io_in = _T_1258 & io_rPort_1_en_0; // @[package.scala 94:16:@9266.4]
  assign RetimeWrapper_7_clock = clock; // @[:@9272.4]
  assign RetimeWrapper_7_reset = reset; // @[:@9273.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@9275.4]
  assign RetimeWrapper_7_io_in = _T_1428 & io_rPort_1_en_0; // @[package.scala 94:16:@9274.4]
  assign RetimeWrapper_8_clock = clock; // @[:@9296.4]
  assign RetimeWrapper_8_reset = reset; // @[:@9297.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9299.4]
  assign RetimeWrapper_8_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@9298.4]
  assign RetimeWrapper_9_clock = clock; // @[:@9304.4]
  assign RetimeWrapper_9_reset = reset; // @[:@9305.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9307.4]
  assign RetimeWrapper_9_io_in = _T_1093 & io_rPort_2_en_0; // @[package.scala 94:16:@9306.4]
  assign RetimeWrapper_10_clock = clock; // @[:@9312.4]
  assign RetimeWrapper_10_reset = reset; // @[:@9313.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9315.4]
  assign RetimeWrapper_10_io_in = _T_1263 & io_rPort_2_en_0; // @[package.scala 94:16:@9314.4]
  assign RetimeWrapper_11_clock = clock; // @[:@9320.4]
  assign RetimeWrapper_11_reset = reset; // @[:@9321.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@9323.4]
  assign RetimeWrapper_11_io_in = _T_1433 & io_rPort_2_en_0; // @[package.scala 94:16:@9322.4]
  assign RetimeWrapper_12_clock = clock; // @[:@9344.4]
  assign RetimeWrapper_12_reset = reset; // @[:@9345.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9347.4]
  assign RetimeWrapper_12_io_in = _T_979 & io_rPort_3_en_0; // @[package.scala 94:16:@9346.4]
  assign RetimeWrapper_13_clock = clock; // @[:@9352.4]
  assign RetimeWrapper_13_reset = reset; // @[:@9353.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9355.4]
  assign RetimeWrapper_13_io_in = _T_1149 & io_rPort_3_en_0; // @[package.scala 94:16:@9354.4]
  assign RetimeWrapper_14_clock = clock; // @[:@9360.4]
  assign RetimeWrapper_14_reset = reset; // @[:@9361.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9363.4]
  assign RetimeWrapper_14_io_in = _T_1319 & io_rPort_3_en_0; // @[package.scala 94:16:@9362.4]
  assign RetimeWrapper_15_clock = clock; // @[:@9368.4]
  assign RetimeWrapper_15_reset = reset; // @[:@9369.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@9371.4]
  assign RetimeWrapper_15_io_in = _T_1489 & io_rPort_3_en_0; // @[package.scala 94:16:@9370.4]
  assign RetimeWrapper_16_clock = clock; // @[:@9392.4]
  assign RetimeWrapper_16_reset = reset; // @[:@9393.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9395.4]
  assign RetimeWrapper_16_io_in = _T_984 & io_rPort_4_en_0; // @[package.scala 94:16:@9394.4]
  assign RetimeWrapper_17_clock = clock; // @[:@9400.4]
  assign RetimeWrapper_17_reset = reset; // @[:@9401.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9403.4]
  assign RetimeWrapper_17_io_in = _T_1154 & io_rPort_4_en_0; // @[package.scala 94:16:@9402.4]
  assign RetimeWrapper_18_clock = clock; // @[:@9408.4]
  assign RetimeWrapper_18_reset = reset; // @[:@9409.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9411.4]
  assign RetimeWrapper_18_io_in = _T_1324 & io_rPort_4_en_0; // @[package.scala 94:16:@9410.4]
  assign RetimeWrapper_19_clock = clock; // @[:@9416.4]
  assign RetimeWrapper_19_reset = reset; // @[:@9417.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@9419.4]
  assign RetimeWrapper_19_io_in = _T_1494 & io_rPort_4_en_0; // @[package.scala 94:16:@9418.4]
  assign RetimeWrapper_20_clock = clock; // @[:@9440.4]
  assign RetimeWrapper_20_reset = reset; // @[:@9441.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9443.4]
  assign RetimeWrapper_20_io_in = _T_928 & io_rPort_5_en_0; // @[package.scala 94:16:@9442.4]
  assign RetimeWrapper_21_clock = clock; // @[:@9448.4]
  assign RetimeWrapper_21_reset = reset; // @[:@9449.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9451.4]
  assign RetimeWrapper_21_io_in = _T_1098 & io_rPort_5_en_0; // @[package.scala 94:16:@9450.4]
  assign RetimeWrapper_22_clock = clock; // @[:@9456.4]
  assign RetimeWrapper_22_reset = reset; // @[:@9457.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9459.4]
  assign RetimeWrapper_22_io_in = _T_1268 & io_rPort_5_en_0; // @[package.scala 94:16:@9458.4]
  assign RetimeWrapper_23_clock = clock; // @[:@9464.4]
  assign RetimeWrapper_23_reset = reset; // @[:@9465.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@9467.4]
  assign RetimeWrapper_23_io_in = _T_1438 & io_rPort_5_en_0; // @[package.scala 94:16:@9466.4]
  assign RetimeWrapper_24_clock = clock; // @[:@9488.4]
  assign RetimeWrapper_24_reset = reset; // @[:@9489.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9491.4]
  assign RetimeWrapper_24_io_in = _T_889 & io_rPort_6_en_0; // @[package.scala 94:16:@9490.4]
  assign RetimeWrapper_25_clock = clock; // @[:@9496.4]
  assign RetimeWrapper_25_reset = reset; // @[:@9497.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9499.4]
  assign RetimeWrapper_25_io_in = _T_1059 & io_rPort_6_en_0; // @[package.scala 94:16:@9498.4]
  assign RetimeWrapper_26_clock = clock; // @[:@9504.4]
  assign RetimeWrapper_26_reset = reset; // @[:@9505.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9507.4]
  assign RetimeWrapper_26_io_in = _T_1229 & io_rPort_6_en_0; // @[package.scala 94:16:@9506.4]
  assign RetimeWrapper_27_clock = clock; // @[:@9512.4]
  assign RetimeWrapper_27_reset = reset; // @[:@9513.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@9515.4]
  assign RetimeWrapper_27_io_in = _T_1399 & io_rPort_6_en_0; // @[package.scala 94:16:@9514.4]
  assign RetimeWrapper_28_clock = clock; // @[:@9536.4]
  assign RetimeWrapper_28_reset = reset; // @[:@9537.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9539.4]
  assign RetimeWrapper_28_io_in = _T_933 & io_rPort_7_en_0; // @[package.scala 94:16:@9538.4]
  assign RetimeWrapper_29_clock = clock; // @[:@9544.4]
  assign RetimeWrapper_29_reset = reset; // @[:@9545.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9547.4]
  assign RetimeWrapper_29_io_in = _T_1103 & io_rPort_7_en_0; // @[package.scala 94:16:@9546.4]
  assign RetimeWrapper_30_clock = clock; // @[:@9552.4]
  assign RetimeWrapper_30_reset = reset; // @[:@9553.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9555.4]
  assign RetimeWrapper_30_io_in = _T_1273 & io_rPort_7_en_0; // @[package.scala 94:16:@9554.4]
  assign RetimeWrapper_31_clock = clock; // @[:@9560.4]
  assign RetimeWrapper_31_reset = reset; // @[:@9561.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@9563.4]
  assign RetimeWrapper_31_io_in = _T_1443 & io_rPort_7_en_0; // @[package.scala 94:16:@9562.4]
  assign RetimeWrapper_32_clock = clock; // @[:@9584.4]
  assign RetimeWrapper_32_reset = reset; // @[:@9585.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9587.4]
  assign RetimeWrapper_32_io_in = _T_938 & io_rPort_8_en_0; // @[package.scala 94:16:@9586.4]
  assign RetimeWrapper_33_clock = clock; // @[:@9592.4]
  assign RetimeWrapper_33_reset = reset; // @[:@9593.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9595.4]
  assign RetimeWrapper_33_io_in = _T_1108 & io_rPort_8_en_0; // @[package.scala 94:16:@9594.4]
  assign RetimeWrapper_34_clock = clock; // @[:@9600.4]
  assign RetimeWrapper_34_reset = reset; // @[:@9601.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9603.4]
  assign RetimeWrapper_34_io_in = _T_1278 & io_rPort_8_en_0; // @[package.scala 94:16:@9602.4]
  assign RetimeWrapper_35_clock = clock; // @[:@9608.4]
  assign RetimeWrapper_35_reset = reset; // @[:@9609.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@9611.4]
  assign RetimeWrapper_35_io_in = _T_1448 & io_rPort_8_en_0; // @[package.scala 94:16:@9610.4]
  assign RetimeWrapper_36_clock = clock; // @[:@9632.4]
  assign RetimeWrapper_36_reset = reset; // @[:@9633.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9635.4]
  assign RetimeWrapper_36_io_in = _T_989 & io_rPort_9_en_0; // @[package.scala 94:16:@9634.4]
  assign RetimeWrapper_37_clock = clock; // @[:@9640.4]
  assign RetimeWrapper_37_reset = reset; // @[:@9641.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9643.4]
  assign RetimeWrapper_37_io_in = _T_1159 & io_rPort_9_en_0; // @[package.scala 94:16:@9642.4]
  assign RetimeWrapper_38_clock = clock; // @[:@9648.4]
  assign RetimeWrapper_38_reset = reset; // @[:@9649.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9651.4]
  assign RetimeWrapper_38_io_in = _T_1329 & io_rPort_9_en_0; // @[package.scala 94:16:@9650.4]
  assign RetimeWrapper_39_clock = clock; // @[:@9656.4]
  assign RetimeWrapper_39_reset = reset; // @[:@9657.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@9659.4]
  assign RetimeWrapper_39_io_in = _T_1499 & io_rPort_9_en_0; // @[package.scala 94:16:@9658.4]
  assign RetimeWrapper_40_clock = clock; // @[:@9680.4]
  assign RetimeWrapper_40_reset = reset; // @[:@9681.4]
  assign RetimeWrapper_40_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9683.4]
  assign RetimeWrapper_40_io_in = _T_894 & io_rPort_10_en_0; // @[package.scala 94:16:@9682.4]
  assign RetimeWrapper_41_clock = clock; // @[:@9688.4]
  assign RetimeWrapper_41_reset = reset; // @[:@9689.4]
  assign RetimeWrapper_41_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9691.4]
  assign RetimeWrapper_41_io_in = _T_1064 & io_rPort_10_en_0; // @[package.scala 94:16:@9690.4]
  assign RetimeWrapper_42_clock = clock; // @[:@9696.4]
  assign RetimeWrapper_42_reset = reset; // @[:@9697.4]
  assign RetimeWrapper_42_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9699.4]
  assign RetimeWrapper_42_io_in = _T_1234 & io_rPort_10_en_0; // @[package.scala 94:16:@9698.4]
  assign RetimeWrapper_43_clock = clock; // @[:@9704.4]
  assign RetimeWrapper_43_reset = reset; // @[:@9705.4]
  assign RetimeWrapper_43_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@9707.4]
  assign RetimeWrapper_43_io_in = _T_1404 & io_rPort_10_en_0; // @[package.scala 94:16:@9706.4]
  assign RetimeWrapper_44_clock = clock; // @[:@9728.4]
  assign RetimeWrapper_44_reset = reset; // @[:@9729.4]
  assign RetimeWrapper_44_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9731.4]
  assign RetimeWrapper_44_io_in = _T_899 & io_rPort_11_en_0; // @[package.scala 94:16:@9730.4]
  assign RetimeWrapper_45_clock = clock; // @[:@9736.4]
  assign RetimeWrapper_45_reset = reset; // @[:@9737.4]
  assign RetimeWrapper_45_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9739.4]
  assign RetimeWrapper_45_io_in = _T_1069 & io_rPort_11_en_0; // @[package.scala 94:16:@9738.4]
  assign RetimeWrapper_46_clock = clock; // @[:@9744.4]
  assign RetimeWrapper_46_reset = reset; // @[:@9745.4]
  assign RetimeWrapper_46_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9747.4]
  assign RetimeWrapper_46_io_in = _T_1239 & io_rPort_11_en_0; // @[package.scala 94:16:@9746.4]
  assign RetimeWrapper_47_clock = clock; // @[:@9752.4]
  assign RetimeWrapper_47_reset = reset; // @[:@9753.4]
  assign RetimeWrapper_47_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@9755.4]
  assign RetimeWrapper_47_io_in = _T_1409 & io_rPort_11_en_0; // @[package.scala 94:16:@9754.4]
  assign RetimeWrapper_48_clock = clock; // @[:@9776.4]
  assign RetimeWrapper_48_reset = reset; // @[:@9777.4]
  assign RetimeWrapper_48_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9779.4]
  assign RetimeWrapper_48_io_in = _T_860 & io_rPort_12_en_0; // @[package.scala 94:16:@9778.4]
  assign RetimeWrapper_49_clock = clock; // @[:@9784.4]
  assign RetimeWrapper_49_reset = reset; // @[:@9785.4]
  assign RetimeWrapper_49_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9787.4]
  assign RetimeWrapper_49_io_in = _T_1030 & io_rPort_12_en_0; // @[package.scala 94:16:@9786.4]
  assign RetimeWrapper_50_clock = clock; // @[:@9792.4]
  assign RetimeWrapper_50_reset = reset; // @[:@9793.4]
  assign RetimeWrapper_50_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9795.4]
  assign RetimeWrapper_50_io_in = _T_1200 & io_rPort_12_en_0; // @[package.scala 94:16:@9794.4]
  assign RetimeWrapper_51_clock = clock; // @[:@9800.4]
  assign RetimeWrapper_51_reset = reset; // @[:@9801.4]
  assign RetimeWrapper_51_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@9803.4]
  assign RetimeWrapper_51_io_in = _T_1370 & io_rPort_12_en_0; // @[package.scala 94:16:@9802.4]
  assign RetimeWrapper_52_clock = clock; // @[:@9824.4]
  assign RetimeWrapper_52_reset = reset; // @[:@9825.4]
  assign RetimeWrapper_52_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9827.4]
  assign RetimeWrapper_52_io_in = _T_865 & io_rPort_13_en_0; // @[package.scala 94:16:@9826.4]
  assign RetimeWrapper_53_clock = clock; // @[:@9832.4]
  assign RetimeWrapper_53_reset = reset; // @[:@9833.4]
  assign RetimeWrapper_53_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9835.4]
  assign RetimeWrapper_53_io_in = _T_1035 & io_rPort_13_en_0; // @[package.scala 94:16:@9834.4]
  assign RetimeWrapper_54_clock = clock; // @[:@9840.4]
  assign RetimeWrapper_54_reset = reset; // @[:@9841.4]
  assign RetimeWrapper_54_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9843.4]
  assign RetimeWrapper_54_io_in = _T_1205 & io_rPort_13_en_0; // @[package.scala 94:16:@9842.4]
  assign RetimeWrapper_55_clock = clock; // @[:@9848.4]
  assign RetimeWrapper_55_reset = reset; // @[:@9849.4]
  assign RetimeWrapper_55_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@9851.4]
  assign RetimeWrapper_55_io_in = _T_1375 & io_rPort_13_en_0; // @[package.scala 94:16:@9850.4]
  assign RetimeWrapper_56_clock = clock; // @[:@9872.4]
  assign RetimeWrapper_56_reset = reset; // @[:@9873.4]
  assign RetimeWrapper_56_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9875.4]
  assign RetimeWrapper_56_io_in = _T_994 & io_rPort_14_en_0; // @[package.scala 94:16:@9874.4]
  assign RetimeWrapper_57_clock = clock; // @[:@9880.4]
  assign RetimeWrapper_57_reset = reset; // @[:@9881.4]
  assign RetimeWrapper_57_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9883.4]
  assign RetimeWrapper_57_io_in = _T_1164 & io_rPort_14_en_0; // @[package.scala 94:16:@9882.4]
  assign RetimeWrapper_58_clock = clock; // @[:@9888.4]
  assign RetimeWrapper_58_reset = reset; // @[:@9889.4]
  assign RetimeWrapper_58_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9891.4]
  assign RetimeWrapper_58_io_in = _T_1334 & io_rPort_14_en_0; // @[package.scala 94:16:@9890.4]
  assign RetimeWrapper_59_clock = clock; // @[:@9896.4]
  assign RetimeWrapper_59_reset = reset; // @[:@9897.4]
  assign RetimeWrapper_59_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@9899.4]
  assign RetimeWrapper_59_io_in = _T_1504 & io_rPort_14_en_0; // @[package.scala 94:16:@9898.4]
  assign RetimeWrapper_60_clock = clock; // @[:@9920.4]
  assign RetimeWrapper_60_reset = reset; // @[:@9921.4]
  assign RetimeWrapper_60_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9923.4]
  assign RetimeWrapper_60_io_in = _T_999 & io_rPort_15_en_0; // @[package.scala 94:16:@9922.4]
  assign RetimeWrapper_61_clock = clock; // @[:@9928.4]
  assign RetimeWrapper_61_reset = reset; // @[:@9929.4]
  assign RetimeWrapper_61_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9931.4]
  assign RetimeWrapper_61_io_in = _T_1169 & io_rPort_15_en_0; // @[package.scala 94:16:@9930.4]
  assign RetimeWrapper_62_clock = clock; // @[:@9936.4]
  assign RetimeWrapper_62_reset = reset; // @[:@9937.4]
  assign RetimeWrapper_62_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9939.4]
  assign RetimeWrapper_62_io_in = _T_1339 & io_rPort_15_en_0; // @[package.scala 94:16:@9938.4]
  assign RetimeWrapper_63_clock = clock; // @[:@9944.4]
  assign RetimeWrapper_63_reset = reset; // @[:@9945.4]
  assign RetimeWrapper_63_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@9947.4]
  assign RetimeWrapper_63_io_in = _T_1509 & io_rPort_15_en_0; // @[package.scala 94:16:@9946.4]
  assign RetimeWrapper_64_clock = clock; // @[:@9968.4]
  assign RetimeWrapper_64_reset = reset; // @[:@9969.4]
  assign RetimeWrapper_64_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9971.4]
  assign RetimeWrapper_64_io_in = _T_870 & io_rPort_16_en_0; // @[package.scala 94:16:@9970.4]
  assign RetimeWrapper_65_clock = clock; // @[:@9976.4]
  assign RetimeWrapper_65_reset = reset; // @[:@9977.4]
  assign RetimeWrapper_65_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9979.4]
  assign RetimeWrapper_65_io_in = _T_1040 & io_rPort_16_en_0; // @[package.scala 94:16:@9978.4]
  assign RetimeWrapper_66_clock = clock; // @[:@9984.4]
  assign RetimeWrapper_66_reset = reset; // @[:@9985.4]
  assign RetimeWrapper_66_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9987.4]
  assign RetimeWrapper_66_io_in = _T_1210 & io_rPort_16_en_0; // @[package.scala 94:16:@9986.4]
  assign RetimeWrapper_67_clock = clock; // @[:@9992.4]
  assign RetimeWrapper_67_reset = reset; // @[:@9993.4]
  assign RetimeWrapper_67_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@9995.4]
  assign RetimeWrapper_67_io_in = _T_1380 & io_rPort_16_en_0; // @[package.scala 94:16:@9994.4]
  assign RetimeWrapper_68_clock = clock; // @[:@10016.4]
  assign RetimeWrapper_68_reset = reset; // @[:@10017.4]
  assign RetimeWrapper_68_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10019.4]
  assign RetimeWrapper_68_io_in = _T_943 & io_rPort_17_en_0; // @[package.scala 94:16:@10018.4]
  assign RetimeWrapper_69_clock = clock; // @[:@10024.4]
  assign RetimeWrapper_69_reset = reset; // @[:@10025.4]
  assign RetimeWrapper_69_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10027.4]
  assign RetimeWrapper_69_io_in = _T_1113 & io_rPort_17_en_0; // @[package.scala 94:16:@10026.4]
  assign RetimeWrapper_70_clock = clock; // @[:@10032.4]
  assign RetimeWrapper_70_reset = reset; // @[:@10033.4]
  assign RetimeWrapper_70_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10035.4]
  assign RetimeWrapper_70_io_in = _T_1283 & io_rPort_17_en_0; // @[package.scala 94:16:@10034.4]
  assign RetimeWrapper_71_clock = clock; // @[:@10040.4]
  assign RetimeWrapper_71_reset = reset; // @[:@10041.4]
  assign RetimeWrapper_71_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@10043.4]
  assign RetimeWrapper_71_io_in = _T_1453 & io_rPort_17_en_0; // @[package.scala 94:16:@10042.4]
endmodule
module StickySelects_16( // @[:@11571.2]
  input   clock, // @[:@11572.4]
  input   reset, // @[:@11573.4]
  input   io_ins_0, // @[:@11574.4]
  input   io_ins_1, // @[:@11574.4]
  output  io_outs_0, // @[:@11574.4]
  output  io_outs_1 // @[:@11574.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@11576.4]
  reg [31:0] _RAND_0;
  wire  _T_21; // @[StickySelects.scala 24:52:@11577.4]
  wire  _T_22; // @[StickySelects.scala 24:21:@11578.4]
  reg  _T_25; // @[StickySelects.scala 21:22:@11580.4]
  reg [31:0] _RAND_1;
  wire  _T_27; // @[StickySelects.scala 24:52:@11581.4]
  wire  _T_28; // @[StickySelects.scala 24:21:@11582.4]
  assign _T_21 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@11577.4]
  assign _T_22 = io_ins_1 ? 1'h0 : _T_21; // @[StickySelects.scala 24:21:@11578.4]
  assign _T_27 = io_ins_1 | _T_25; // @[StickySelects.scala 24:52:@11581.4]
  assign _T_28 = io_ins_0 ? 1'h0 : _T_27; // @[StickySelects.scala 24:21:@11582.4]
  assign io_outs_0 = io_ins_1 ? 1'h0 : _T_21; // @[StickySelects.scala 28:52:@11584.4]
  assign io_outs_1 = io_ins_0 ? 1'h0 : _T_27; // @[StickySelects.scala 28:52:@11585.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_25 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_ins_1) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_21;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (io_ins_0) begin
        _T_25 <= 1'h0;
      end else begin
        _T_25 <= _T_27;
      end
    end
  end
endmodule
module StickySelects_19( // @[:@11619.2]
  input   clock, // @[:@11620.4]
  input   reset, // @[:@11621.4]
  input   io_ins_0, // @[:@11622.4]
  input   io_ins_1, // @[:@11622.4]
  input   io_ins_2, // @[:@11622.4]
  input   io_ins_3, // @[:@11622.4]
  output  io_outs_0, // @[:@11622.4]
  output  io_outs_1, // @[:@11622.4]
  output  io_outs_2, // @[:@11622.4]
  output  io_outs_3 // @[:@11622.4]
);
  reg  _T_19; // @[StickySelects.scala 21:22:@11624.4]
  reg [31:0] _RAND_0;
  wire  _T_20; // @[StickySelects.scala 22:54:@11625.4]
  wire  _T_21; // @[StickySelects.scala 22:54:@11626.4]
  wire  _T_23; // @[StickySelects.scala 24:52:@11627.4]
  wire  _T_24; // @[StickySelects.scala 24:21:@11628.4]
  reg  _T_27; // @[StickySelects.scala 21:22:@11630.4]
  reg [31:0] _RAND_1;
  wire  _T_28; // @[StickySelects.scala 22:54:@11631.4]
  wire  _T_29; // @[StickySelects.scala 22:54:@11632.4]
  wire  _T_31; // @[StickySelects.scala 24:52:@11633.4]
  wire  _T_32; // @[StickySelects.scala 24:21:@11634.4]
  reg  _T_35; // @[StickySelects.scala 21:22:@11636.4]
  reg [31:0] _RAND_2;
  wire  _T_36; // @[StickySelects.scala 22:54:@11637.4]
  wire  _T_37; // @[StickySelects.scala 22:54:@11638.4]
  wire  _T_39; // @[StickySelects.scala 24:52:@11639.4]
  wire  _T_40; // @[StickySelects.scala 24:21:@11640.4]
  reg  _T_43; // @[StickySelects.scala 21:22:@11642.4]
  reg [31:0] _RAND_3;
  wire  _T_45; // @[StickySelects.scala 22:54:@11644.4]
  wire  _T_47; // @[StickySelects.scala 24:52:@11645.4]
  wire  _T_48; // @[StickySelects.scala 24:21:@11646.4]
  assign _T_20 = io_ins_1 | io_ins_2; // @[StickySelects.scala 22:54:@11625.4]
  assign _T_21 = _T_20 | io_ins_3; // @[StickySelects.scala 22:54:@11626.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 24:52:@11627.4]
  assign _T_24 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 24:21:@11628.4]
  assign _T_28 = io_ins_0 | io_ins_2; // @[StickySelects.scala 22:54:@11631.4]
  assign _T_29 = _T_28 | io_ins_3; // @[StickySelects.scala 22:54:@11632.4]
  assign _T_31 = io_ins_1 | _T_27; // @[StickySelects.scala 24:52:@11633.4]
  assign _T_32 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 24:21:@11634.4]
  assign _T_36 = io_ins_0 | io_ins_1; // @[StickySelects.scala 22:54:@11637.4]
  assign _T_37 = _T_36 | io_ins_3; // @[StickySelects.scala 22:54:@11638.4]
  assign _T_39 = io_ins_2 | _T_35; // @[StickySelects.scala 24:52:@11639.4]
  assign _T_40 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 24:21:@11640.4]
  assign _T_45 = _T_36 | io_ins_2; // @[StickySelects.scala 22:54:@11644.4]
  assign _T_47 = io_ins_3 | _T_43; // @[StickySelects.scala 24:52:@11645.4]
  assign _T_48 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 24:21:@11646.4]
  assign io_outs_0 = _T_21 ? 1'h0 : _T_23; // @[StickySelects.scala 28:52:@11648.4]
  assign io_outs_1 = _T_29 ? 1'h0 : _T_31; // @[StickySelects.scala 28:52:@11649.4]
  assign io_outs_2 = _T_37 ? 1'h0 : _T_39; // @[StickySelects.scala 28:52:@11650.4]
  assign io_outs_3 = _T_45 ? 1'h0 : _T_47; // @[StickySelects.scala 28:52:@11651.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_27 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_35 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_43 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_21) begin
        _T_19 <= 1'h0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_27 <= 1'h0;
    end else begin
      if (_T_29) begin
        _T_27 <= 1'h0;
      end else begin
        _T_27 <= _T_31;
      end
    end
    if (reset) begin
      _T_35 <= 1'h0;
    end else begin
      if (_T_37) begin
        _T_35 <= 1'h0;
      end else begin
        _T_35 <= _T_39;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_45) begin
        _T_43 <= 1'h0;
      end else begin
        _T_43 <= _T_47;
      end
    end
  end
endmodule
module x387_lb2_0( // @[:@13179.2]
  input        clock, // @[:@13180.4]
  input        reset, // @[:@13181.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@13182.4]
  input        io_rPort_9_ofs_0, // @[:@13182.4]
  input        io_rPort_9_en_0, // @[:@13182.4]
  input        io_rPort_9_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_9_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@13182.4]
  input        io_rPort_8_ofs_0, // @[:@13182.4]
  input        io_rPort_8_en_0, // @[:@13182.4]
  input        io_rPort_8_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_8_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@13182.4]
  input        io_rPort_7_ofs_0, // @[:@13182.4]
  input        io_rPort_7_en_0, // @[:@13182.4]
  input        io_rPort_7_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_7_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@13182.4]
  input        io_rPort_6_ofs_0, // @[:@13182.4]
  input        io_rPort_6_en_0, // @[:@13182.4]
  input        io_rPort_6_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_6_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@13182.4]
  input        io_rPort_5_ofs_0, // @[:@13182.4]
  input        io_rPort_5_en_0, // @[:@13182.4]
  input        io_rPort_5_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_5_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@13182.4]
  input        io_rPort_4_ofs_0, // @[:@13182.4]
  input        io_rPort_4_en_0, // @[:@13182.4]
  input        io_rPort_4_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_4_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@13182.4]
  input        io_rPort_3_ofs_0, // @[:@13182.4]
  input        io_rPort_3_en_0, // @[:@13182.4]
  input        io_rPort_3_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_3_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@13182.4]
  input        io_rPort_2_ofs_0, // @[:@13182.4]
  input        io_rPort_2_en_0, // @[:@13182.4]
  input        io_rPort_2_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_2_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@13182.4]
  input        io_rPort_1_ofs_0, // @[:@13182.4]
  input        io_rPort_1_en_0, // @[:@13182.4]
  input        io_rPort_1_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_1_output_0, // @[:@13182.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@13182.4]
  input        io_rPort_0_ofs_0, // @[:@13182.4]
  input        io_rPort_0_en_0, // @[:@13182.4]
  input        io_rPort_0_backpressure, // @[:@13182.4]
  output [7:0] io_rPort_0_output_0, // @[:@13182.4]
  input  [2:0] io_wPort_3_banks_0, // @[:@13182.4]
  input        io_wPort_3_ofs_0, // @[:@13182.4]
  input  [7:0] io_wPort_3_data_0, // @[:@13182.4]
  input        io_wPort_3_en_0, // @[:@13182.4]
  input  [2:0] io_wPort_2_banks_0, // @[:@13182.4]
  input        io_wPort_2_ofs_0, // @[:@13182.4]
  input  [7:0] io_wPort_2_data_0, // @[:@13182.4]
  input        io_wPort_2_en_0, // @[:@13182.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@13182.4]
  input        io_wPort_1_ofs_0, // @[:@13182.4]
  input  [7:0] io_wPort_1_data_0, // @[:@13182.4]
  input        io_wPort_1_en_0, // @[:@13182.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@13182.4]
  input        io_wPort_0_ofs_0, // @[:@13182.4]
  input  [7:0] io_wPort_0_data_0, // @[:@13182.4]
  input        io_wPort_0_en_0 // @[:@13182.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@13277.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@13277.4]
  wire  Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13277.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13277.4]
  wire  Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13277.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@13277.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@13277.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@13277.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@13293.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@13293.4]
  wire  Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13293.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13293.4]
  wire  Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13293.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@13293.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@13293.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@13293.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@13309.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@13309.4]
  wire  Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13309.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13309.4]
  wire  Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13309.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@13309.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@13309.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@13309.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@13325.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@13325.4]
  wire  Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13325.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13325.4]
  wire  Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13325.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@13325.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@13325.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@13325.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@13341.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@13341.4]
  wire  Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13341.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13341.4]
  wire  Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13341.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@13341.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@13341.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@13341.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@13357.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@13357.4]
  wire  Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13357.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13357.4]
  wire  Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13357.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@13357.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@13357.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@13357.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@13373.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@13373.4]
  wire  Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13373.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13373.4]
  wire  Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13373.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@13373.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@13373.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@13373.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@13389.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@13389.4]
  wire  Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13389.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13389.4]
  wire  Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13389.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@13389.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@13389.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@13389.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@13405.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@13405.4]
  wire  Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13405.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13405.4]
  wire  Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13405.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@13405.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@13405.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@13405.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@13421.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@13421.4]
  wire  Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13421.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13421.4]
  wire  Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13421.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@13421.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@13421.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@13421.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@13437.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@13437.4]
  wire  Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13437.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13437.4]
  wire  Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13437.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@13437.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@13437.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@13437.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@13453.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@13453.4]
  wire  Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13453.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13453.4]
  wire  Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13453.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@13453.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@13453.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@13453.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@13469.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@13469.4]
  wire  Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13469.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13469.4]
  wire  Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13469.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@13469.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@13469.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@13469.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@13485.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@13485.4]
  wire  Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13485.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13485.4]
  wire  Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13485.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@13485.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@13485.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@13485.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@13501.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@13501.4]
  wire  Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13501.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13501.4]
  wire  Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13501.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@13501.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@13501.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@13501.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@13517.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@13517.4]
  wire  Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13517.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13517.4]
  wire  Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13517.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@13517.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@13517.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@13517.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@13739.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@13739.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@13739.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@13739.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@13739.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@13739.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@13763.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@13763.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@13763.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@13763.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@13763.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@13763.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@13793.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@13827.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@13827.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@13827.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@13827.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@13827.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@13827.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@13851.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@13851.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@13851.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@13851.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@13851.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@13851.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@13875.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@13875.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@13875.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@13875.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@13875.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@13875.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@13905.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@13939.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@13939.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@13939.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@13939.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@13939.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@13939.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@13987.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@13987.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@13987.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@13987.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@13987.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@13987.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@14017.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@14051.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@14051.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@14051.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@14051.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@14051.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@14051.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@14075.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@14075.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@14075.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@14075.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@14075.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@14075.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@14099.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@14099.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@14099.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@14099.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@14099.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@14099.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@14129.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14170.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14170.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14170.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14170.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14170.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14178.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14178.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14178.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14178.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14178.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14186.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14186.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14186.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14186.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14186.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14194.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14194.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14194.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14194.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14194.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14218.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14218.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14218.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14218.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14218.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14226.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14226.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14226.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14226.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14226.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14234.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14234.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14234.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14234.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14234.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14242.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14242.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14242.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14242.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14242.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14266.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14266.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14266.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14266.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14266.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14274.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14274.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14274.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14274.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14274.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14282.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14282.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14282.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14282.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14282.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14290.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14290.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14290.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14290.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14290.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14314.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14314.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14314.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14314.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14314.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14322.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14322.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14322.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14322.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14322.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14330.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14330.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14330.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14330.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14330.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14338.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14338.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14338.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14338.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14338.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14362.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14362.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14362.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14362.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14362.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14370.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14370.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14370.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14370.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14370.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14378.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14378.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14378.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14378.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14378.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14386.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14386.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14386.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14386.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14386.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14410.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14410.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14410.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14410.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14410.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14418.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14418.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14418.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14418.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14418.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14426.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14426.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14426.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14426.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14426.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14434.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14434.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14434.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14434.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14434.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14458.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14458.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14458.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14458.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14458.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14466.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14466.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14466.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14466.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14466.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14474.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14474.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14474.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14474.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14474.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14482.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14482.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14482.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14482.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14482.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14506.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14506.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14506.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14506.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14506.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14514.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14514.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14514.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14514.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14514.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14522.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14522.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14522.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14522.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14522.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14530.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14530.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14530.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14530.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14530.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14554.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14554.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14554.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14554.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14554.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14562.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14562.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14562.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14562.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14562.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14570.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14570.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14570.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14570.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14570.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14578.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14578.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14578.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14578.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14578.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14602.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14602.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14602.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14602.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14602.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14610.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14610.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14610.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14610.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14610.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14618.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14618.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14618.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14618.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14618.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14626.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14626.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14626.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14626.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14626.4]
  wire  _T_460; // @[MemPrimitives.scala 82:210:@13533.4]
  wire  _T_463; // @[MemPrimitives.scala 83:102:@13535.4]
  wire [9:0] _T_465; // @[Cat.scala 30:58:@13537.4]
  wire  _T_470; // @[MemPrimitives.scala 82:210:@13544.4]
  wire  _T_473; // @[MemPrimitives.scala 83:102:@13546.4]
  wire [9:0] _T_475; // @[Cat.scala 30:58:@13548.4]
  wire  _T_480; // @[MemPrimitives.scala 82:210:@13555.4]
  wire  _T_483; // @[MemPrimitives.scala 83:102:@13557.4]
  wire [9:0] _T_485; // @[Cat.scala 30:58:@13559.4]
  wire  _T_490; // @[MemPrimitives.scala 82:210:@13566.4]
  wire  _T_493; // @[MemPrimitives.scala 83:102:@13568.4]
  wire [9:0] _T_495; // @[Cat.scala 30:58:@13570.4]
  wire  _T_500; // @[MemPrimitives.scala 82:210:@13577.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@13579.4]
  wire [9:0] _T_505; // @[Cat.scala 30:58:@13581.4]
  wire  _T_510; // @[MemPrimitives.scala 82:210:@13588.4]
  wire  _T_513; // @[MemPrimitives.scala 83:102:@13590.4]
  wire [9:0] _T_515; // @[Cat.scala 30:58:@13592.4]
  wire  _T_520; // @[MemPrimitives.scala 82:210:@13599.4]
  wire  _T_523; // @[MemPrimitives.scala 83:102:@13601.4]
  wire [9:0] _T_525; // @[Cat.scala 30:58:@13603.4]
  wire  _T_530; // @[MemPrimitives.scala 82:210:@13610.4]
  wire  _T_533; // @[MemPrimitives.scala 83:102:@13612.4]
  wire [9:0] _T_535; // @[Cat.scala 30:58:@13614.4]
  wire  _T_540; // @[MemPrimitives.scala 82:210:@13621.4]
  wire  _T_543; // @[MemPrimitives.scala 83:102:@13623.4]
  wire [9:0] _T_545; // @[Cat.scala 30:58:@13625.4]
  wire  _T_550; // @[MemPrimitives.scala 82:210:@13632.4]
  wire  _T_553; // @[MemPrimitives.scala 83:102:@13634.4]
  wire [9:0] _T_555; // @[Cat.scala 30:58:@13636.4]
  wire  _T_560; // @[MemPrimitives.scala 82:210:@13643.4]
  wire  _T_563; // @[MemPrimitives.scala 83:102:@13645.4]
  wire [9:0] _T_565; // @[Cat.scala 30:58:@13647.4]
  wire  _T_570; // @[MemPrimitives.scala 82:210:@13654.4]
  wire  _T_573; // @[MemPrimitives.scala 83:102:@13656.4]
  wire [9:0] _T_575; // @[Cat.scala 30:58:@13658.4]
  wire  _T_580; // @[MemPrimitives.scala 82:210:@13665.4]
  wire  _T_583; // @[MemPrimitives.scala 83:102:@13667.4]
  wire [9:0] _T_585; // @[Cat.scala 30:58:@13669.4]
  wire  _T_590; // @[MemPrimitives.scala 82:210:@13676.4]
  wire  _T_593; // @[MemPrimitives.scala 83:102:@13678.4]
  wire [9:0] _T_595; // @[Cat.scala 30:58:@13680.4]
  wire  _T_600; // @[MemPrimitives.scala 82:210:@13687.4]
  wire  _T_603; // @[MemPrimitives.scala 83:102:@13689.4]
  wire [9:0] _T_605; // @[Cat.scala 30:58:@13691.4]
  wire  _T_610; // @[MemPrimitives.scala 82:210:@13698.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@13700.4]
  wire [9:0] _T_615; // @[Cat.scala 30:58:@13702.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@13709.4]
  wire  _T_625; // @[MemPrimitives.scala 110:210:@13712.4]
  wire  _T_629; // @[MemPrimitives.scala 123:41:@13720.4]
  wire  _T_630; // @[MemPrimitives.scala 123:41:@13721.4]
  wire [2:0] _T_632; // @[Cat.scala 30:58:@13723.4]
  wire [2:0] _T_634; // @[Cat.scala 30:58:@13725.4]
  wire [2:0] _T_635; // @[Mux.scala 31:69:@13726.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13733.4]
  wire  _T_645; // @[MemPrimitives.scala 110:210:@13736.4]
  wire  _T_649; // @[MemPrimitives.scala 123:41:@13744.4]
  wire  _T_650; // @[MemPrimitives.scala 123:41:@13745.4]
  wire [2:0] _T_652; // @[Cat.scala 30:58:@13747.4]
  wire [2:0] _T_654; // @[Cat.scala 30:58:@13749.4]
  wire [2:0] _T_655; // @[Mux.scala 31:69:@13750.4]
  wire  _T_660; // @[MemPrimitives.scala 110:210:@13757.4]
  wire  _T_665; // @[MemPrimitives.scala 110:210:@13760.4]
  wire  _T_669; // @[MemPrimitives.scala 123:41:@13768.4]
  wire  _T_670; // @[MemPrimitives.scala 123:41:@13769.4]
  wire [2:0] _T_672; // @[Cat.scala 30:58:@13771.4]
  wire [2:0] _T_674; // @[Cat.scala 30:58:@13773.4]
  wire [2:0] _T_675; // @[Mux.scala 31:69:@13774.4]
  wire  _T_680; // @[MemPrimitives.scala 110:210:@13781.4]
  wire  _T_685; // @[MemPrimitives.scala 110:210:@13784.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@13787.4]
  wire  _T_695; // @[MemPrimitives.scala 110:210:@13790.4]
  wire  _T_699; // @[MemPrimitives.scala 123:41:@13800.4]
  wire  _T_700; // @[MemPrimitives.scala 123:41:@13801.4]
  wire  _T_701; // @[MemPrimitives.scala 123:41:@13802.4]
  wire  _T_702; // @[MemPrimitives.scala 123:41:@13803.4]
  wire [2:0] _T_704; // @[Cat.scala 30:58:@13805.4]
  wire [2:0] _T_706; // @[Cat.scala 30:58:@13807.4]
  wire [2:0] _T_708; // @[Cat.scala 30:58:@13809.4]
  wire [2:0] _T_710; // @[Cat.scala 30:58:@13811.4]
  wire [2:0] _T_711; // @[Mux.scala 31:69:@13812.4]
  wire [2:0] _T_712; // @[Mux.scala 31:69:@13813.4]
  wire [2:0] _T_713; // @[Mux.scala 31:69:@13814.4]
  wire  _T_718; // @[MemPrimitives.scala 110:210:@13821.4]
  wire  _T_723; // @[MemPrimitives.scala 110:210:@13824.4]
  wire  _T_727; // @[MemPrimitives.scala 123:41:@13832.4]
  wire  _T_728; // @[MemPrimitives.scala 123:41:@13833.4]
  wire [2:0] _T_730; // @[Cat.scala 30:58:@13835.4]
  wire [2:0] _T_732; // @[Cat.scala 30:58:@13837.4]
  wire [2:0] _T_733; // @[Mux.scala 31:69:@13838.4]
  wire  _T_738; // @[MemPrimitives.scala 110:210:@13845.4]
  wire  _T_743; // @[MemPrimitives.scala 110:210:@13848.4]
  wire  _T_747; // @[MemPrimitives.scala 123:41:@13856.4]
  wire  _T_748; // @[MemPrimitives.scala 123:41:@13857.4]
  wire [2:0] _T_750; // @[Cat.scala 30:58:@13859.4]
  wire [2:0] _T_752; // @[Cat.scala 30:58:@13861.4]
  wire [2:0] _T_753; // @[Mux.scala 31:69:@13862.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@13869.4]
  wire  _T_763; // @[MemPrimitives.scala 110:210:@13872.4]
  wire  _T_767; // @[MemPrimitives.scala 123:41:@13880.4]
  wire  _T_768; // @[MemPrimitives.scala 123:41:@13881.4]
  wire [2:0] _T_770; // @[Cat.scala 30:58:@13883.4]
  wire [2:0] _T_772; // @[Cat.scala 30:58:@13885.4]
  wire [2:0] _T_773; // @[Mux.scala 31:69:@13886.4]
  wire  _T_778; // @[MemPrimitives.scala 110:210:@13893.4]
  wire  _T_783; // @[MemPrimitives.scala 110:210:@13896.4]
  wire  _T_788; // @[MemPrimitives.scala 110:210:@13899.4]
  wire  _T_793; // @[MemPrimitives.scala 110:210:@13902.4]
  wire  _T_797; // @[MemPrimitives.scala 123:41:@13912.4]
  wire  _T_798; // @[MemPrimitives.scala 123:41:@13913.4]
  wire  _T_799; // @[MemPrimitives.scala 123:41:@13914.4]
  wire  _T_800; // @[MemPrimitives.scala 123:41:@13915.4]
  wire [2:0] _T_802; // @[Cat.scala 30:58:@13917.4]
  wire [2:0] _T_804; // @[Cat.scala 30:58:@13919.4]
  wire [2:0] _T_806; // @[Cat.scala 30:58:@13921.4]
  wire [2:0] _T_808; // @[Cat.scala 30:58:@13923.4]
  wire [2:0] _T_809; // @[Mux.scala 31:69:@13924.4]
  wire [2:0] _T_810; // @[Mux.scala 31:69:@13925.4]
  wire [2:0] _T_811; // @[Mux.scala 31:69:@13926.4]
  wire  _T_816; // @[MemPrimitives.scala 110:210:@13933.4]
  wire  _T_821; // @[MemPrimitives.scala 110:210:@13936.4]
  wire  _T_825; // @[MemPrimitives.scala 123:41:@13944.4]
  wire  _T_826; // @[MemPrimitives.scala 123:41:@13945.4]
  wire [2:0] _T_828; // @[Cat.scala 30:58:@13947.4]
  wire [2:0] _T_830; // @[Cat.scala 30:58:@13949.4]
  wire [2:0] _T_831; // @[Mux.scala 31:69:@13950.4]
  wire  _T_836; // @[MemPrimitives.scala 110:210:@13957.4]
  wire  _T_841; // @[MemPrimitives.scala 110:210:@13960.4]
  wire  _T_845; // @[MemPrimitives.scala 123:41:@13968.4]
  wire  _T_846; // @[MemPrimitives.scala 123:41:@13969.4]
  wire [2:0] _T_848; // @[Cat.scala 30:58:@13971.4]
  wire [2:0] _T_850; // @[Cat.scala 30:58:@13973.4]
  wire [2:0] _T_851; // @[Mux.scala 31:69:@13974.4]
  wire  _T_856; // @[MemPrimitives.scala 110:210:@13981.4]
  wire  _T_861; // @[MemPrimitives.scala 110:210:@13984.4]
  wire  _T_865; // @[MemPrimitives.scala 123:41:@13992.4]
  wire  _T_866; // @[MemPrimitives.scala 123:41:@13993.4]
  wire [2:0] _T_868; // @[Cat.scala 30:58:@13995.4]
  wire [2:0] _T_870; // @[Cat.scala 30:58:@13997.4]
  wire [2:0] _T_871; // @[Mux.scala 31:69:@13998.4]
  wire  _T_876; // @[MemPrimitives.scala 110:210:@14005.4]
  wire  _T_881; // @[MemPrimitives.scala 110:210:@14008.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@14011.4]
  wire  _T_891; // @[MemPrimitives.scala 110:210:@14014.4]
  wire  _T_895; // @[MemPrimitives.scala 123:41:@14024.4]
  wire  _T_896; // @[MemPrimitives.scala 123:41:@14025.4]
  wire  _T_897; // @[MemPrimitives.scala 123:41:@14026.4]
  wire  _T_898; // @[MemPrimitives.scala 123:41:@14027.4]
  wire [2:0] _T_900; // @[Cat.scala 30:58:@14029.4]
  wire [2:0] _T_902; // @[Cat.scala 30:58:@14031.4]
  wire [2:0] _T_904; // @[Cat.scala 30:58:@14033.4]
  wire [2:0] _T_906; // @[Cat.scala 30:58:@14035.4]
  wire [2:0] _T_907; // @[Mux.scala 31:69:@14036.4]
  wire [2:0] _T_908; // @[Mux.scala 31:69:@14037.4]
  wire [2:0] _T_909; // @[Mux.scala 31:69:@14038.4]
  wire  _T_914; // @[MemPrimitives.scala 110:210:@14045.4]
  wire  _T_919; // @[MemPrimitives.scala 110:210:@14048.4]
  wire  _T_923; // @[MemPrimitives.scala 123:41:@14056.4]
  wire  _T_924; // @[MemPrimitives.scala 123:41:@14057.4]
  wire [2:0] _T_926; // @[Cat.scala 30:58:@14059.4]
  wire [2:0] _T_928; // @[Cat.scala 30:58:@14061.4]
  wire [2:0] _T_929; // @[Mux.scala 31:69:@14062.4]
  wire  _T_934; // @[MemPrimitives.scala 110:210:@14069.4]
  wire  _T_939; // @[MemPrimitives.scala 110:210:@14072.4]
  wire  _T_943; // @[MemPrimitives.scala 123:41:@14080.4]
  wire  _T_944; // @[MemPrimitives.scala 123:41:@14081.4]
  wire [2:0] _T_946; // @[Cat.scala 30:58:@14083.4]
  wire [2:0] _T_948; // @[Cat.scala 30:58:@14085.4]
  wire [2:0] _T_949; // @[Mux.scala 31:69:@14086.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@14093.4]
  wire  _T_959; // @[MemPrimitives.scala 110:210:@14096.4]
  wire  _T_963; // @[MemPrimitives.scala 123:41:@14104.4]
  wire  _T_964; // @[MemPrimitives.scala 123:41:@14105.4]
  wire [2:0] _T_966; // @[Cat.scala 30:58:@14107.4]
  wire [2:0] _T_968; // @[Cat.scala 30:58:@14109.4]
  wire [2:0] _T_969; // @[Mux.scala 31:69:@14110.4]
  wire  _T_974; // @[MemPrimitives.scala 110:210:@14117.4]
  wire  _T_979; // @[MemPrimitives.scala 110:210:@14120.4]
  wire  _T_984; // @[MemPrimitives.scala 110:210:@14123.4]
  wire  _T_989; // @[MemPrimitives.scala 110:210:@14126.4]
  wire  _T_993; // @[MemPrimitives.scala 123:41:@14136.4]
  wire  _T_994; // @[MemPrimitives.scala 123:41:@14137.4]
  wire  _T_995; // @[MemPrimitives.scala 123:41:@14138.4]
  wire  _T_996; // @[MemPrimitives.scala 123:41:@14139.4]
  wire [2:0] _T_998; // @[Cat.scala 30:58:@14141.4]
  wire [2:0] _T_1000; // @[Cat.scala 30:58:@14143.4]
  wire [2:0] _T_1002; // @[Cat.scala 30:58:@14145.4]
  wire [2:0] _T_1004; // @[Cat.scala 30:58:@14147.4]
  wire [2:0] _T_1005; // @[Mux.scala 31:69:@14148.4]
  wire [2:0] _T_1006; // @[Mux.scala 31:69:@14149.4]
  wire [2:0] _T_1007; // @[Mux.scala 31:69:@14150.4]
  wire  _T_1039; // @[package.scala 96:25:@14191.4 package.scala 96:25:@14192.4]
  wire [7:0] _T_1043; // @[Mux.scala 31:69:@14201.4]
  wire  _T_1036; // @[package.scala 96:25:@14183.4 package.scala 96:25:@14184.4]
  wire [7:0] _T_1044; // @[Mux.scala 31:69:@14202.4]
  wire  _T_1033; // @[package.scala 96:25:@14175.4 package.scala 96:25:@14176.4]
  wire  _T_1074; // @[package.scala 96:25:@14239.4 package.scala 96:25:@14240.4]
  wire [7:0] _T_1078; // @[Mux.scala 31:69:@14249.4]
  wire  _T_1071; // @[package.scala 96:25:@14231.4 package.scala 96:25:@14232.4]
  wire [7:0] _T_1079; // @[Mux.scala 31:69:@14250.4]
  wire  _T_1068; // @[package.scala 96:25:@14223.4 package.scala 96:25:@14224.4]
  wire  _T_1109; // @[package.scala 96:25:@14287.4 package.scala 96:25:@14288.4]
  wire [7:0] _T_1113; // @[Mux.scala 31:69:@14297.4]
  wire  _T_1106; // @[package.scala 96:25:@14279.4 package.scala 96:25:@14280.4]
  wire [7:0] _T_1114; // @[Mux.scala 31:69:@14298.4]
  wire  _T_1103; // @[package.scala 96:25:@14271.4 package.scala 96:25:@14272.4]
  wire  _T_1144; // @[package.scala 96:25:@14335.4 package.scala 96:25:@14336.4]
  wire [7:0] _T_1148; // @[Mux.scala 31:69:@14345.4]
  wire  _T_1141; // @[package.scala 96:25:@14327.4 package.scala 96:25:@14328.4]
  wire [7:0] _T_1149; // @[Mux.scala 31:69:@14346.4]
  wire  _T_1138; // @[package.scala 96:25:@14319.4 package.scala 96:25:@14320.4]
  wire  _T_1179; // @[package.scala 96:25:@14383.4 package.scala 96:25:@14384.4]
  wire [7:0] _T_1183; // @[Mux.scala 31:69:@14393.4]
  wire  _T_1176; // @[package.scala 96:25:@14375.4 package.scala 96:25:@14376.4]
  wire [7:0] _T_1184; // @[Mux.scala 31:69:@14394.4]
  wire  _T_1173; // @[package.scala 96:25:@14367.4 package.scala 96:25:@14368.4]
  wire  _T_1214; // @[package.scala 96:25:@14431.4 package.scala 96:25:@14432.4]
  wire [7:0] _T_1218; // @[Mux.scala 31:69:@14441.4]
  wire  _T_1211; // @[package.scala 96:25:@14423.4 package.scala 96:25:@14424.4]
  wire [7:0] _T_1219; // @[Mux.scala 31:69:@14442.4]
  wire  _T_1208; // @[package.scala 96:25:@14415.4 package.scala 96:25:@14416.4]
  wire  _T_1249; // @[package.scala 96:25:@14479.4 package.scala 96:25:@14480.4]
  wire [7:0] _T_1253; // @[Mux.scala 31:69:@14489.4]
  wire  _T_1246; // @[package.scala 96:25:@14471.4 package.scala 96:25:@14472.4]
  wire [7:0] _T_1254; // @[Mux.scala 31:69:@14490.4]
  wire  _T_1243; // @[package.scala 96:25:@14463.4 package.scala 96:25:@14464.4]
  wire  _T_1284; // @[package.scala 96:25:@14527.4 package.scala 96:25:@14528.4]
  wire [7:0] _T_1288; // @[Mux.scala 31:69:@14537.4]
  wire  _T_1281; // @[package.scala 96:25:@14519.4 package.scala 96:25:@14520.4]
  wire [7:0] _T_1289; // @[Mux.scala 31:69:@14538.4]
  wire  _T_1278; // @[package.scala 96:25:@14511.4 package.scala 96:25:@14512.4]
  wire  _T_1319; // @[package.scala 96:25:@14575.4 package.scala 96:25:@14576.4]
  wire [7:0] _T_1323; // @[Mux.scala 31:69:@14585.4]
  wire  _T_1316; // @[package.scala 96:25:@14567.4 package.scala 96:25:@14568.4]
  wire [7:0] _T_1324; // @[Mux.scala 31:69:@14586.4]
  wire  _T_1313; // @[package.scala 96:25:@14559.4 package.scala 96:25:@14560.4]
  wire  _T_1354; // @[package.scala 96:25:@14623.4 package.scala 96:25:@14624.4]
  wire [7:0] _T_1358; // @[Mux.scala 31:69:@14633.4]
  wire  _T_1351; // @[package.scala 96:25:@14615.4 package.scala 96:25:@14616.4]
  wire [7:0] _T_1359; // @[Mux.scala 31:69:@14634.4]
  wire  _T_1348; // @[package.scala 96:25:@14607.4 package.scala 96:25:@14608.4]
  Mem1D_4 Mem1D ( // @[MemPrimitives.scala 64:21:@13277.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_4 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@13293.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_4 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@13309.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_4 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@13325.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_4 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@13341.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_4 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@13357.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_4 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@13373.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_4 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@13389.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_4 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@13405.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_4 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@13421.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_4 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@13437.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_4 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@13453.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_4 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@13469.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_4 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@13485.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_4 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@13501.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_4 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@13517.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_16 StickySelects ( // @[MemPrimitives.scala 121:29:@13715.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1)
  );
  StickySelects_16 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@13739.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1)
  );
  StickySelects_16 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@13763.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1)
  );
  StickySelects_19 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@13793.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3)
  );
  StickySelects_16 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@13827.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1)
  );
  StickySelects_16 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@13851.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1)
  );
  StickySelects_16 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@13875.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1)
  );
  StickySelects_19 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@13905.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3)
  );
  StickySelects_16 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@13939.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1)
  );
  StickySelects_16 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@13963.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1)
  );
  StickySelects_16 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@13987.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1)
  );
  StickySelects_19 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@14017.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3)
  );
  StickySelects_16 StickySelects_12 ( // @[MemPrimitives.scala 121:29:@14051.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1)
  );
  StickySelects_16 StickySelects_13 ( // @[MemPrimitives.scala 121:29:@14075.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1)
  );
  StickySelects_16 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@14099.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1)
  );
  StickySelects_19 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@14129.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@14170.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_1 ( // @[package.scala 93:22:@14178.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_2 ( // @[package.scala 93:22:@14186.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_3 ( // @[package.scala 93:22:@14194.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_4 ( // @[package.scala 93:22:@14218.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_5 ( // @[package.scala 93:22:@14226.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_6 ( // @[package.scala 93:22:@14234.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_7 ( // @[package.scala 93:22:@14242.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_8 ( // @[package.scala 93:22:@14266.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_9 ( // @[package.scala 93:22:@14274.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_10 ( // @[package.scala 93:22:@14282.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_11 ( // @[package.scala 93:22:@14290.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_12 ( // @[package.scala 93:22:@14314.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_13 ( // @[package.scala 93:22:@14322.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_14 ( // @[package.scala 93:22:@14330.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_15 ( // @[package.scala 93:22:@14338.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_16 ( // @[package.scala 93:22:@14362.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_17 ( // @[package.scala 93:22:@14370.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_18 ( // @[package.scala 93:22:@14378.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_19 ( // @[package.scala 93:22:@14386.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_20 ( // @[package.scala 93:22:@14410.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_21 ( // @[package.scala 93:22:@14418.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_22 ( // @[package.scala 93:22:@14426.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_23 ( // @[package.scala 93:22:@14434.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_24 ( // @[package.scala 93:22:@14458.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_25 ( // @[package.scala 93:22:@14466.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_26 ( // @[package.scala 93:22:@14474.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_27 ( // @[package.scala 93:22:@14482.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_28 ( // @[package.scala 93:22:@14506.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_29 ( // @[package.scala 93:22:@14514.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_30 ( // @[package.scala 93:22:@14522.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_31 ( // @[package.scala 93:22:@14530.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_32 ( // @[package.scala 93:22:@14554.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_33 ( // @[package.scala 93:22:@14562.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_34 ( // @[package.scala 93:22:@14570.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_35 ( // @[package.scala 93:22:@14578.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_36 ( // @[package.scala 93:22:@14602.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_37 ( // @[package.scala 93:22:@14610.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@14618.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_39 ( // @[package.scala 93:22:@14626.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  assign _T_460 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13533.4]
  assign _T_463 = io_wPort_0_en_0 & _T_460; // @[MemPrimitives.scala 83:102:@13535.4]
  assign _T_465 = {_T_463,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13537.4]
  assign _T_470 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13544.4]
  assign _T_473 = io_wPort_1_en_0 & _T_470; // @[MemPrimitives.scala 83:102:@13546.4]
  assign _T_475 = {_T_473,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13548.4]
  assign _T_480 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13555.4]
  assign _T_483 = io_wPort_2_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@13557.4]
  assign _T_485 = {_T_483,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@13559.4]
  assign _T_490 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13566.4]
  assign _T_493 = io_wPort_3_en_0 & _T_490; // @[MemPrimitives.scala 83:102:@13568.4]
  assign _T_495 = {_T_493,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@13570.4]
  assign _T_500 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13577.4]
  assign _T_503 = io_wPort_0_en_0 & _T_500; // @[MemPrimitives.scala 83:102:@13579.4]
  assign _T_505 = {_T_503,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13581.4]
  assign _T_510 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13588.4]
  assign _T_513 = io_wPort_1_en_0 & _T_510; // @[MemPrimitives.scala 83:102:@13590.4]
  assign _T_515 = {_T_513,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13592.4]
  assign _T_520 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13599.4]
  assign _T_523 = io_wPort_2_en_0 & _T_520; // @[MemPrimitives.scala 83:102:@13601.4]
  assign _T_525 = {_T_523,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@13603.4]
  assign _T_530 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13610.4]
  assign _T_533 = io_wPort_3_en_0 & _T_530; // @[MemPrimitives.scala 83:102:@13612.4]
  assign _T_535 = {_T_533,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@13614.4]
  assign _T_540 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13621.4]
  assign _T_543 = io_wPort_0_en_0 & _T_540; // @[MemPrimitives.scala 83:102:@13623.4]
  assign _T_545 = {_T_543,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13625.4]
  assign _T_550 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13632.4]
  assign _T_553 = io_wPort_1_en_0 & _T_550; // @[MemPrimitives.scala 83:102:@13634.4]
  assign _T_555 = {_T_553,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13636.4]
  assign _T_560 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13643.4]
  assign _T_563 = io_wPort_2_en_0 & _T_560; // @[MemPrimitives.scala 83:102:@13645.4]
  assign _T_565 = {_T_563,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@13647.4]
  assign _T_570 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13654.4]
  assign _T_573 = io_wPort_3_en_0 & _T_570; // @[MemPrimitives.scala 83:102:@13656.4]
  assign _T_575 = {_T_573,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@13658.4]
  assign _T_580 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13665.4]
  assign _T_583 = io_wPort_0_en_0 & _T_580; // @[MemPrimitives.scala 83:102:@13667.4]
  assign _T_585 = {_T_583,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13669.4]
  assign _T_590 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13676.4]
  assign _T_593 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@13678.4]
  assign _T_595 = {_T_593,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13680.4]
  assign _T_600 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13687.4]
  assign _T_603 = io_wPort_2_en_0 & _T_600; // @[MemPrimitives.scala 83:102:@13689.4]
  assign _T_605 = {_T_603,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@13691.4]
  assign _T_610 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13698.4]
  assign _T_613 = io_wPort_3_en_0 & _T_610; // @[MemPrimitives.scala 83:102:@13700.4]
  assign _T_615 = {_T_613,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@13702.4]
  assign _T_620 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13709.4]
  assign _T_625 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13712.4]
  assign _T_629 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@13720.4]
  assign _T_630 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@13721.4]
  assign _T_632 = {_T_629,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13723.4]
  assign _T_634 = {_T_630,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13725.4]
  assign _T_635 = _T_629 ? _T_632 : _T_634; // @[Mux.scala 31:69:@13726.4]
  assign _T_640 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13733.4]
  assign _T_645 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13736.4]
  assign _T_649 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@13744.4]
  assign _T_650 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@13745.4]
  assign _T_652 = {_T_649,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13747.4]
  assign _T_654 = {_T_650,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13749.4]
  assign _T_655 = _T_649 ? _T_652 : _T_654; // @[Mux.scala 31:69:@13750.4]
  assign _T_660 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13757.4]
  assign _T_665 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13760.4]
  assign _T_669 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@13768.4]
  assign _T_670 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@13769.4]
  assign _T_672 = {_T_669,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13771.4]
  assign _T_674 = {_T_670,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13773.4]
  assign _T_675 = _T_669 ? _T_672 : _T_674; // @[Mux.scala 31:69:@13774.4]
  assign _T_680 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13781.4]
  assign _T_685 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13784.4]
  assign _T_690 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13787.4]
  assign _T_695 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13790.4]
  assign _T_699 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@13800.4]
  assign _T_700 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@13801.4]
  assign _T_701 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@13802.4]
  assign _T_702 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@13803.4]
  assign _T_704 = {_T_699,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13805.4]
  assign _T_706 = {_T_700,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13807.4]
  assign _T_708 = {_T_701,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13809.4]
  assign _T_710 = {_T_702,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13811.4]
  assign _T_711 = _T_701 ? _T_708 : _T_710; // @[Mux.scala 31:69:@13812.4]
  assign _T_712 = _T_700 ? _T_706 : _T_711; // @[Mux.scala 31:69:@13813.4]
  assign _T_713 = _T_699 ? _T_704 : _T_712; // @[Mux.scala 31:69:@13814.4]
  assign _T_718 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13821.4]
  assign _T_723 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13824.4]
  assign _T_727 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@13832.4]
  assign _T_728 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@13833.4]
  assign _T_730 = {_T_727,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13835.4]
  assign _T_732 = {_T_728,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13837.4]
  assign _T_733 = _T_727 ? _T_730 : _T_732; // @[Mux.scala 31:69:@13838.4]
  assign _T_738 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13845.4]
  assign _T_743 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13848.4]
  assign _T_747 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@13856.4]
  assign _T_748 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@13857.4]
  assign _T_750 = {_T_747,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13859.4]
  assign _T_752 = {_T_748,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13861.4]
  assign _T_753 = _T_747 ? _T_750 : _T_752; // @[Mux.scala 31:69:@13862.4]
  assign _T_758 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13869.4]
  assign _T_763 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13872.4]
  assign _T_767 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@13880.4]
  assign _T_768 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@13881.4]
  assign _T_770 = {_T_767,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13883.4]
  assign _T_772 = {_T_768,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13885.4]
  assign _T_773 = _T_767 ? _T_770 : _T_772; // @[Mux.scala 31:69:@13886.4]
  assign _T_778 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13893.4]
  assign _T_783 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13896.4]
  assign _T_788 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13899.4]
  assign _T_793 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13902.4]
  assign _T_797 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@13912.4]
  assign _T_798 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@13913.4]
  assign _T_799 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@13914.4]
  assign _T_800 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@13915.4]
  assign _T_802 = {_T_797,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13917.4]
  assign _T_804 = {_T_798,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13919.4]
  assign _T_806 = {_T_799,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13921.4]
  assign _T_808 = {_T_800,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13923.4]
  assign _T_809 = _T_799 ? _T_806 : _T_808; // @[Mux.scala 31:69:@13924.4]
  assign _T_810 = _T_798 ? _T_804 : _T_809; // @[Mux.scala 31:69:@13925.4]
  assign _T_811 = _T_797 ? _T_802 : _T_810; // @[Mux.scala 31:69:@13926.4]
  assign _T_816 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13933.4]
  assign _T_821 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13936.4]
  assign _T_825 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@13944.4]
  assign _T_826 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@13945.4]
  assign _T_828 = {_T_825,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13947.4]
  assign _T_830 = {_T_826,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13949.4]
  assign _T_831 = _T_825 ? _T_828 : _T_830; // @[Mux.scala 31:69:@13950.4]
  assign _T_836 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13957.4]
  assign _T_841 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13960.4]
  assign _T_845 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@13968.4]
  assign _T_846 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@13969.4]
  assign _T_848 = {_T_845,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13971.4]
  assign _T_850 = {_T_846,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13973.4]
  assign _T_851 = _T_845 ? _T_848 : _T_850; // @[Mux.scala 31:69:@13974.4]
  assign _T_856 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13981.4]
  assign _T_861 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13984.4]
  assign _T_865 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@13992.4]
  assign _T_866 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@13993.4]
  assign _T_868 = {_T_865,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13995.4]
  assign _T_870 = {_T_866,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13997.4]
  assign _T_871 = _T_865 ? _T_868 : _T_870; // @[Mux.scala 31:69:@13998.4]
  assign _T_876 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@14005.4]
  assign _T_881 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@14008.4]
  assign _T_886 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@14011.4]
  assign _T_891 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@14014.4]
  assign _T_895 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@14024.4]
  assign _T_896 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@14025.4]
  assign _T_897 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@14026.4]
  assign _T_898 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@14027.4]
  assign _T_900 = {_T_895,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14029.4]
  assign _T_902 = {_T_896,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14031.4]
  assign _T_904 = {_T_897,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14033.4]
  assign _T_906 = {_T_898,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14035.4]
  assign _T_907 = _T_897 ? _T_904 : _T_906; // @[Mux.scala 31:69:@14036.4]
  assign _T_908 = _T_896 ? _T_902 : _T_907; // @[Mux.scala 31:69:@14037.4]
  assign _T_909 = _T_895 ? _T_900 : _T_908; // @[Mux.scala 31:69:@14038.4]
  assign _T_914 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14045.4]
  assign _T_919 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14048.4]
  assign _T_923 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@14056.4]
  assign _T_924 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@14057.4]
  assign _T_926 = {_T_923,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14059.4]
  assign _T_928 = {_T_924,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14061.4]
  assign _T_929 = _T_923 ? _T_926 : _T_928; // @[Mux.scala 31:69:@14062.4]
  assign _T_934 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14069.4]
  assign _T_939 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14072.4]
  assign _T_943 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@14080.4]
  assign _T_944 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@14081.4]
  assign _T_946 = {_T_943,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14083.4]
  assign _T_948 = {_T_944,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14085.4]
  assign _T_949 = _T_943 ? _T_946 : _T_948; // @[Mux.scala 31:69:@14086.4]
  assign _T_954 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14093.4]
  assign _T_959 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14096.4]
  assign _T_963 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@14104.4]
  assign _T_964 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@14105.4]
  assign _T_966 = {_T_963,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14107.4]
  assign _T_968 = {_T_964,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14109.4]
  assign _T_969 = _T_963 ? _T_966 : _T_968; // @[Mux.scala 31:69:@14110.4]
  assign _T_974 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14117.4]
  assign _T_979 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14120.4]
  assign _T_984 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14123.4]
  assign _T_989 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14126.4]
  assign _T_993 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@14136.4]
  assign _T_994 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@14137.4]
  assign _T_995 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@14138.4]
  assign _T_996 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@14139.4]
  assign _T_998 = {_T_993,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14141.4]
  assign _T_1000 = {_T_994,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14143.4]
  assign _T_1002 = {_T_995,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14145.4]
  assign _T_1004 = {_T_996,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14147.4]
  assign _T_1005 = _T_995 ? _T_1002 : _T_1004; // @[Mux.scala 31:69:@14148.4]
  assign _T_1006 = _T_994 ? _T_1000 : _T_1005; // @[Mux.scala 31:69:@14149.4]
  assign _T_1007 = _T_993 ? _T_998 : _T_1006; // @[Mux.scala 31:69:@14150.4]
  assign _T_1039 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14191.4 package.scala 96:25:@14192.4]
  assign _T_1043 = _T_1039 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@14201.4]
  assign _T_1036 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14183.4 package.scala 96:25:@14184.4]
  assign _T_1044 = _T_1036 ? Mem1D_5_io_output : _T_1043; // @[Mux.scala 31:69:@14202.4]
  assign _T_1033 = RetimeWrapper_io_out; // @[package.scala 96:25:@14175.4 package.scala 96:25:@14176.4]
  assign _T_1074 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14239.4 package.scala 96:25:@14240.4]
  assign _T_1078 = _T_1074 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14249.4]
  assign _T_1071 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14231.4 package.scala 96:25:@14232.4]
  assign _T_1079 = _T_1071 ? Mem1D_7_io_output : _T_1078; // @[Mux.scala 31:69:@14250.4]
  assign _T_1068 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14223.4 package.scala 96:25:@14224.4]
  assign _T_1109 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14287.4 package.scala 96:25:@14288.4]
  assign _T_1113 = _T_1109 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14297.4]
  assign _T_1106 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14279.4 package.scala 96:25:@14280.4]
  assign _T_1114 = _T_1106 ? Mem1D_7_io_output : _T_1113; // @[Mux.scala 31:69:@14298.4]
  assign _T_1103 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14271.4 package.scala 96:25:@14272.4]
  assign _T_1144 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14335.4 package.scala 96:25:@14336.4]
  assign _T_1148 = _T_1144 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14345.4]
  assign _T_1141 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14327.4 package.scala 96:25:@14328.4]
  assign _T_1149 = _T_1141 ? Mem1D_6_io_output : _T_1148; // @[Mux.scala 31:69:@14346.4]
  assign _T_1138 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14319.4 package.scala 96:25:@14320.4]
  assign _T_1179 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14383.4 package.scala 96:25:@14384.4]
  assign _T_1183 = _T_1179 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14393.4]
  assign _T_1176 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14375.4 package.scala 96:25:@14376.4]
  assign _T_1184 = _T_1176 ? Mem1D_7_io_output : _T_1183; // @[Mux.scala 31:69:@14394.4]
  assign _T_1173 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14367.4 package.scala 96:25:@14368.4]
  assign _T_1214 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14431.4 package.scala 96:25:@14432.4]
  assign _T_1218 = _T_1214 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@14441.4]
  assign _T_1211 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14423.4 package.scala 96:25:@14424.4]
  assign _T_1219 = _T_1211 ? Mem1D_4_io_output : _T_1218; // @[Mux.scala 31:69:@14442.4]
  assign _T_1208 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14415.4 package.scala 96:25:@14416.4]
  assign _T_1249 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14479.4 package.scala 96:25:@14480.4]
  assign _T_1253 = _T_1249 ? Mem1D_8_io_output : Mem1D_12_io_output; // @[Mux.scala 31:69:@14489.4]
  assign _T_1246 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14471.4 package.scala 96:25:@14472.4]
  assign _T_1254 = _T_1246 ? Mem1D_4_io_output : _T_1253; // @[Mux.scala 31:69:@14490.4]
  assign _T_1243 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14463.4 package.scala 96:25:@14464.4]
  assign _T_1284 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14527.4 package.scala 96:25:@14528.4]
  assign _T_1288 = _T_1284 ? Mem1D_9_io_output : Mem1D_13_io_output; // @[Mux.scala 31:69:@14537.4]
  assign _T_1281 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14519.4 package.scala 96:25:@14520.4]
  assign _T_1289 = _T_1281 ? Mem1D_5_io_output : _T_1288; // @[Mux.scala 31:69:@14538.4]
  assign _T_1278 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14511.4 package.scala 96:25:@14512.4]
  assign _T_1319 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14575.4 package.scala 96:25:@14576.4]
  assign _T_1323 = _T_1319 ? Mem1D_11_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14585.4]
  assign _T_1316 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14567.4 package.scala 96:25:@14568.4]
  assign _T_1324 = _T_1316 ? Mem1D_7_io_output : _T_1323; // @[Mux.scala 31:69:@14586.4]
  assign _T_1313 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14559.4 package.scala 96:25:@14560.4]
  assign _T_1354 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14623.4 package.scala 96:25:@14624.4]
  assign _T_1358 = _T_1354 ? Mem1D_10_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14633.4]
  assign _T_1351 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14615.4 package.scala 96:25:@14616.4]
  assign _T_1359 = _T_1351 ? Mem1D_6_io_output : _T_1358; // @[Mux.scala 31:69:@14634.4]
  assign _T_1348 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14607.4 package.scala 96:25:@14608.4]
  assign io_rPort_9_output_0 = _T_1348 ? Mem1D_2_io_output : _T_1359; // @[MemPrimitives.scala 148:13:@14636.4]
  assign io_rPort_8_output_0 = _T_1313 ? Mem1D_3_io_output : _T_1324; // @[MemPrimitives.scala 148:13:@14588.4]
  assign io_rPort_7_output_0 = _T_1278 ? Mem1D_1_io_output : _T_1289; // @[MemPrimitives.scala 148:13:@14540.4]
  assign io_rPort_6_output_0 = _T_1243 ? Mem1D_io_output : _T_1254; // @[MemPrimitives.scala 148:13:@14492.4]
  assign io_rPort_5_output_0 = _T_1208 ? Mem1D_io_output : _T_1219; // @[MemPrimitives.scala 148:13:@14444.4]
  assign io_rPort_4_output_0 = _T_1173 ? Mem1D_3_io_output : _T_1184; // @[MemPrimitives.scala 148:13:@14396.4]
  assign io_rPort_3_output_0 = _T_1138 ? Mem1D_2_io_output : _T_1149; // @[MemPrimitives.scala 148:13:@14348.4]
  assign io_rPort_2_output_0 = _T_1103 ? Mem1D_3_io_output : _T_1114; // @[MemPrimitives.scala 148:13:@14300.4]
  assign io_rPort_1_output_0 = _T_1068 ? Mem1D_3_io_output : _T_1079; // @[MemPrimitives.scala 148:13:@14252.4]
  assign io_rPort_0_output_0 = _T_1033 ? Mem1D_1_io_output : _T_1044; // @[MemPrimitives.scala 148:13:@14204.4]
  assign Mem1D_clock = clock; // @[:@13278.4]
  assign Mem1D_reset = reset; // @[:@13279.4]
  assign Mem1D_io_r_ofs_0 = _T_635[0]; // @[MemPrimitives.scala 127:28:@13730.4]
  assign Mem1D_io_r_backpressure = _T_635[1]; // @[MemPrimitives.scala 128:32:@13731.4]
  assign Mem1D_io_w_ofs_0 = _T_465[0]; // @[MemPrimitives.scala 94:28:@13541.4]
  assign Mem1D_io_w_data_0 = _T_465[8:1]; // @[MemPrimitives.scala 95:29:@13542.4]
  assign Mem1D_io_w_en_0 = _T_465[9]; // @[MemPrimitives.scala 96:27:@13543.4]
  assign Mem1D_1_clock = clock; // @[:@13294.4]
  assign Mem1D_1_reset = reset; // @[:@13295.4]
  assign Mem1D_1_io_r_ofs_0 = _T_655[0]; // @[MemPrimitives.scala 127:28:@13754.4]
  assign Mem1D_1_io_r_backpressure = _T_655[1]; // @[MemPrimitives.scala 128:32:@13755.4]
  assign Mem1D_1_io_w_ofs_0 = _T_475[0]; // @[MemPrimitives.scala 94:28:@13552.4]
  assign Mem1D_1_io_w_data_0 = _T_475[8:1]; // @[MemPrimitives.scala 95:29:@13553.4]
  assign Mem1D_1_io_w_en_0 = _T_475[9]; // @[MemPrimitives.scala 96:27:@13554.4]
  assign Mem1D_2_clock = clock; // @[:@13310.4]
  assign Mem1D_2_reset = reset; // @[:@13311.4]
  assign Mem1D_2_io_r_ofs_0 = _T_675[0]; // @[MemPrimitives.scala 127:28:@13778.4]
  assign Mem1D_2_io_r_backpressure = _T_675[1]; // @[MemPrimitives.scala 128:32:@13779.4]
  assign Mem1D_2_io_w_ofs_0 = _T_485[0]; // @[MemPrimitives.scala 94:28:@13563.4]
  assign Mem1D_2_io_w_data_0 = _T_485[8:1]; // @[MemPrimitives.scala 95:29:@13564.4]
  assign Mem1D_2_io_w_en_0 = _T_485[9]; // @[MemPrimitives.scala 96:27:@13565.4]
  assign Mem1D_3_clock = clock; // @[:@13326.4]
  assign Mem1D_3_reset = reset; // @[:@13327.4]
  assign Mem1D_3_io_r_ofs_0 = _T_713[0]; // @[MemPrimitives.scala 127:28:@13818.4]
  assign Mem1D_3_io_r_backpressure = _T_713[1]; // @[MemPrimitives.scala 128:32:@13819.4]
  assign Mem1D_3_io_w_ofs_0 = _T_495[0]; // @[MemPrimitives.scala 94:28:@13574.4]
  assign Mem1D_3_io_w_data_0 = _T_495[8:1]; // @[MemPrimitives.scala 95:29:@13575.4]
  assign Mem1D_3_io_w_en_0 = _T_495[9]; // @[MemPrimitives.scala 96:27:@13576.4]
  assign Mem1D_4_clock = clock; // @[:@13342.4]
  assign Mem1D_4_reset = reset; // @[:@13343.4]
  assign Mem1D_4_io_r_ofs_0 = _T_733[0]; // @[MemPrimitives.scala 127:28:@13842.4]
  assign Mem1D_4_io_r_backpressure = _T_733[1]; // @[MemPrimitives.scala 128:32:@13843.4]
  assign Mem1D_4_io_w_ofs_0 = _T_505[0]; // @[MemPrimitives.scala 94:28:@13585.4]
  assign Mem1D_4_io_w_data_0 = _T_505[8:1]; // @[MemPrimitives.scala 95:29:@13586.4]
  assign Mem1D_4_io_w_en_0 = _T_505[9]; // @[MemPrimitives.scala 96:27:@13587.4]
  assign Mem1D_5_clock = clock; // @[:@13358.4]
  assign Mem1D_5_reset = reset; // @[:@13359.4]
  assign Mem1D_5_io_r_ofs_0 = _T_753[0]; // @[MemPrimitives.scala 127:28:@13866.4]
  assign Mem1D_5_io_r_backpressure = _T_753[1]; // @[MemPrimitives.scala 128:32:@13867.4]
  assign Mem1D_5_io_w_ofs_0 = _T_515[0]; // @[MemPrimitives.scala 94:28:@13596.4]
  assign Mem1D_5_io_w_data_0 = _T_515[8:1]; // @[MemPrimitives.scala 95:29:@13597.4]
  assign Mem1D_5_io_w_en_0 = _T_515[9]; // @[MemPrimitives.scala 96:27:@13598.4]
  assign Mem1D_6_clock = clock; // @[:@13374.4]
  assign Mem1D_6_reset = reset; // @[:@13375.4]
  assign Mem1D_6_io_r_ofs_0 = _T_773[0]; // @[MemPrimitives.scala 127:28:@13890.4]
  assign Mem1D_6_io_r_backpressure = _T_773[1]; // @[MemPrimitives.scala 128:32:@13891.4]
  assign Mem1D_6_io_w_ofs_0 = _T_525[0]; // @[MemPrimitives.scala 94:28:@13607.4]
  assign Mem1D_6_io_w_data_0 = _T_525[8:1]; // @[MemPrimitives.scala 95:29:@13608.4]
  assign Mem1D_6_io_w_en_0 = _T_525[9]; // @[MemPrimitives.scala 96:27:@13609.4]
  assign Mem1D_7_clock = clock; // @[:@13390.4]
  assign Mem1D_7_reset = reset; // @[:@13391.4]
  assign Mem1D_7_io_r_ofs_0 = _T_811[0]; // @[MemPrimitives.scala 127:28:@13930.4]
  assign Mem1D_7_io_r_backpressure = _T_811[1]; // @[MemPrimitives.scala 128:32:@13931.4]
  assign Mem1D_7_io_w_ofs_0 = _T_535[0]; // @[MemPrimitives.scala 94:28:@13618.4]
  assign Mem1D_7_io_w_data_0 = _T_535[8:1]; // @[MemPrimitives.scala 95:29:@13619.4]
  assign Mem1D_7_io_w_en_0 = _T_535[9]; // @[MemPrimitives.scala 96:27:@13620.4]
  assign Mem1D_8_clock = clock; // @[:@13406.4]
  assign Mem1D_8_reset = reset; // @[:@13407.4]
  assign Mem1D_8_io_r_ofs_0 = _T_831[0]; // @[MemPrimitives.scala 127:28:@13954.4]
  assign Mem1D_8_io_r_backpressure = _T_831[1]; // @[MemPrimitives.scala 128:32:@13955.4]
  assign Mem1D_8_io_w_ofs_0 = _T_545[0]; // @[MemPrimitives.scala 94:28:@13629.4]
  assign Mem1D_8_io_w_data_0 = _T_545[8:1]; // @[MemPrimitives.scala 95:29:@13630.4]
  assign Mem1D_8_io_w_en_0 = _T_545[9]; // @[MemPrimitives.scala 96:27:@13631.4]
  assign Mem1D_9_clock = clock; // @[:@13422.4]
  assign Mem1D_9_reset = reset; // @[:@13423.4]
  assign Mem1D_9_io_r_ofs_0 = _T_851[0]; // @[MemPrimitives.scala 127:28:@13978.4]
  assign Mem1D_9_io_r_backpressure = _T_851[1]; // @[MemPrimitives.scala 128:32:@13979.4]
  assign Mem1D_9_io_w_ofs_0 = _T_555[0]; // @[MemPrimitives.scala 94:28:@13640.4]
  assign Mem1D_9_io_w_data_0 = _T_555[8:1]; // @[MemPrimitives.scala 95:29:@13641.4]
  assign Mem1D_9_io_w_en_0 = _T_555[9]; // @[MemPrimitives.scala 96:27:@13642.4]
  assign Mem1D_10_clock = clock; // @[:@13438.4]
  assign Mem1D_10_reset = reset; // @[:@13439.4]
  assign Mem1D_10_io_r_ofs_0 = _T_871[0]; // @[MemPrimitives.scala 127:28:@14002.4]
  assign Mem1D_10_io_r_backpressure = _T_871[1]; // @[MemPrimitives.scala 128:32:@14003.4]
  assign Mem1D_10_io_w_ofs_0 = _T_565[0]; // @[MemPrimitives.scala 94:28:@13651.4]
  assign Mem1D_10_io_w_data_0 = _T_565[8:1]; // @[MemPrimitives.scala 95:29:@13652.4]
  assign Mem1D_10_io_w_en_0 = _T_565[9]; // @[MemPrimitives.scala 96:27:@13653.4]
  assign Mem1D_11_clock = clock; // @[:@13454.4]
  assign Mem1D_11_reset = reset; // @[:@13455.4]
  assign Mem1D_11_io_r_ofs_0 = _T_909[0]; // @[MemPrimitives.scala 127:28:@14042.4]
  assign Mem1D_11_io_r_backpressure = _T_909[1]; // @[MemPrimitives.scala 128:32:@14043.4]
  assign Mem1D_11_io_w_ofs_0 = _T_575[0]; // @[MemPrimitives.scala 94:28:@13662.4]
  assign Mem1D_11_io_w_data_0 = _T_575[8:1]; // @[MemPrimitives.scala 95:29:@13663.4]
  assign Mem1D_11_io_w_en_0 = _T_575[9]; // @[MemPrimitives.scala 96:27:@13664.4]
  assign Mem1D_12_clock = clock; // @[:@13470.4]
  assign Mem1D_12_reset = reset; // @[:@13471.4]
  assign Mem1D_12_io_r_ofs_0 = _T_929[0]; // @[MemPrimitives.scala 127:28:@14066.4]
  assign Mem1D_12_io_r_backpressure = _T_929[1]; // @[MemPrimitives.scala 128:32:@14067.4]
  assign Mem1D_12_io_w_ofs_0 = _T_585[0]; // @[MemPrimitives.scala 94:28:@13673.4]
  assign Mem1D_12_io_w_data_0 = _T_585[8:1]; // @[MemPrimitives.scala 95:29:@13674.4]
  assign Mem1D_12_io_w_en_0 = _T_585[9]; // @[MemPrimitives.scala 96:27:@13675.4]
  assign Mem1D_13_clock = clock; // @[:@13486.4]
  assign Mem1D_13_reset = reset; // @[:@13487.4]
  assign Mem1D_13_io_r_ofs_0 = _T_949[0]; // @[MemPrimitives.scala 127:28:@14090.4]
  assign Mem1D_13_io_r_backpressure = _T_949[1]; // @[MemPrimitives.scala 128:32:@14091.4]
  assign Mem1D_13_io_w_ofs_0 = _T_595[0]; // @[MemPrimitives.scala 94:28:@13684.4]
  assign Mem1D_13_io_w_data_0 = _T_595[8:1]; // @[MemPrimitives.scala 95:29:@13685.4]
  assign Mem1D_13_io_w_en_0 = _T_595[9]; // @[MemPrimitives.scala 96:27:@13686.4]
  assign Mem1D_14_clock = clock; // @[:@13502.4]
  assign Mem1D_14_reset = reset; // @[:@13503.4]
  assign Mem1D_14_io_r_ofs_0 = _T_969[0]; // @[MemPrimitives.scala 127:28:@14114.4]
  assign Mem1D_14_io_r_backpressure = _T_969[1]; // @[MemPrimitives.scala 128:32:@14115.4]
  assign Mem1D_14_io_w_ofs_0 = _T_605[0]; // @[MemPrimitives.scala 94:28:@13695.4]
  assign Mem1D_14_io_w_data_0 = _T_605[8:1]; // @[MemPrimitives.scala 95:29:@13696.4]
  assign Mem1D_14_io_w_en_0 = _T_605[9]; // @[MemPrimitives.scala 96:27:@13697.4]
  assign Mem1D_15_clock = clock; // @[:@13518.4]
  assign Mem1D_15_reset = reset; // @[:@13519.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1007[0]; // @[MemPrimitives.scala 127:28:@14154.4]
  assign Mem1D_15_io_r_backpressure = _T_1007[1]; // @[MemPrimitives.scala 128:32:@14155.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[0]; // @[MemPrimitives.scala 94:28:@13706.4]
  assign Mem1D_15_io_w_data_0 = _T_615[8:1]; // @[MemPrimitives.scala 95:29:@13707.4]
  assign Mem1D_15_io_w_en_0 = _T_615[9]; // @[MemPrimitives.scala 96:27:@13708.4]
  assign StickySelects_clock = clock; // @[:@13716.4]
  assign StickySelects_reset = reset; // @[:@13717.4]
  assign StickySelects_io_ins_0 = io_rPort_5_en_0 & _T_620; // @[MemPrimitives.scala 122:60:@13718.4]
  assign StickySelects_io_ins_1 = io_rPort_6_en_0 & _T_625; // @[MemPrimitives.scala 122:60:@13719.4]
  assign StickySelects_1_clock = clock; // @[:@13740.4]
  assign StickySelects_1_reset = reset; // @[:@13741.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_640; // @[MemPrimitives.scala 122:60:@13742.4]
  assign StickySelects_1_io_ins_1 = io_rPort_7_en_0 & _T_645; // @[MemPrimitives.scala 122:60:@13743.4]
  assign StickySelects_2_clock = clock; // @[:@13764.4]
  assign StickySelects_2_reset = reset; // @[:@13765.4]
  assign StickySelects_2_io_ins_0 = io_rPort_3_en_0 & _T_660; // @[MemPrimitives.scala 122:60:@13766.4]
  assign StickySelects_2_io_ins_1 = io_rPort_9_en_0 & _T_665; // @[MemPrimitives.scala 122:60:@13767.4]
  assign StickySelects_3_clock = clock; // @[:@13794.4]
  assign StickySelects_3_reset = reset; // @[:@13795.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_680; // @[MemPrimitives.scala 122:60:@13796.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_685; // @[MemPrimitives.scala 122:60:@13797.4]
  assign StickySelects_3_io_ins_2 = io_rPort_4_en_0 & _T_690; // @[MemPrimitives.scala 122:60:@13798.4]
  assign StickySelects_3_io_ins_3 = io_rPort_8_en_0 & _T_695; // @[MemPrimitives.scala 122:60:@13799.4]
  assign StickySelects_4_clock = clock; // @[:@13828.4]
  assign StickySelects_4_reset = reset; // @[:@13829.4]
  assign StickySelects_4_io_ins_0 = io_rPort_5_en_0 & _T_718; // @[MemPrimitives.scala 122:60:@13830.4]
  assign StickySelects_4_io_ins_1 = io_rPort_6_en_0 & _T_723; // @[MemPrimitives.scala 122:60:@13831.4]
  assign StickySelects_5_clock = clock; // @[:@13852.4]
  assign StickySelects_5_reset = reset; // @[:@13853.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_738; // @[MemPrimitives.scala 122:60:@13854.4]
  assign StickySelects_5_io_ins_1 = io_rPort_7_en_0 & _T_743; // @[MemPrimitives.scala 122:60:@13855.4]
  assign StickySelects_6_clock = clock; // @[:@13876.4]
  assign StickySelects_6_reset = reset; // @[:@13877.4]
  assign StickySelects_6_io_ins_0 = io_rPort_3_en_0 & _T_758; // @[MemPrimitives.scala 122:60:@13878.4]
  assign StickySelects_6_io_ins_1 = io_rPort_9_en_0 & _T_763; // @[MemPrimitives.scala 122:60:@13879.4]
  assign StickySelects_7_clock = clock; // @[:@13906.4]
  assign StickySelects_7_reset = reset; // @[:@13907.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_778; // @[MemPrimitives.scala 122:60:@13908.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_783; // @[MemPrimitives.scala 122:60:@13909.4]
  assign StickySelects_7_io_ins_2 = io_rPort_4_en_0 & _T_788; // @[MemPrimitives.scala 122:60:@13910.4]
  assign StickySelects_7_io_ins_3 = io_rPort_8_en_0 & _T_793; // @[MemPrimitives.scala 122:60:@13911.4]
  assign StickySelects_8_clock = clock; // @[:@13940.4]
  assign StickySelects_8_reset = reset; // @[:@13941.4]
  assign StickySelects_8_io_ins_0 = io_rPort_5_en_0 & _T_816; // @[MemPrimitives.scala 122:60:@13942.4]
  assign StickySelects_8_io_ins_1 = io_rPort_6_en_0 & _T_821; // @[MemPrimitives.scala 122:60:@13943.4]
  assign StickySelects_9_clock = clock; // @[:@13964.4]
  assign StickySelects_9_reset = reset; // @[:@13965.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_836; // @[MemPrimitives.scala 122:60:@13966.4]
  assign StickySelects_9_io_ins_1 = io_rPort_7_en_0 & _T_841; // @[MemPrimitives.scala 122:60:@13967.4]
  assign StickySelects_10_clock = clock; // @[:@13988.4]
  assign StickySelects_10_reset = reset; // @[:@13989.4]
  assign StickySelects_10_io_ins_0 = io_rPort_3_en_0 & _T_856; // @[MemPrimitives.scala 122:60:@13990.4]
  assign StickySelects_10_io_ins_1 = io_rPort_9_en_0 & _T_861; // @[MemPrimitives.scala 122:60:@13991.4]
  assign StickySelects_11_clock = clock; // @[:@14018.4]
  assign StickySelects_11_reset = reset; // @[:@14019.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_876; // @[MemPrimitives.scala 122:60:@14020.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_881; // @[MemPrimitives.scala 122:60:@14021.4]
  assign StickySelects_11_io_ins_2 = io_rPort_4_en_0 & _T_886; // @[MemPrimitives.scala 122:60:@14022.4]
  assign StickySelects_11_io_ins_3 = io_rPort_8_en_0 & _T_891; // @[MemPrimitives.scala 122:60:@14023.4]
  assign StickySelects_12_clock = clock; // @[:@14052.4]
  assign StickySelects_12_reset = reset; // @[:@14053.4]
  assign StickySelects_12_io_ins_0 = io_rPort_5_en_0 & _T_914; // @[MemPrimitives.scala 122:60:@14054.4]
  assign StickySelects_12_io_ins_1 = io_rPort_6_en_0 & _T_919; // @[MemPrimitives.scala 122:60:@14055.4]
  assign StickySelects_13_clock = clock; // @[:@14076.4]
  assign StickySelects_13_reset = reset; // @[:@14077.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_934; // @[MemPrimitives.scala 122:60:@14078.4]
  assign StickySelects_13_io_ins_1 = io_rPort_7_en_0 & _T_939; // @[MemPrimitives.scala 122:60:@14079.4]
  assign StickySelects_14_clock = clock; // @[:@14100.4]
  assign StickySelects_14_reset = reset; // @[:@14101.4]
  assign StickySelects_14_io_ins_0 = io_rPort_3_en_0 & _T_954; // @[MemPrimitives.scala 122:60:@14102.4]
  assign StickySelects_14_io_ins_1 = io_rPort_9_en_0 & _T_959; // @[MemPrimitives.scala 122:60:@14103.4]
  assign StickySelects_15_clock = clock; // @[:@14130.4]
  assign StickySelects_15_reset = reset; // @[:@14131.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_974; // @[MemPrimitives.scala 122:60:@14132.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_979; // @[MemPrimitives.scala 122:60:@14133.4]
  assign StickySelects_15_io_ins_2 = io_rPort_4_en_0 & _T_984; // @[MemPrimitives.scala 122:60:@14134.4]
  assign StickySelects_15_io_ins_3 = io_rPort_8_en_0 & _T_989; // @[MemPrimitives.scala 122:60:@14135.4]
  assign RetimeWrapper_clock = clock; // @[:@14171.4]
  assign RetimeWrapper_reset = reset; // @[:@14172.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14174.4]
  assign RetimeWrapper_io_in = _T_640 & io_rPort_0_en_0; // @[package.scala 94:16:@14173.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14179.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14180.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14182.4]
  assign RetimeWrapper_1_io_in = _T_738 & io_rPort_0_en_0; // @[package.scala 94:16:@14181.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14187.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14188.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14190.4]
  assign RetimeWrapper_2_io_in = _T_836 & io_rPort_0_en_0; // @[package.scala 94:16:@14189.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14195.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14196.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14198.4]
  assign RetimeWrapper_3_io_in = _T_934 & io_rPort_0_en_0; // @[package.scala 94:16:@14197.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14219.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14220.4]
  assign RetimeWrapper_4_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14222.4]
  assign RetimeWrapper_4_io_in = _T_680 & io_rPort_1_en_0; // @[package.scala 94:16:@14221.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14227.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14228.4]
  assign RetimeWrapper_5_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14230.4]
  assign RetimeWrapper_5_io_in = _T_778 & io_rPort_1_en_0; // @[package.scala 94:16:@14229.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14235.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14236.4]
  assign RetimeWrapper_6_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14238.4]
  assign RetimeWrapper_6_io_in = _T_876 & io_rPort_1_en_0; // @[package.scala 94:16:@14237.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14243.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14244.4]
  assign RetimeWrapper_7_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14246.4]
  assign RetimeWrapper_7_io_in = _T_974 & io_rPort_1_en_0; // @[package.scala 94:16:@14245.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14267.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14268.4]
  assign RetimeWrapper_8_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14270.4]
  assign RetimeWrapper_8_io_in = _T_685 & io_rPort_2_en_0; // @[package.scala 94:16:@14269.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14275.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14276.4]
  assign RetimeWrapper_9_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14278.4]
  assign RetimeWrapper_9_io_in = _T_783 & io_rPort_2_en_0; // @[package.scala 94:16:@14277.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14283.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14284.4]
  assign RetimeWrapper_10_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14286.4]
  assign RetimeWrapper_10_io_in = _T_881 & io_rPort_2_en_0; // @[package.scala 94:16:@14285.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14291.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14292.4]
  assign RetimeWrapper_11_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14294.4]
  assign RetimeWrapper_11_io_in = _T_979 & io_rPort_2_en_0; // @[package.scala 94:16:@14293.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14315.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14316.4]
  assign RetimeWrapper_12_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14318.4]
  assign RetimeWrapper_12_io_in = _T_660 & io_rPort_3_en_0; // @[package.scala 94:16:@14317.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14323.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14324.4]
  assign RetimeWrapper_13_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14326.4]
  assign RetimeWrapper_13_io_in = _T_758 & io_rPort_3_en_0; // @[package.scala 94:16:@14325.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14331.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14332.4]
  assign RetimeWrapper_14_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14334.4]
  assign RetimeWrapper_14_io_in = _T_856 & io_rPort_3_en_0; // @[package.scala 94:16:@14333.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14339.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14340.4]
  assign RetimeWrapper_15_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14342.4]
  assign RetimeWrapper_15_io_in = _T_954 & io_rPort_3_en_0; // @[package.scala 94:16:@14341.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14363.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14364.4]
  assign RetimeWrapper_16_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14366.4]
  assign RetimeWrapper_16_io_in = _T_690 & io_rPort_4_en_0; // @[package.scala 94:16:@14365.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14371.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14372.4]
  assign RetimeWrapper_17_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14374.4]
  assign RetimeWrapper_17_io_in = _T_788 & io_rPort_4_en_0; // @[package.scala 94:16:@14373.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14379.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14380.4]
  assign RetimeWrapper_18_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14382.4]
  assign RetimeWrapper_18_io_in = _T_886 & io_rPort_4_en_0; // @[package.scala 94:16:@14381.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14387.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14388.4]
  assign RetimeWrapper_19_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14390.4]
  assign RetimeWrapper_19_io_in = _T_984 & io_rPort_4_en_0; // @[package.scala 94:16:@14389.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14411.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14412.4]
  assign RetimeWrapper_20_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14414.4]
  assign RetimeWrapper_20_io_in = _T_620 & io_rPort_5_en_0; // @[package.scala 94:16:@14413.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14419.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14420.4]
  assign RetimeWrapper_21_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14422.4]
  assign RetimeWrapper_21_io_in = _T_718 & io_rPort_5_en_0; // @[package.scala 94:16:@14421.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14427.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14428.4]
  assign RetimeWrapper_22_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14430.4]
  assign RetimeWrapper_22_io_in = _T_816 & io_rPort_5_en_0; // @[package.scala 94:16:@14429.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14435.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14436.4]
  assign RetimeWrapper_23_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14438.4]
  assign RetimeWrapper_23_io_in = _T_914 & io_rPort_5_en_0; // @[package.scala 94:16:@14437.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14459.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14460.4]
  assign RetimeWrapper_24_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14462.4]
  assign RetimeWrapper_24_io_in = _T_625 & io_rPort_6_en_0; // @[package.scala 94:16:@14461.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14467.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14468.4]
  assign RetimeWrapper_25_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14470.4]
  assign RetimeWrapper_25_io_in = _T_723 & io_rPort_6_en_0; // @[package.scala 94:16:@14469.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14475.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14476.4]
  assign RetimeWrapper_26_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14478.4]
  assign RetimeWrapper_26_io_in = _T_821 & io_rPort_6_en_0; // @[package.scala 94:16:@14477.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14483.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14484.4]
  assign RetimeWrapper_27_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14486.4]
  assign RetimeWrapper_27_io_in = _T_919 & io_rPort_6_en_0; // @[package.scala 94:16:@14485.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14507.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14508.4]
  assign RetimeWrapper_28_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14510.4]
  assign RetimeWrapper_28_io_in = _T_645 & io_rPort_7_en_0; // @[package.scala 94:16:@14509.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14515.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14516.4]
  assign RetimeWrapper_29_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14518.4]
  assign RetimeWrapper_29_io_in = _T_743 & io_rPort_7_en_0; // @[package.scala 94:16:@14517.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14523.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14524.4]
  assign RetimeWrapper_30_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14526.4]
  assign RetimeWrapper_30_io_in = _T_841 & io_rPort_7_en_0; // @[package.scala 94:16:@14525.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14531.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14532.4]
  assign RetimeWrapper_31_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14534.4]
  assign RetimeWrapper_31_io_in = _T_939 & io_rPort_7_en_0; // @[package.scala 94:16:@14533.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14555.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14556.4]
  assign RetimeWrapper_32_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14558.4]
  assign RetimeWrapper_32_io_in = _T_695 & io_rPort_8_en_0; // @[package.scala 94:16:@14557.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14563.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14564.4]
  assign RetimeWrapper_33_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14566.4]
  assign RetimeWrapper_33_io_in = _T_793 & io_rPort_8_en_0; // @[package.scala 94:16:@14565.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14571.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14572.4]
  assign RetimeWrapper_34_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14574.4]
  assign RetimeWrapper_34_io_in = _T_891 & io_rPort_8_en_0; // @[package.scala 94:16:@14573.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14579.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14580.4]
  assign RetimeWrapper_35_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14582.4]
  assign RetimeWrapper_35_io_in = _T_989 & io_rPort_8_en_0; // @[package.scala 94:16:@14581.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14603.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14604.4]
  assign RetimeWrapper_36_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14606.4]
  assign RetimeWrapper_36_io_in = _T_665 & io_rPort_9_en_0; // @[package.scala 94:16:@14605.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14611.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14612.4]
  assign RetimeWrapper_37_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14614.4]
  assign RetimeWrapper_37_io_in = _T_763 & io_rPort_9_en_0; // @[package.scala 94:16:@14613.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14619.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14620.4]
  assign RetimeWrapper_38_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14622.4]
  assign RetimeWrapper_38_io_in = _T_861 & io_rPort_9_en_0; // @[package.scala 94:16:@14621.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14627.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14628.4]
  assign RetimeWrapper_39_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14630.4]
  assign RetimeWrapper_39_io_in = _T_959 & io_rPort_9_en_0; // @[package.scala 94:16:@14629.4]
endmodule
module RetimeWrapper_196( // @[:@14650.2]
  input         clock, // @[:@14651.4]
  input         reset, // @[:@14652.4]
  input         io_flow, // @[:@14653.4]
  input  [31:0] io_in, // @[:@14653.4]
  output [31:0] io_out // @[:@14653.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14655.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14655.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14655.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14655.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14655.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14655.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@14655.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14668.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14667.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14666.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14665.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14664.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14662.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@14670.2]
  input  [31:0] io_a, // @[:@14673.4]
  output [32:0] io_b // @[:@14673.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@14680.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@14680.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@14685.4]
endmodule
module __2( // @[:@14687.2]
  input  [31:0] io_b, // @[:@14690.4]
  output [32:0] io_result // @[:@14690.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@14695.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@14695.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@14695.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@14708.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@14703.4]
endmodule
module fix2fixBox( // @[:@14782.2]
  input         clock, // @[:@14783.4]
  input         reset, // @[:@14784.4]
  input  [32:0] io_a, // @[:@14785.4]
  input         io_flow, // @[:@14785.4]
  output [31:0] io_b // @[:@14785.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14795.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14795.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14795.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@14795.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@14795.4]
  RetimeWrapper_196 RetimeWrapper ( // @[package.scala 93:22:@14795.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@14802.4]
  assign RetimeWrapper_clock = clock; // @[:@14796.4]
  assign RetimeWrapper_reset = reset; // @[:@14797.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@14799.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@14798.4]
endmodule
module x401_sum( // @[:@14804.2]
  input         clock, // @[:@14805.4]
  input         reset, // @[:@14806.4]
  input  [31:0] io_a, // @[:@14807.4]
  input  [31:0] io_b, // @[:@14807.4]
  input         io_flow, // @[:@14807.4]
  output [31:0] io_result // @[:@14807.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@14815.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@14815.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@14822.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@14822.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@14840.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@14840.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@14840.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@14840.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@14840.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@14820.4 Math.scala 713:14:@14821.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@14827.4 Math.scala 713:14:@14828.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@14829.4]
  __2 _ ( // @[Math.scala 709:24:@14815.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@14822.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@14840.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@14820.4 Math.scala 713:14:@14821.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@14827.4 Math.scala 713:14:@14828.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@14829.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@14848.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@14818.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@14825.4]
  assign fix2fixBox_clock = clock; // @[:@14841.4]
  assign fix2fixBox_reset = reset; // @[:@14842.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@14843.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@14846.4]
endmodule
module RetimeWrapper_198( // @[:@14862.2]
  input   clock, // @[:@14863.4]
  input   reset, // @[:@14864.4]
  input   io_flow, // @[:@14865.4]
  input   io_in, // @[:@14865.4]
  output  io_out // @[:@14865.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@14867.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@14867.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@14867.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14867.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14867.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14867.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@14867.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14880.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14879.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@14878.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14877.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14876.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14874.4]
endmodule
module RetimeWrapper_200( // @[:@14926.2]
  input        clock, // @[:@14927.4]
  input        reset, // @[:@14928.4]
  input        io_flow, // @[:@14929.4]
  input  [7:0] io_in, // @[:@14929.4]
  output [7:0] io_out // @[:@14929.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14931.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14931.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14931.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14931.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14931.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14931.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@14931.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14944.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14943.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@14942.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14941.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14940.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14938.4]
endmodule
module RetimeWrapper_201( // @[:@14958.2]
  input         clock, // @[:@14959.4]
  input         reset, // @[:@14960.4]
  input         io_flow, // @[:@14961.4]
  input  [31:0] io_in, // @[:@14961.4]
  output [31:0] io_out // @[:@14961.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14963.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14963.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14963.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14963.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14963.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14963.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@14963.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@14976.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@14975.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@14974.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@14973.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@14972.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@14970.4]
endmodule
module RetimeWrapper_202( // @[:@14990.2]
  input         clock, // @[:@14991.4]
  input         reset, // @[:@14992.4]
  input         io_flow, // @[:@14993.4]
  input  [31:0] io_in, // @[:@14993.4]
  output [31:0] io_out // @[:@14993.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@14995.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@14995.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@14995.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@14995.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@14995.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@14995.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@14995.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15008.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15007.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15006.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15005.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15004.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15002.4]
endmodule
module RetimeWrapper_208( // @[:@15478.2]
  input         clock, // @[:@15479.4]
  input         reset, // @[:@15480.4]
  input         io_flow, // @[:@15481.4]
  input  [31:0] io_in, // @[:@15481.4]
  output [31:0] io_out // @[:@15481.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15483.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15483.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15483.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15483.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15483.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15483.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15483.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15496.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15495.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15494.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15493.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15492.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15490.4]
endmodule
module RetimeWrapper_220( // @[:@16454.2]
  input         clock, // @[:@16455.4]
  input         reset, // @[:@16456.4]
  input         io_flow, // @[:@16457.4]
  input  [31:0] io_in, // @[:@16457.4]
  output [31:0] io_out // @[:@16457.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16459.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16459.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16459.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16459.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16459.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16459.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@16459.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16472.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16471.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16470.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16469.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16468.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16466.4]
endmodule
module RetimeWrapper_226( // @[:@16794.2]
  input   clock, // @[:@16795.4]
  input   reset, // @[:@16796.4]
  input   io_flow, // @[:@16797.4]
  input   io_in, // @[:@16797.4]
  output  io_out // @[:@16797.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@16799.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@16799.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@16799.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16799.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16799.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16799.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@16799.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16812.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16811.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@16810.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16809.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16808.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16806.4]
endmodule
module x496_rdrow( // @[:@18880.2]
  input         clock, // @[:@18881.4]
  input         reset, // @[:@18882.4]
  input  [31:0] io_a, // @[:@18883.4]
  input  [31:0] io_b, // @[:@18883.4]
  input         io_flow, // @[:@18883.4]
  output [31:0] io_result // @[:@18883.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@18891.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@18891.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@18898.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@18898.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@18917.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@18917.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@18917.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@18917.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@18917.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@18896.4 Math.scala 713:14:@18897.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@18903.4 Math.scala 713:14:@18904.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@18905.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@18906.4]
  __2 _ ( // @[Math.scala 709:24:@18891.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@18898.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@18917.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@18896.4 Math.scala 713:14:@18897.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@18903.4 Math.scala 713:14:@18904.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@18905.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@18906.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@18925.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@18894.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@18901.4]
  assign fix2fixBox_clock = clock; // @[:@18918.4]
  assign fix2fixBox_reset = reset; // @[:@18919.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@18920.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@18923.4]
endmodule
module RetimeWrapper_267( // @[:@19735.2]
  input         clock, // @[:@19736.4]
  input         reset, // @[:@19737.4]
  input         io_flow, // @[:@19738.4]
  input  [31:0] io_in, // @[:@19738.4]
  output [31:0] io_out // @[:@19738.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@19740.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@19740.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@19740.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@19740.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@19740.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@19740.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@19740.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@19753.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@19752.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@19751.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@19750.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@19749.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@19747.4]
endmodule
module SimBlackBoxesfix2fixBox_60( // @[:@22164.2]
  input  [7:0] io_a, // @[:@22167.4]
  output [8:0] io_b // @[:@22167.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@22178.4]
endmodule
module __60( // @[:@22180.2]
  input  [7:0] io_b, // @[:@22183.4]
  output [8:0] io_result // @[:@22183.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@22188.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@22188.4]
  SimBlackBoxesfix2fixBox_60 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@22188.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@22201.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@22196.4]
endmodule
module fix2fixBox_29( // @[:@22274.2]
  input        clock, // @[:@22275.4]
  input        reset, // @[:@22276.4]
  input  [8:0] io_a, // @[:@22277.4]
  input        io_flow, // @[:@22277.4]
  output [7:0] io_b // @[:@22277.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22287.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22287.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22287.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@22287.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@22287.4]
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@22287.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@22294.4]
  assign RetimeWrapper_clock = clock; // @[:@22288.4]
  assign RetimeWrapper_reset = reset; // @[:@22289.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@22291.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@22290.4]
endmodule
module x597_x23( // @[:@22296.2]
  input        clock, // @[:@22297.4]
  input        reset, // @[:@22298.4]
  input  [7:0] io_a, // @[:@22299.4]
  input  [7:0] io_b, // @[:@22299.4]
  input        io_flow, // @[:@22299.4]
  output [7:0] io_result // @[:@22299.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22307.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22307.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22314.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22314.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@22324.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@22324.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22324.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@22324.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22324.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22312.4 Math.scala 713:14:@22313.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22319.4 Math.scala 713:14:@22320.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22321.4]
  __60 _ ( // @[Math.scala 709:24:@22307.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __60 __1 ( // @[Math.scala 709:24:@22314.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_29 fix2fixBox ( // @[Math.scala 141:30:@22324.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22312.4 Math.scala 713:14:@22313.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22319.4 Math.scala 713:14:@22320.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22321.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22332.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22310.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22317.4]
  assign fix2fixBox_clock = clock; // @[:@22325.4]
  assign fix2fixBox_reset = reset; // @[:@22326.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22327.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@22330.4]
endmodule
module fix2fixBox_33( // @[:@22922.2]
  input  [8:0] io_a, // @[:@22925.4]
  output [7:0] io_b // @[:@22925.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@22935.4]
endmodule
module x601_x23( // @[:@22937.2]
  input  [7:0] io_a, // @[:@22940.4]
  input  [7:0] io_b, // @[:@22940.4]
  output [7:0] io_result // @[:@22940.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22948.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22948.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22955.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22955.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22965.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22965.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22953.4 Math.scala 713:14:@22954.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22960.4 Math.scala 713:14:@22961.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22962.4]
  __60 _ ( // @[Math.scala 709:24:@22948.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __60 __1 ( // @[Math.scala 709:24:@22955.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_33 fix2fixBox ( // @[Math.scala 141:30:@22965.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22953.4 Math.scala 713:14:@22954.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22960.4 Math.scala 713:14:@22961.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22962.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22973.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22951.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22958.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22968.4]
endmodule
module RetimeWrapper_321( // @[:@27248.2]
  input   clock, // @[:@27249.4]
  input   reset, // @[:@27250.4]
  input   io_flow, // @[:@27251.4]
  input   io_in, // @[:@27251.4]
  output  io_out // @[:@27251.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@27253.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@27253.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@27253.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27253.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27253.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27253.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@27253.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27266.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27265.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@27264.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27263.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27262.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27260.4]
endmodule
module RetimeWrapper_323( // @[:@27312.2]
  input         clock, // @[:@27313.4]
  input         reset, // @[:@27314.4]
  input         io_flow, // @[:@27315.4]
  input  [31:0] io_in, // @[:@27315.4]
  output [31:0] io_out // @[:@27315.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27317.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27317.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27317.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27317.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27317.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27317.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@27317.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27330.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27329.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27328.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27327.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27326.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27324.4]
endmodule
module RetimeWrapper_324( // @[:@27344.2]
  input         clock, // @[:@27345.4]
  input         reset, // @[:@27346.4]
  input         io_flow, // @[:@27347.4]
  input  [31:0] io_in, // @[:@27347.4]
  output [31:0] io_out // @[:@27347.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27349.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27349.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27349.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27349.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27349.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27349.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@27349.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27362.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27361.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27360.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27359.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27358.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27356.4]
endmodule
module RetimeWrapper_326( // @[:@27408.2]
  input         clock, // @[:@27409.4]
  input         reset, // @[:@27410.4]
  input         io_flow, // @[:@27411.4]
  input  [31:0] io_in, // @[:@27411.4]
  output [31:0] io_out // @[:@27411.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27413.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27413.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27413.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27413.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27413.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27413.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@27413.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27426.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27425.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27424.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27423.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27422.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27420.4]
endmodule
module RetimeWrapper_333( // @[:@27632.2]
  input   clock, // @[:@27633.4]
  input   reset, // @[:@27634.4]
  input   io_flow, // @[:@27635.4]
  input   io_in, // @[:@27635.4]
  output  io_out // @[:@27635.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@27637.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@27637.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@27637.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27637.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27637.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27637.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@27637.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27650.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27649.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@27648.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27647.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27646.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27644.4]
endmodule
module RetimeWrapper_342( // @[:@27920.2]
  input         clock, // @[:@27921.4]
  input         reset, // @[:@27922.4]
  input         io_flow, // @[:@27923.4]
  input  [31:0] io_in, // @[:@27923.4]
  output [31:0] io_out // @[:@27923.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@27925.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@27925.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@27925.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27925.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27925.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27925.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@27925.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27938.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27937.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@27936.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27935.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27934.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27932.4]
endmodule
module RetimeWrapper_343( // @[:@27952.2]
  input   clock, // @[:@27953.4]
  input   reset, // @[:@27954.4]
  input   io_flow, // @[:@27955.4]
  input   io_in, // @[:@27955.4]
  output  io_out // @[:@27955.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@27957.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@27957.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@27957.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@27957.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@27957.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@27957.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@27957.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@27970.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@27969.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@27968.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@27967.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@27966.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@27964.4]
endmodule
module RetimeWrapper_364( // @[:@29017.2]
  input        clock, // @[:@29018.4]
  input        reset, // @[:@29019.4]
  input        io_flow, // @[:@29020.4]
  input  [7:0] io_in, // @[:@29020.4]
  output [7:0] io_out // @[:@29020.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@29022.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@29022.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@29022.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@29022.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@29022.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@29022.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@29022.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@29035.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@29034.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@29033.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@29032.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@29031.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@29029.4]
endmodule
module SimBlackBoxesfix2fixBox_130( // @[:@29037.2]
  input  [7:0] io_a, // @[:@29040.4]
  output [7:0] io_b // @[:@29040.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@29050.4]
endmodule
module __130( // @[:@29052.2]
  input  [7:0] io_b, // @[:@29055.4]
  output [7:0] io_result // @[:@29055.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@29060.4]
  wire [7:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@29060.4]
  SimBlackBoxesfix2fixBox_130 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@29060.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@29073.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@29068.4]
endmodule
module x677_div( // @[:@29075.2]
  input        clock, // @[:@29076.4]
  input        reset, // @[:@29077.4]
  input  [7:0] io_a, // @[:@29078.4]
  input        io_flow, // @[:@29078.4]
  output [7:0] io_result // @[:@29078.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29085.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29085.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29085.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@29085.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@29085.4]
  wire [7:0] __io_b; // @[Math.scala 709:24:@29095.4]
  wire [7:0] __io_result; // @[Math.scala 709:24:@29095.4]
  RetimeWrapper_364 RetimeWrapper ( // @[package.scala 93:22:@29085.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  __130 _ ( // @[Math.scala 709:24:@29095.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign io_result = __io_result; // @[Math.scala 291:34:@29103.4]
  assign RetimeWrapper_clock = clock; // @[:@29086.4]
  assign RetimeWrapper_reset = reset; // @[:@29087.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@29089.4]
  assign RetimeWrapper_io_in = io_a / 8'h6; // @[package.scala 94:16:@29088.4]
  assign __io_b = RetimeWrapper_io_out; // @[Math.scala 710:17:@29098.4]
endmodule
module RetimeWrapper_369( // @[:@30628.2]
  input   clock, // @[:@30629.4]
  input   reset, // @[:@30630.4]
  input   io_flow, // @[:@30631.4]
  input   io_in, // @[:@30631.4]
  output  io_out // @[:@30631.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30633.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30633.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30633.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30633.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30633.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30633.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@30633.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30646.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30645.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30644.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30643.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30642.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30640.4]
endmodule
module x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@30712.2]
  input          clock, // @[:@30713.4]
  input          reset, // @[:@30714.4]
  output         io_in_x374_TVALID, // @[:@30715.4]
  input          io_in_x374_TREADY, // @[:@30715.4]
  output [255:0] io_in_x374_TDATA, // @[:@30715.4]
  output         io_in_x373_TREADY, // @[:@30715.4]
  input  [255:0] io_in_x373_TDATA, // @[:@30715.4]
  input  [7:0]   io_in_x373_TID, // @[:@30715.4]
  input  [7:0]   io_in_x373_TDEST, // @[:@30715.4]
  input          io_sigsIn_backpressure, // @[:@30715.4]
  input          io_sigsIn_datapathEn, // @[:@30715.4]
  input          io_sigsIn_break, // @[:@30715.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@30715.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@30715.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@30715.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@30715.4]
  input          io_rr // @[:@30715.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@30729.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@30729.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@30741.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@30741.4]
  wire  x386_lb_0_clock; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_reset; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_17_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_17_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_17_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_17_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_17_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_16_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_16_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_16_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_16_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_16_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_15_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_15_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_15_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_15_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_15_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_14_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_14_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_14_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_14_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_14_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_13_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_13_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_13_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_13_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_13_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_12_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_12_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_12_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_12_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_12_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_11_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_11_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_11_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_11_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_11_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_10_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_10_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_10_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_10_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_10_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_9_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_9_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_9_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_9_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_9_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_8_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_8_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_8_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_8_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_8_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_7_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_7_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_7_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_7_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_7_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_6_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_6_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_6_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_6_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_6_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_5_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_5_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_5_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_5_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_5_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_4_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_4_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_4_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_4_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_4_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_3_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_3_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_3_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_3_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_3_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_2_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_2_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_2_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_2_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_2_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_1_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_1_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_1_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_1_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_1_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_rPort_0_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_0_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_0_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_rPort_0_backpressure; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_rPort_0_output_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_wPort_3_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_3_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_wPort_3_data_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_3_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_wPort_2_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_2_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_wPort_2_data_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_2_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_wPort_1_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_1_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_wPort_1_data_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_1_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [2:0] x386_lb_0_io_wPort_0_banks_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_0_ofs_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire [7:0] x386_lb_0_io_wPort_0_data_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x386_lb_0_io_wPort_0_en_0; // @[m_x386_lb_0.scala 47:17:@30751.4]
  wire  x387_lb2_0_clock; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_reset; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_9_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_9_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_9_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_9_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_9_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_8_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_8_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_8_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_8_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_8_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_7_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_7_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_7_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_7_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_7_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_6_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_6_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_6_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_6_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_6_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_5_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_5_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_5_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_5_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_5_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_4_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_4_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_4_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_4_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_4_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_3_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_3_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_3_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_3_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_3_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_2_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_2_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_2_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_2_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_2_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_1_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_1_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_1_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_1_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_1_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_rPort_0_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_0_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_0_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_rPort_0_backpressure; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_rPort_0_output_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_wPort_3_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_3_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_wPort_3_data_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_3_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_wPort_2_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_2_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_wPort_2_data_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_2_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_wPort_1_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_1_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_wPort_1_data_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_1_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [2:0] x387_lb2_0_io_wPort_0_banks_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_0_ofs_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire [7:0] x387_lb2_0_io_wPort_0_data_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  x387_lb2_0_io_wPort_0_en_0; // @[m_x387_lb2_0.scala 39:17:@30896.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31006.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31006.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31006.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@31006.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@31006.4]
  wire  x401_sum_1_clock; // @[Math.scala 150:24:@31106.4]
  wire  x401_sum_1_reset; // @[Math.scala 150:24:@31106.4]
  wire [31:0] x401_sum_1_io_a; // @[Math.scala 150:24:@31106.4]
  wire [31:0] x401_sum_1_io_b; // @[Math.scala 150:24:@31106.4]
  wire  x401_sum_1_io_flow; // @[Math.scala 150:24:@31106.4]
  wire [31:0] x401_sum_1_io_result; // @[Math.scala 150:24:@31106.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31116.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31116.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31116.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31116.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31116.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31125.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31125.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31125.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31125.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31125.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31134.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31134.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31134.4]
  wire [7:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@31134.4]
  wire [7:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@31134.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31143.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31143.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31143.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@31143.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@31143.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@31152.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@31152.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@31152.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@31152.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@31152.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@31165.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@31165.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@31165.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@31165.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@31165.4]
  wire  x407_rdcol_1_clock; // @[Math.scala 150:24:@31188.4]
  wire  x407_rdcol_1_reset; // @[Math.scala 150:24:@31188.4]
  wire [31:0] x407_rdcol_1_io_a; // @[Math.scala 150:24:@31188.4]
  wire [31:0] x407_rdcol_1_io_b; // @[Math.scala 150:24:@31188.4]
  wire  x407_rdcol_1_io_flow; // @[Math.scala 150:24:@31188.4]
  wire [31:0] x407_rdcol_1_io_result; // @[Math.scala 150:24:@31188.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@31209.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@31209.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@31209.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@31209.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@31209.4]
  wire  x411_sum_1_clock; // @[Math.scala 150:24:@31218.4]
  wire  x411_sum_1_reset; // @[Math.scala 150:24:@31218.4]
  wire [31:0] x411_sum_1_io_a; // @[Math.scala 150:24:@31218.4]
  wire [31:0] x411_sum_1_io_b; // @[Math.scala 150:24:@31218.4]
  wire  x411_sum_1_io_flow; // @[Math.scala 150:24:@31218.4]
  wire [31:0] x411_sum_1_io_result; // @[Math.scala 150:24:@31218.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@31228.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@31228.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@31228.4]
  wire [7:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@31228.4]
  wire [7:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@31228.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@31237.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@31237.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@31237.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@31237.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@31237.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@31250.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@31250.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@31250.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@31250.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@31250.4]
  wire  x416_rdcol_1_clock; // @[Math.scala 150:24:@31273.4]
  wire  x416_rdcol_1_reset; // @[Math.scala 150:24:@31273.4]
  wire [31:0] x416_rdcol_1_io_a; // @[Math.scala 150:24:@31273.4]
  wire [31:0] x416_rdcol_1_io_b; // @[Math.scala 150:24:@31273.4]
  wire  x416_rdcol_1_io_flow; // @[Math.scala 150:24:@31273.4]
  wire [31:0] x416_rdcol_1_io_result; // @[Math.scala 150:24:@31273.4]
  wire  x420_sum_1_clock; // @[Math.scala 150:24:@31294.4]
  wire  x420_sum_1_reset; // @[Math.scala 150:24:@31294.4]
  wire [31:0] x420_sum_1_io_a; // @[Math.scala 150:24:@31294.4]
  wire [31:0] x420_sum_1_io_b; // @[Math.scala 150:24:@31294.4]
  wire  x420_sum_1_io_flow; // @[Math.scala 150:24:@31294.4]
  wire [31:0] x420_sum_1_io_result; // @[Math.scala 150:24:@31294.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@31304.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@31304.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@31304.4]
  wire [7:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@31304.4]
  wire [7:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@31304.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@31313.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@31313.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@31313.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@31313.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@31313.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@31326.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@31326.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@31326.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@31326.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@31326.4]
  wire  x425_rdcol_1_clock; // @[Math.scala 150:24:@31349.4]
  wire  x425_rdcol_1_reset; // @[Math.scala 150:24:@31349.4]
  wire [31:0] x425_rdcol_1_io_a; // @[Math.scala 150:24:@31349.4]
  wire [31:0] x425_rdcol_1_io_b; // @[Math.scala 150:24:@31349.4]
  wire  x425_rdcol_1_io_flow; // @[Math.scala 150:24:@31349.4]
  wire [31:0] x425_rdcol_1_io_result; // @[Math.scala 150:24:@31349.4]
  wire  x429_sum_1_clock; // @[Math.scala 150:24:@31370.4]
  wire  x429_sum_1_reset; // @[Math.scala 150:24:@31370.4]
  wire [31:0] x429_sum_1_io_a; // @[Math.scala 150:24:@31370.4]
  wire [31:0] x429_sum_1_io_b; // @[Math.scala 150:24:@31370.4]
  wire  x429_sum_1_io_flow; // @[Math.scala 150:24:@31370.4]
  wire [31:0] x429_sum_1_io_result; // @[Math.scala 150:24:@31370.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@31380.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@31380.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@31380.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@31380.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@31380.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@31389.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@31389.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@31389.4]
  wire [7:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@31389.4]
  wire [7:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@31389.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@31402.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@31402.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@31402.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@31402.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@31402.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@31423.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@31423.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@31423.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@31423.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@31423.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@31450.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@31450.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@31450.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@31450.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@31450.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@31468.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@31468.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@31468.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@31468.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@31468.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@31503.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@31503.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@31503.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@31503.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@31503.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@31512.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@31512.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@31512.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@31512.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@31512.4]
  wire  x442_sum_1_clock; // @[Math.scala 150:24:@31521.4]
  wire  x442_sum_1_reset; // @[Math.scala 150:24:@31521.4]
  wire [31:0] x442_sum_1_io_a; // @[Math.scala 150:24:@31521.4]
  wire [31:0] x442_sum_1_io_b; // @[Math.scala 150:24:@31521.4]
  wire  x442_sum_1_io_flow; // @[Math.scala 150:24:@31521.4]
  wire [31:0] x442_sum_1_io_result; // @[Math.scala 150:24:@31521.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@31531.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@31531.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@31531.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@31531.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@31531.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@31540.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@31540.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@31540.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@31540.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@31540.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@31549.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@31549.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@31549.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@31549.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@31549.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@31558.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@31558.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@31558.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@31558.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@31558.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@31572.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@31572.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@31572.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@31572.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@31572.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@31593.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@31593.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@31593.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@31615.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@31615.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@31615.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@31615.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@31615.4]
  wire  x451_sum_1_clock; // @[Math.scala 150:24:@31624.4]
  wire  x451_sum_1_reset; // @[Math.scala 150:24:@31624.4]
  wire [31:0] x451_sum_1_io_a; // @[Math.scala 150:24:@31624.4]
  wire [31:0] x451_sum_1_io_b; // @[Math.scala 150:24:@31624.4]
  wire  x451_sum_1_io_flow; // @[Math.scala 150:24:@31624.4]
  wire [31:0] x451_sum_1_io_result; // @[Math.scala 150:24:@31624.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@31634.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@31634.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@31634.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@31634.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@31634.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@31648.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@31648.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@31648.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@31648.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@31648.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@31669.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@31669.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@31669.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@31669.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@31669.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@31691.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@31691.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@31691.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@31691.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@31691.4]
  wire  x459_sum_1_clock; // @[Math.scala 150:24:@31700.4]
  wire  x459_sum_1_reset; // @[Math.scala 150:24:@31700.4]
  wire [31:0] x459_sum_1_io_a; // @[Math.scala 150:24:@31700.4]
  wire [31:0] x459_sum_1_io_b; // @[Math.scala 150:24:@31700.4]
  wire  x459_sum_1_io_flow; // @[Math.scala 150:24:@31700.4]
  wire [31:0] x459_sum_1_io_result; // @[Math.scala 150:24:@31700.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@31710.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@31710.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@31710.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@31710.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@31710.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@31724.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@31724.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@31724.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@31724.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@31724.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@31745.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@31745.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@31745.4]
  wire [31:0] RetimeWrapper_35_io_in; // @[package.scala 93:22:@31745.4]
  wire [31:0] RetimeWrapper_35_io_out; // @[package.scala 93:22:@31745.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@31767.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@31767.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@31767.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@31767.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@31767.4]
  wire  x467_sum_1_clock; // @[Math.scala 150:24:@31776.4]
  wire  x467_sum_1_reset; // @[Math.scala 150:24:@31776.4]
  wire [31:0] x467_sum_1_io_a; // @[Math.scala 150:24:@31776.4]
  wire [31:0] x467_sum_1_io_b; // @[Math.scala 150:24:@31776.4]
  wire  x467_sum_1_io_flow; // @[Math.scala 150:24:@31776.4]
  wire [31:0] x467_sum_1_io_result; // @[Math.scala 150:24:@31776.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@31786.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@31786.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@31786.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@31786.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@31786.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@31795.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@31795.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@31795.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@31795.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@31795.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@31809.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@31809.4]
  wire  x472_rdcol_1_clock; // @[Math.scala 150:24:@31832.4]
  wire  x472_rdcol_1_reset; // @[Math.scala 150:24:@31832.4]
  wire [31:0] x472_rdcol_1_io_a; // @[Math.scala 150:24:@31832.4]
  wire [31:0] x472_rdcol_1_io_b; // @[Math.scala 150:24:@31832.4]
  wire  x472_rdcol_1_io_flow; // @[Math.scala 150:24:@31832.4]
  wire [31:0] x472_rdcol_1_io_result; // @[Math.scala 150:24:@31832.4]
  wire  x478_sum_1_clock; // @[Math.scala 150:24:@31864.4]
  wire  x478_sum_1_reset; // @[Math.scala 150:24:@31864.4]
  wire [31:0] x478_sum_1_io_a; // @[Math.scala 150:24:@31864.4]
  wire [31:0] x478_sum_1_io_b; // @[Math.scala 150:24:@31864.4]
  wire  x478_sum_1_io_flow; // @[Math.scala 150:24:@31864.4]
  wire [31:0] x478_sum_1_io_result; // @[Math.scala 150:24:@31864.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@31874.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@31874.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@31874.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@31874.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@31874.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@31888.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@31888.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@31888.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@31888.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@31888.4]
  wire  x484_rdcol_1_clock; // @[Math.scala 150:24:@31913.4]
  wire  x484_rdcol_1_reset; // @[Math.scala 150:24:@31913.4]
  wire [31:0] x484_rdcol_1_io_a; // @[Math.scala 150:24:@31913.4]
  wire [31:0] x484_rdcol_1_io_b; // @[Math.scala 150:24:@31913.4]
  wire  x484_rdcol_1_io_flow; // @[Math.scala 150:24:@31913.4]
  wire [31:0] x484_rdcol_1_io_result; // @[Math.scala 150:24:@31913.4]
  wire  x490_sum_1_clock; // @[Math.scala 150:24:@31945.4]
  wire  x490_sum_1_reset; // @[Math.scala 150:24:@31945.4]
  wire [31:0] x490_sum_1_io_a; // @[Math.scala 150:24:@31945.4]
  wire [31:0] x490_sum_1_io_b; // @[Math.scala 150:24:@31945.4]
  wire  x490_sum_1_io_flow; // @[Math.scala 150:24:@31945.4]
  wire [31:0] x490_sum_1_io_result; // @[Math.scala 150:24:@31945.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@31955.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@31955.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@31955.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@31955.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@31955.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@31969.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@31969.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@31969.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@31969.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@31969.4]
  wire  x496_rdrow_1_clock; // @[Math.scala 191:24:@31992.4]
  wire  x496_rdrow_1_reset; // @[Math.scala 191:24:@31992.4]
  wire [31:0] x496_rdrow_1_io_a; // @[Math.scala 191:24:@31992.4]
  wire [31:0] x496_rdrow_1_io_b; // @[Math.scala 191:24:@31992.4]
  wire  x496_rdrow_1_io_flow; // @[Math.scala 191:24:@31992.4]
  wire [31:0] x496_rdrow_1_io_result; // @[Math.scala 191:24:@31992.4]
  wire  x503_sum_1_clock; // @[Math.scala 150:24:@32046.4]
  wire  x503_sum_1_reset; // @[Math.scala 150:24:@32046.4]
  wire [31:0] x503_sum_1_io_a; // @[Math.scala 150:24:@32046.4]
  wire [31:0] x503_sum_1_io_b; // @[Math.scala 150:24:@32046.4]
  wire  x503_sum_1_io_flow; // @[Math.scala 150:24:@32046.4]
  wire [31:0] x503_sum_1_io_result; // @[Math.scala 150:24:@32046.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@32056.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@32056.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@32056.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@32056.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@32056.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@32065.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@32065.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@32065.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@32065.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@32065.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@32079.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@32079.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@32079.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@32079.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@32079.4]
  wire  x511_sum_1_clock; // @[Math.scala 150:24:@32106.4]
  wire  x511_sum_1_reset; // @[Math.scala 150:24:@32106.4]
  wire [31:0] x511_sum_1_io_a; // @[Math.scala 150:24:@32106.4]
  wire [31:0] x511_sum_1_io_b; // @[Math.scala 150:24:@32106.4]
  wire  x511_sum_1_io_flow; // @[Math.scala 150:24:@32106.4]
  wire [31:0] x511_sum_1_io_result; // @[Math.scala 150:24:@32106.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@32116.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@32116.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@32116.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@32116.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@32116.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@32130.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@32130.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@32130.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@32130.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@32130.4]
  wire  x518_sum_1_clock; // @[Math.scala 150:24:@32157.4]
  wire  x518_sum_1_reset; // @[Math.scala 150:24:@32157.4]
  wire [31:0] x518_sum_1_io_a; // @[Math.scala 150:24:@32157.4]
  wire [31:0] x518_sum_1_io_b; // @[Math.scala 150:24:@32157.4]
  wire  x518_sum_1_io_flow; // @[Math.scala 150:24:@32157.4]
  wire [31:0] x518_sum_1_io_result; // @[Math.scala 150:24:@32157.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@32167.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@32167.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@32167.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@32167.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@32167.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@32181.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@32181.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@32181.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@32181.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@32181.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@32202.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@32202.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@32202.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@32202.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@32202.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@32217.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@32217.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@32217.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@32217.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@32217.4]
  wire  x525_sum_1_clock; // @[Math.scala 150:24:@32226.4]
  wire  x525_sum_1_reset; // @[Math.scala 150:24:@32226.4]
  wire [31:0] x525_sum_1_io_a; // @[Math.scala 150:24:@32226.4]
  wire [31:0] x525_sum_1_io_b; // @[Math.scala 150:24:@32226.4]
  wire  x525_sum_1_io_flow; // @[Math.scala 150:24:@32226.4]
  wire [31:0] x525_sum_1_io_result; // @[Math.scala 150:24:@32226.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@32236.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@32236.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@32236.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@32236.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@32236.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@32250.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@32250.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@32250.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@32250.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@32250.4]
  wire  x532_sum_1_clock; // @[Math.scala 150:24:@32277.4]
  wire  x532_sum_1_reset; // @[Math.scala 150:24:@32277.4]
  wire [31:0] x532_sum_1_io_a; // @[Math.scala 150:24:@32277.4]
  wire [31:0] x532_sum_1_io_b; // @[Math.scala 150:24:@32277.4]
  wire  x532_sum_1_io_flow; // @[Math.scala 150:24:@32277.4]
  wire [31:0] x532_sum_1_io_result; // @[Math.scala 150:24:@32277.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@32287.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@32287.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@32287.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@32287.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@32287.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@32301.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@32301.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@32301.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@32301.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@32301.4]
  wire  x539_sum_1_clock; // @[Math.scala 150:24:@32330.4]
  wire  x539_sum_1_reset; // @[Math.scala 150:24:@32330.4]
  wire [31:0] x539_sum_1_io_a; // @[Math.scala 150:24:@32330.4]
  wire [31:0] x539_sum_1_io_b; // @[Math.scala 150:24:@32330.4]
  wire  x539_sum_1_io_flow; // @[Math.scala 150:24:@32330.4]
  wire [31:0] x539_sum_1_io_result; // @[Math.scala 150:24:@32330.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@32340.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@32340.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@32340.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@32340.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@32340.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@32354.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@32354.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@32354.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@32354.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@32354.4]
  wire  x544_rdrow_1_clock; // @[Math.scala 191:24:@32377.4]
  wire  x544_rdrow_1_reset; // @[Math.scala 191:24:@32377.4]
  wire [31:0] x544_rdrow_1_io_a; // @[Math.scala 191:24:@32377.4]
  wire [31:0] x544_rdrow_1_io_b; // @[Math.scala 191:24:@32377.4]
  wire  x544_rdrow_1_io_flow; // @[Math.scala 191:24:@32377.4]
  wire [31:0] x544_rdrow_1_io_result; // @[Math.scala 191:24:@32377.4]
  wire  x551_sum_1_clock; // @[Math.scala 150:24:@32431.4]
  wire  x551_sum_1_reset; // @[Math.scala 150:24:@32431.4]
  wire [31:0] x551_sum_1_io_a; // @[Math.scala 150:24:@32431.4]
  wire [31:0] x551_sum_1_io_b; // @[Math.scala 150:24:@32431.4]
  wire  x551_sum_1_io_flow; // @[Math.scala 150:24:@32431.4]
  wire [31:0] x551_sum_1_io_result; // @[Math.scala 150:24:@32431.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@32441.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@32441.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@32441.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@32441.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@32441.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@32450.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@32464.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@32464.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@32464.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@32464.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@32464.4]
  wire  x559_sum_1_clock; // @[Math.scala 150:24:@32491.4]
  wire  x559_sum_1_reset; // @[Math.scala 150:24:@32491.4]
  wire [31:0] x559_sum_1_io_a; // @[Math.scala 150:24:@32491.4]
  wire [31:0] x559_sum_1_io_b; // @[Math.scala 150:24:@32491.4]
  wire  x559_sum_1_io_flow; // @[Math.scala 150:24:@32491.4]
  wire [31:0] x559_sum_1_io_result; // @[Math.scala 150:24:@32491.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@32501.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@32501.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@32501.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@32501.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@32501.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@32515.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@32515.4]
  wire  x566_sum_1_clock; // @[Math.scala 150:24:@32542.4]
  wire  x566_sum_1_reset; // @[Math.scala 150:24:@32542.4]
  wire [31:0] x566_sum_1_io_a; // @[Math.scala 150:24:@32542.4]
  wire [31:0] x566_sum_1_io_b; // @[Math.scala 150:24:@32542.4]
  wire  x566_sum_1_io_flow; // @[Math.scala 150:24:@32542.4]
  wire [31:0] x566_sum_1_io_result; // @[Math.scala 150:24:@32542.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@32552.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@32552.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@32552.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@32552.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@32552.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@32566.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@32566.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@32566.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@32566.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@32566.4]
  wire  x573_sum_1_clock; // @[Math.scala 150:24:@32593.4]
  wire  x573_sum_1_reset; // @[Math.scala 150:24:@32593.4]
  wire [31:0] x573_sum_1_io_a; // @[Math.scala 150:24:@32593.4]
  wire [31:0] x573_sum_1_io_b; // @[Math.scala 150:24:@32593.4]
  wire  x573_sum_1_io_flow; // @[Math.scala 150:24:@32593.4]
  wire [31:0] x573_sum_1_io_result; // @[Math.scala 150:24:@32593.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@32603.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@32603.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@32603.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@32603.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@32603.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@32617.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@32617.4]
  wire  x580_sum_1_clock; // @[Math.scala 150:24:@32644.4]
  wire  x580_sum_1_reset; // @[Math.scala 150:24:@32644.4]
  wire [31:0] x580_sum_1_io_a; // @[Math.scala 150:24:@32644.4]
  wire [31:0] x580_sum_1_io_b; // @[Math.scala 150:24:@32644.4]
  wire  x580_sum_1_io_flow; // @[Math.scala 150:24:@32644.4]
  wire [31:0] x580_sum_1_io_result; // @[Math.scala 150:24:@32644.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@32654.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@32654.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@32654.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@32654.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@32654.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@32668.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@32668.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@32668.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@32668.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@32668.4]
  wire  x587_sum_1_clock; // @[Math.scala 150:24:@32695.4]
  wire  x587_sum_1_reset; // @[Math.scala 150:24:@32695.4]
  wire [31:0] x587_sum_1_io_a; // @[Math.scala 150:24:@32695.4]
  wire [31:0] x587_sum_1_io_b; // @[Math.scala 150:24:@32695.4]
  wire  x587_sum_1_io_flow; // @[Math.scala 150:24:@32695.4]
  wire [31:0] x587_sum_1_io_result; // @[Math.scala 150:24:@32695.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@32705.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@32705.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@32705.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@32705.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@32705.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@32719.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@32719.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@32719.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@32719.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@32719.4]
  wire  x597_x23_1_clock; // @[Math.scala 150:24:@32767.4]
  wire  x597_x23_1_reset; // @[Math.scala 150:24:@32767.4]
  wire [7:0] x597_x23_1_io_a; // @[Math.scala 150:24:@32767.4]
  wire [7:0] x597_x23_1_io_b; // @[Math.scala 150:24:@32767.4]
  wire  x597_x23_1_io_flow; // @[Math.scala 150:24:@32767.4]
  wire [7:0] x597_x23_1_io_result; // @[Math.scala 150:24:@32767.4]
  wire  x598_x24_1_clock; // @[Math.scala 150:24:@32777.4]
  wire  x598_x24_1_reset; // @[Math.scala 150:24:@32777.4]
  wire [7:0] x598_x24_1_io_a; // @[Math.scala 150:24:@32777.4]
  wire [7:0] x598_x24_1_io_b; // @[Math.scala 150:24:@32777.4]
  wire  x598_x24_1_io_flow; // @[Math.scala 150:24:@32777.4]
  wire [7:0] x598_x24_1_io_result; // @[Math.scala 150:24:@32777.4]
  wire  x599_x23_1_clock; // @[Math.scala 150:24:@32787.4]
  wire  x599_x23_1_reset; // @[Math.scala 150:24:@32787.4]
  wire [7:0] x599_x23_1_io_a; // @[Math.scala 150:24:@32787.4]
  wire [7:0] x599_x23_1_io_b; // @[Math.scala 150:24:@32787.4]
  wire  x599_x23_1_io_flow; // @[Math.scala 150:24:@32787.4]
  wire [7:0] x599_x23_1_io_result; // @[Math.scala 150:24:@32787.4]
  wire  x600_x24_1_clock; // @[Math.scala 150:24:@32797.4]
  wire  x600_x24_1_reset; // @[Math.scala 150:24:@32797.4]
  wire [7:0] x600_x24_1_io_a; // @[Math.scala 150:24:@32797.4]
  wire [7:0] x600_x24_1_io_b; // @[Math.scala 150:24:@32797.4]
  wire  x600_x24_1_io_flow; // @[Math.scala 150:24:@32797.4]
  wire [7:0] x600_x24_1_io_result; // @[Math.scala 150:24:@32797.4]
  wire [7:0] x601_x23_1_io_a; // @[Math.scala 150:24:@32807.4]
  wire [7:0] x601_x23_1_io_b; // @[Math.scala 150:24:@32807.4]
  wire [7:0] x601_x23_1_io_result; // @[Math.scala 150:24:@32807.4]
  wire [7:0] x602_x24_1_io_a; // @[Math.scala 150:24:@32817.4]
  wire [7:0] x602_x24_1_io_b; // @[Math.scala 150:24:@32817.4]
  wire [7:0] x602_x24_1_io_result; // @[Math.scala 150:24:@32817.4]
  wire [7:0] x603_x23_1_io_a; // @[Math.scala 150:24:@32827.4]
  wire [7:0] x603_x23_1_io_b; // @[Math.scala 150:24:@32827.4]
  wire [7:0] x603_x23_1_io_result; // @[Math.scala 150:24:@32827.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@32837.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@32837.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@32837.4]
  wire [7:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@32837.4]
  wire [7:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@32837.4]
  wire [7:0] x604_sum_1_io_a; // @[Math.scala 150:24:@32846.4]
  wire [7:0] x604_sum_1_io_b; // @[Math.scala 150:24:@32846.4]
  wire [7:0] x604_sum_1_io_result; // @[Math.scala 150:24:@32846.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@32860.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@32860.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@32860.4]
  wire [7:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@32860.4]
  wire [7:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@32860.4]
  wire  x611_x23_1_clock; // @[Math.scala 150:24:@32895.4]
  wire  x611_x23_1_reset; // @[Math.scala 150:24:@32895.4]
  wire [7:0] x611_x23_1_io_a; // @[Math.scala 150:24:@32895.4]
  wire [7:0] x611_x23_1_io_b; // @[Math.scala 150:24:@32895.4]
  wire  x611_x23_1_io_flow; // @[Math.scala 150:24:@32895.4]
  wire [7:0] x611_x23_1_io_result; // @[Math.scala 150:24:@32895.4]
  wire  x612_x24_1_clock; // @[Math.scala 150:24:@32905.4]
  wire  x612_x24_1_reset; // @[Math.scala 150:24:@32905.4]
  wire [7:0] x612_x24_1_io_a; // @[Math.scala 150:24:@32905.4]
  wire [7:0] x612_x24_1_io_b; // @[Math.scala 150:24:@32905.4]
  wire  x612_x24_1_io_flow; // @[Math.scala 150:24:@32905.4]
  wire [7:0] x612_x24_1_io_result; // @[Math.scala 150:24:@32905.4]
  wire  x613_x23_1_clock; // @[Math.scala 150:24:@32915.4]
  wire  x613_x23_1_reset; // @[Math.scala 150:24:@32915.4]
  wire [7:0] x613_x23_1_io_a; // @[Math.scala 150:24:@32915.4]
  wire [7:0] x613_x23_1_io_b; // @[Math.scala 150:24:@32915.4]
  wire  x613_x23_1_io_flow; // @[Math.scala 150:24:@32915.4]
  wire [7:0] x613_x23_1_io_result; // @[Math.scala 150:24:@32915.4]
  wire  x614_x24_1_clock; // @[Math.scala 150:24:@32925.4]
  wire  x614_x24_1_reset; // @[Math.scala 150:24:@32925.4]
  wire [7:0] x614_x24_1_io_a; // @[Math.scala 150:24:@32925.4]
  wire [7:0] x614_x24_1_io_b; // @[Math.scala 150:24:@32925.4]
  wire  x614_x24_1_io_flow; // @[Math.scala 150:24:@32925.4]
  wire [7:0] x614_x24_1_io_result; // @[Math.scala 150:24:@32925.4]
  wire [7:0] x615_x23_1_io_a; // @[Math.scala 150:24:@32935.4]
  wire [7:0] x615_x23_1_io_b; // @[Math.scala 150:24:@32935.4]
  wire [7:0] x615_x23_1_io_result; // @[Math.scala 150:24:@32935.4]
  wire [7:0] x616_x24_1_io_a; // @[Math.scala 150:24:@32945.4]
  wire [7:0] x616_x24_1_io_b; // @[Math.scala 150:24:@32945.4]
  wire [7:0] x616_x24_1_io_result; // @[Math.scala 150:24:@32945.4]
  wire [7:0] x617_x23_1_io_a; // @[Math.scala 150:24:@32955.4]
  wire [7:0] x617_x23_1_io_b; // @[Math.scala 150:24:@32955.4]
  wire [7:0] x617_x23_1_io_result; // @[Math.scala 150:24:@32955.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@32965.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@32965.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@32965.4]
  wire [7:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@32965.4]
  wire [7:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@32965.4]
  wire [7:0] x618_sum_1_io_a; // @[Math.scala 150:24:@32974.4]
  wire [7:0] x618_sum_1_io_b; // @[Math.scala 150:24:@32974.4]
  wire [7:0] x618_sum_1_io_result; // @[Math.scala 150:24:@32974.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@32988.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@32988.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@32988.4]
  wire [7:0] RetimeWrapper_75_io_in; // @[package.scala 93:22:@32988.4]
  wire [7:0] RetimeWrapper_75_io_out; // @[package.scala 93:22:@32988.4]
  wire  x624_x23_1_clock; // @[Math.scala 150:24:@33018.4]
  wire  x624_x23_1_reset; // @[Math.scala 150:24:@33018.4]
  wire [7:0] x624_x23_1_io_a; // @[Math.scala 150:24:@33018.4]
  wire [7:0] x624_x23_1_io_b; // @[Math.scala 150:24:@33018.4]
  wire  x624_x23_1_io_flow; // @[Math.scala 150:24:@33018.4]
  wire [7:0] x624_x23_1_io_result; // @[Math.scala 150:24:@33018.4]
  wire  x625_x24_1_clock; // @[Math.scala 150:24:@33028.4]
  wire  x625_x24_1_reset; // @[Math.scala 150:24:@33028.4]
  wire [7:0] x625_x24_1_io_a; // @[Math.scala 150:24:@33028.4]
  wire [7:0] x625_x24_1_io_b; // @[Math.scala 150:24:@33028.4]
  wire  x625_x24_1_io_flow; // @[Math.scala 150:24:@33028.4]
  wire [7:0] x625_x24_1_io_result; // @[Math.scala 150:24:@33028.4]
  wire  x626_x23_1_clock; // @[Math.scala 150:24:@33038.4]
  wire  x626_x23_1_reset; // @[Math.scala 150:24:@33038.4]
  wire [7:0] x626_x23_1_io_a; // @[Math.scala 150:24:@33038.4]
  wire [7:0] x626_x23_1_io_b; // @[Math.scala 150:24:@33038.4]
  wire  x626_x23_1_io_flow; // @[Math.scala 150:24:@33038.4]
  wire [7:0] x626_x23_1_io_result; // @[Math.scala 150:24:@33038.4]
  wire  x627_x24_1_clock; // @[Math.scala 150:24:@33048.4]
  wire  x627_x24_1_reset; // @[Math.scala 150:24:@33048.4]
  wire [7:0] x627_x24_1_io_a; // @[Math.scala 150:24:@33048.4]
  wire [7:0] x627_x24_1_io_b; // @[Math.scala 150:24:@33048.4]
  wire  x627_x24_1_io_flow; // @[Math.scala 150:24:@33048.4]
  wire [7:0] x627_x24_1_io_result; // @[Math.scala 150:24:@33048.4]
  wire [7:0] x628_x23_1_io_a; // @[Math.scala 150:24:@33058.4]
  wire [7:0] x628_x23_1_io_b; // @[Math.scala 150:24:@33058.4]
  wire [7:0] x628_x23_1_io_result; // @[Math.scala 150:24:@33058.4]
  wire [7:0] x629_x24_1_io_a; // @[Math.scala 150:24:@33068.4]
  wire [7:0] x629_x24_1_io_b; // @[Math.scala 150:24:@33068.4]
  wire [7:0] x629_x24_1_io_result; // @[Math.scala 150:24:@33068.4]
  wire [7:0] x630_x23_1_io_a; // @[Math.scala 150:24:@33078.4]
  wire [7:0] x630_x23_1_io_b; // @[Math.scala 150:24:@33078.4]
  wire [7:0] x630_x23_1_io_result; // @[Math.scala 150:24:@33078.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@33088.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@33088.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@33088.4]
  wire [7:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@33088.4]
  wire [7:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@33088.4]
  wire [7:0] x631_sum_1_io_a; // @[Math.scala 150:24:@33097.4]
  wire [7:0] x631_sum_1_io_b; // @[Math.scala 150:24:@33097.4]
  wire [7:0] x631_sum_1_io_result; // @[Math.scala 150:24:@33097.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@33111.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@33111.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@33111.4]
  wire [7:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@33111.4]
  wire [7:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@33111.4]
  wire  x637_x23_1_clock; // @[Math.scala 150:24:@33141.4]
  wire  x637_x23_1_reset; // @[Math.scala 150:24:@33141.4]
  wire [7:0] x637_x23_1_io_a; // @[Math.scala 150:24:@33141.4]
  wire [7:0] x637_x23_1_io_b; // @[Math.scala 150:24:@33141.4]
  wire  x637_x23_1_io_flow; // @[Math.scala 150:24:@33141.4]
  wire [7:0] x637_x23_1_io_result; // @[Math.scala 150:24:@33141.4]
  wire  x638_x24_1_clock; // @[Math.scala 150:24:@33153.4]
  wire  x638_x24_1_reset; // @[Math.scala 150:24:@33153.4]
  wire [7:0] x638_x24_1_io_a; // @[Math.scala 150:24:@33153.4]
  wire [7:0] x638_x24_1_io_b; // @[Math.scala 150:24:@33153.4]
  wire  x638_x24_1_io_flow; // @[Math.scala 150:24:@33153.4]
  wire [7:0] x638_x24_1_io_result; // @[Math.scala 150:24:@33153.4]
  wire  x639_x23_1_clock; // @[Math.scala 150:24:@33163.4]
  wire  x639_x23_1_reset; // @[Math.scala 150:24:@33163.4]
  wire [7:0] x639_x23_1_io_a; // @[Math.scala 150:24:@33163.4]
  wire [7:0] x639_x23_1_io_b; // @[Math.scala 150:24:@33163.4]
  wire  x639_x23_1_io_flow; // @[Math.scala 150:24:@33163.4]
  wire [7:0] x639_x23_1_io_result; // @[Math.scala 150:24:@33163.4]
  wire  x640_x24_1_clock; // @[Math.scala 150:24:@33173.4]
  wire  x640_x24_1_reset; // @[Math.scala 150:24:@33173.4]
  wire [7:0] x640_x24_1_io_a; // @[Math.scala 150:24:@33173.4]
  wire [7:0] x640_x24_1_io_b; // @[Math.scala 150:24:@33173.4]
  wire  x640_x24_1_io_flow; // @[Math.scala 150:24:@33173.4]
  wire [7:0] x640_x24_1_io_result; // @[Math.scala 150:24:@33173.4]
  wire [7:0] x641_x23_1_io_a; // @[Math.scala 150:24:@33183.4]
  wire [7:0] x641_x23_1_io_b; // @[Math.scala 150:24:@33183.4]
  wire [7:0] x641_x23_1_io_result; // @[Math.scala 150:24:@33183.4]
  wire [7:0] x642_x24_1_io_a; // @[Math.scala 150:24:@33193.4]
  wire [7:0] x642_x24_1_io_b; // @[Math.scala 150:24:@33193.4]
  wire [7:0] x642_x24_1_io_result; // @[Math.scala 150:24:@33193.4]
  wire [7:0] x643_x23_1_io_a; // @[Math.scala 150:24:@33203.4]
  wire [7:0] x643_x23_1_io_b; // @[Math.scala 150:24:@33203.4]
  wire [7:0] x643_x23_1_io_result; // @[Math.scala 150:24:@33203.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@33213.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@33213.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@33213.4]
  wire [7:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@33213.4]
  wire [7:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@33213.4]
  wire [7:0] x644_sum_1_io_a; // @[Math.scala 150:24:@33222.4]
  wire [7:0] x644_sum_1_io_b; // @[Math.scala 150:24:@33222.4]
  wire [7:0] x644_sum_1_io_result; // @[Math.scala 150:24:@33222.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@33236.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@33236.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@33236.4]
  wire [7:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@33236.4]
  wire [7:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@33236.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@33246.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@33246.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@33246.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@33246.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@33246.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@33255.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@33255.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@33255.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@33255.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@33255.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@33264.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@33264.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@33264.4]
  wire [31:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@33264.4]
  wire [31:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@33264.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@33273.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@33273.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@33273.4]
  wire [31:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@33273.4]
  wire [31:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@33273.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@33286.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@33286.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@33286.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@33286.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@33286.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@33307.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@33307.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@33307.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@33320.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@33341.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@33341.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@33341.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@33341.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@33341.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@33375.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@33375.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@33375.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@33375.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@33375.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@33388.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@33388.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@33388.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@33388.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@33388.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@33409.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@33409.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@33409.4]
  wire [31:0] RetimeWrapper_91_io_in; // @[package.scala 93:22:@33409.4]
  wire [31:0] RetimeWrapper_91_io_out; // @[package.scala 93:22:@33409.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@33418.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@33427.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@33427.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@33427.4]
  wire [31:0] RetimeWrapper_93_io_in; // @[package.scala 93:22:@33427.4]
  wire [31:0] RetimeWrapper_93_io_out; // @[package.scala 93:22:@33427.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@33441.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@33441.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@33441.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@33441.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@33441.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@33462.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@33462.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@33462.4]
  wire [31:0] RetimeWrapper_95_io_in; // @[package.scala 93:22:@33462.4]
  wire [31:0] RetimeWrapper_95_io_out; // @[package.scala 93:22:@33462.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@33471.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@33471.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@33471.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@33471.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@33471.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@33485.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@33485.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@33485.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@33485.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@33485.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@33506.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@33506.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@33506.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@33506.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@33506.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@33515.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@33515.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@33515.4]
  wire [31:0] RetimeWrapper_99_io_in; // @[package.scala 93:22:@33515.4]
  wire [31:0] RetimeWrapper_99_io_out; // @[package.scala 93:22:@33515.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@33529.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@33529.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@33529.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@33529.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@33529.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@33550.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@33550.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@33550.4]
  wire [31:0] RetimeWrapper_101_io_in; // @[package.scala 93:22:@33550.4]
  wire [31:0] RetimeWrapper_101_io_out; // @[package.scala 93:22:@33550.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@33559.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@33559.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@33559.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@33559.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@33559.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@33573.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@33573.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@33573.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@33573.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@33573.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@33594.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@33594.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@33594.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@33594.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@33594.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@33603.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@33603.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@33603.4]
  wire [31:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@33603.4]
  wire [31:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@33603.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@33617.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@33617.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@33617.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@33617.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@33617.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@33638.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@33638.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@33638.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@33638.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@33638.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@33647.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@33647.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@33647.4]
  wire [31:0] RetimeWrapper_108_io_in; // @[package.scala 93:22:@33647.4]
  wire [31:0] RetimeWrapper_108_io_out; // @[package.scala 93:22:@33647.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@33656.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@33656.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@33656.4]
  wire [31:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@33656.4]
  wire [31:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@33656.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@33670.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@33670.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@33670.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@33670.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@33670.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@33691.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@33691.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@33691.4]
  wire [31:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@33691.4]
  wire [31:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@33691.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@33700.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@33700.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@33700.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@33700.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@33700.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@33714.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@33714.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@33714.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@33714.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@33714.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@33735.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@33735.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@33735.4]
  wire [31:0] RetimeWrapper_114_io_in; // @[package.scala 93:22:@33735.4]
  wire [31:0] RetimeWrapper_114_io_out; // @[package.scala 93:22:@33735.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@33744.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@33744.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@33744.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@33744.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@33744.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@33758.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@33779.4]
  wire [31:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@33779.4]
  wire [31:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@33779.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@33788.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@33788.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@33788.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@33788.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@33788.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@33802.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@33802.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@33802.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@33802.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@33802.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@33823.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@33823.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@33823.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@33823.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@33823.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@33832.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@33832.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@33832.4]
  wire [31:0] RetimeWrapper_121_io_in; // @[package.scala 93:22:@33832.4]
  wire [31:0] RetimeWrapper_121_io_out; // @[package.scala 93:22:@33832.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@33846.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@33846.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@33846.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@33846.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@33846.4]
  wire [7:0] x674_x25_1_io_a; // @[Math.scala 150:24:@33879.4]
  wire [7:0] x674_x25_1_io_b; // @[Math.scala 150:24:@33879.4]
  wire [7:0] x674_x25_1_io_result; // @[Math.scala 150:24:@33879.4]
  wire [7:0] x675_x26_1_io_a; // @[Math.scala 150:24:@33889.4]
  wire [7:0] x675_x26_1_io_b; // @[Math.scala 150:24:@33889.4]
  wire [7:0] x675_x26_1_io_result; // @[Math.scala 150:24:@33889.4]
  wire [7:0] x676_sum_1_io_a; // @[Math.scala 150:24:@33899.4]
  wire [7:0] x676_sum_1_io_b; // @[Math.scala 150:24:@33899.4]
  wire [7:0] x676_sum_1_io_result; // @[Math.scala 150:24:@33899.4]
  wire  x677_div_1_clock; // @[Math.scala 327:24:@33911.4]
  wire  x677_div_1_reset; // @[Math.scala 327:24:@33911.4]
  wire [7:0] x677_div_1_io_a; // @[Math.scala 327:24:@33911.4]
  wire  x677_div_1_io_flow; // @[Math.scala 327:24:@33911.4]
  wire [7:0] x677_div_1_io_result; // @[Math.scala 327:24:@33911.4]
  wire [7:0] x680_x25_1_io_a; // @[Math.scala 150:24:@33931.4]
  wire [7:0] x680_x25_1_io_b; // @[Math.scala 150:24:@33931.4]
  wire [7:0] x680_x25_1_io_result; // @[Math.scala 150:24:@33931.4]
  wire [7:0] x681_x26_1_io_a; // @[Math.scala 150:24:@33941.4]
  wire [7:0] x681_x26_1_io_b; // @[Math.scala 150:24:@33941.4]
  wire [7:0] x681_x26_1_io_result; // @[Math.scala 150:24:@33941.4]
  wire [7:0] x682_sum_1_io_a; // @[Math.scala 150:24:@33951.4]
  wire [7:0] x682_sum_1_io_b; // @[Math.scala 150:24:@33951.4]
  wire [7:0] x682_sum_1_io_result; // @[Math.scala 150:24:@33951.4]
  wire  x683_div_1_clock; // @[Math.scala 327:24:@33963.4]
  wire  x683_div_1_reset; // @[Math.scala 327:24:@33963.4]
  wire [7:0] x683_div_1_io_a; // @[Math.scala 327:24:@33963.4]
  wire  x683_div_1_io_flow; // @[Math.scala 327:24:@33963.4]
  wire [7:0] x683_div_1_io_result; // @[Math.scala 327:24:@33963.4]
  wire [7:0] x686_x25_1_io_a; // @[Math.scala 150:24:@33983.4]
  wire [7:0] x686_x25_1_io_b; // @[Math.scala 150:24:@33983.4]
  wire [7:0] x686_x25_1_io_result; // @[Math.scala 150:24:@33983.4]
  wire [7:0] x687_x26_1_io_a; // @[Math.scala 150:24:@33993.4]
  wire [7:0] x687_x26_1_io_b; // @[Math.scala 150:24:@33993.4]
  wire [7:0] x687_x26_1_io_result; // @[Math.scala 150:24:@33993.4]
  wire [7:0] x688_sum_1_io_a; // @[Math.scala 150:24:@34003.4]
  wire [7:0] x688_sum_1_io_b; // @[Math.scala 150:24:@34003.4]
  wire [7:0] x688_sum_1_io_result; // @[Math.scala 150:24:@34003.4]
  wire  x689_div_1_clock; // @[Math.scala 327:24:@34015.4]
  wire  x689_div_1_reset; // @[Math.scala 327:24:@34015.4]
  wire [7:0] x689_div_1_io_a; // @[Math.scala 327:24:@34015.4]
  wire  x689_div_1_io_flow; // @[Math.scala 327:24:@34015.4]
  wire [7:0] x689_div_1_io_result; // @[Math.scala 327:24:@34015.4]
  wire [7:0] x692_x25_1_io_a; // @[Math.scala 150:24:@34035.4]
  wire [7:0] x692_x25_1_io_b; // @[Math.scala 150:24:@34035.4]
  wire [7:0] x692_x25_1_io_result; // @[Math.scala 150:24:@34035.4]
  wire [7:0] x693_x26_1_io_a; // @[Math.scala 150:24:@34045.4]
  wire [7:0] x693_x26_1_io_b; // @[Math.scala 150:24:@34045.4]
  wire [7:0] x693_x26_1_io_result; // @[Math.scala 150:24:@34045.4]
  wire [7:0] x694_sum_1_io_a; // @[Math.scala 150:24:@34055.4]
  wire [7:0] x694_sum_1_io_b; // @[Math.scala 150:24:@34055.4]
  wire [7:0] x694_sum_1_io_result; // @[Math.scala 150:24:@34055.4]
  wire  x695_div_1_clock; // @[Math.scala 327:24:@34067.4]
  wire  x695_div_1_reset; // @[Math.scala 327:24:@34067.4]
  wire [7:0] x695_div_1_io_a; // @[Math.scala 327:24:@34067.4]
  wire  x695_div_1_io_flow; // @[Math.scala 327:24:@34067.4]
  wire [7:0] x695_div_1_io_result; // @[Math.scala 327:24:@34067.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@34087.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@34087.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@34087.4]
  wire [31:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@34087.4]
  wire [31:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@34087.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@34096.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@34096.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@34096.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@34096.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@34096.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@34105.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@34114.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@34114.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@34114.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@34114.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@34114.4]
  wire  b384; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 62:18:@30749.4]
  wire  b385; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 63:18:@30750.4]
  wire  _T_207; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 69:30:@30994.4]
  wire  _T_208; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 69:37:@30995.4]
  wire  _T_212; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:76:@31000.4]
  wire  _T_213; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:62:@31001.4]
  wire  _T_215; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:101:@31002.4]
  wire [31:0] x775_x388_D1_0_number; // @[package.scala 96:25:@31011.4 package.scala 96:25:@31012.4]
  wire [31:0] b382_number; // @[Math.scala 712:22:@30734.4 Math.scala 713:14:@30735.4]
  wire [31:0] _T_247; // @[Math.scala 499:52:@31031.4]
  wire  x392; // @[Math.scala 499:44:@31039.4]
  wire  x393; // @[Math.scala 499:44:@31046.4]
  wire  x394; // @[Math.scala 499:44:@31053.4]
  wire [31:0] _T_294; // @[Mux.scala 19:72:@31065.4]
  wire [31:0] _T_296; // @[Mux.scala 19:72:@31066.4]
  wire [31:0] _T_298; // @[Mux.scala 19:72:@31067.4]
  wire [31:0] _T_300; // @[Mux.scala 19:72:@31069.4]
  wire [31:0] x395_number; // @[Mux.scala 19:72:@31070.4]
  wire [31:0] _T_312; // @[Math.scala 406:49:@31080.4]
  wire [31:0] _T_314; // @[Math.scala 406:56:@31082.4]
  wire [31:0] _T_315; // @[Math.scala 406:56:@31083.4]
  wire  _T_320; // @[FixedPoint.scala 50:25:@31089.4]
  wire [1:0] _T_324; // @[Bitwise.scala 72:12:@31091.4]
  wire [29:0] _T_325; // @[FixedPoint.scala 18:52:@31092.4]
  wire [31:0] b383_number; // @[Math.scala 712:22:@30746.4 Math.scala 713:14:@30747.4]
  wire  _T_330; // @[FixedPoint.scala 50:25:@31098.4]
  wire [1:0] _T_334; // @[Bitwise.scala 72:12:@31100.4]
  wire [29:0] _T_335; // @[FixedPoint.scala 18:52:@31101.4]
  wire  _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:101:@31162.4]
  wire  _T_364; // @[package.scala 96:25:@31170.4 package.scala 96:25:@31171.4]
  wire  _T_366; // @[implicits.scala 55:10:@31172.4]
  wire  _T_367; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:118:@31173.4]
  wire  _T_369; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:205:@31175.4]
  wire  _T_370; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:224:@31176.4]
  wire  x777_b384_D4; // @[package.scala 96:25:@31130.4 package.scala 96:25:@31131.4]
  wire  _T_371; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:250:@31177.4]
  wire  x776_b385_D4; // @[package.scala 96:25:@31121.4 package.scala 96:25:@31122.4]
  wire [31:0] x407_rdcol_number; // @[Math.scala 154:22:@31194.4 Math.scala 155:14:@31195.4]
  wire  _T_384; // @[FixedPoint.scala 50:25:@31201.4]
  wire [1:0] _T_388; // @[Bitwise.scala 72:12:@31203.4]
  wire [29:0] _T_389; // @[FixedPoint.scala 18:52:@31204.4]
  wire  _T_412; // @[package.scala 96:25:@31255.4 package.scala 96:25:@31256.4]
  wire  _T_414; // @[implicits.scala 55:10:@31257.4]
  wire  _T_415; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:118:@31258.4]
  wire  _T_417; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:205:@31260.4]
  wire  _T_418; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:224:@31261.4]
  wire  _T_419; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:250:@31262.4]
  wire [31:0] x416_rdcol_number; // @[Math.scala 154:22:@31279.4 Math.scala 155:14:@31280.4]
  wire  _T_432; // @[FixedPoint.scala 50:25:@31286.4]
  wire [1:0] _T_436; // @[Bitwise.scala 72:12:@31288.4]
  wire [29:0] _T_437; // @[FixedPoint.scala 18:52:@31289.4]
  wire  _T_457; // @[package.scala 96:25:@31331.4 package.scala 96:25:@31332.4]
  wire  _T_459; // @[implicits.scala 55:10:@31333.4]
  wire  _T_460; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:118:@31334.4]
  wire  _T_462; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:205:@31336.4]
  wire  _T_463; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:224:@31337.4]
  wire  _T_464; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:250:@31338.4]
  wire [31:0] x425_rdcol_number; // @[Math.scala 154:22:@31355.4 Math.scala 155:14:@31356.4]
  wire  _T_477; // @[FixedPoint.scala 50:25:@31362.4]
  wire [1:0] _T_481; // @[Bitwise.scala 72:12:@31364.4]
  wire [29:0] _T_482; // @[FixedPoint.scala 18:52:@31365.4]
  wire  _T_502; // @[package.scala 96:25:@31407.4 package.scala 96:25:@31408.4]
  wire  _T_504; // @[implicits.scala 55:10:@31409.4]
  wire  _T_505; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:118:@31410.4]
  wire  _T_507; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:205:@31412.4]
  wire  _T_508; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:224:@31413.4]
  wire  _T_509; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:250:@31414.4]
  wire [31:0] x788_b382_D6_number; // @[package.scala 96:25:@31428.4 package.scala 96:25:@31429.4]
  wire [31:0] _T_521; // @[Math.scala 406:49:@31435.4]
  wire [31:0] _T_523; // @[Math.scala 406:56:@31437.4]
  wire [31:0] _T_524; // @[Math.scala 406:56:@31438.4]
  wire [31:0] x769_number; // @[implicits.scala 133:21:@31439.4]
  wire  x436; // @[Math.scala 465:44:@31447.4]
  wire [31:0] x789_x425_rdcol_D6_number; // @[package.scala 96:25:@31455.4 package.scala 96:25:@31456.4]
  wire [31:0] _T_544; // @[Math.scala 465:37:@31463.4]
  wire  x437; // @[Math.scala 465:44:@31465.4]
  wire  x790_x436_D1; // @[package.scala 96:25:@31473.4 package.scala 96:25:@31474.4]
  wire  x438; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 190:24:@31477.4]
  wire [31:0] _T_561; // @[Math.scala 406:49:@31486.4]
  wire [31:0] _T_563; // @[Math.scala 406:56:@31488.4]
  wire [31:0] _T_564; // @[Math.scala 406:56:@31489.4]
  wire  _T_569; // @[FixedPoint.scala 50:25:@31495.4]
  wire [1:0] _T_573; // @[Bitwise.scala 72:12:@31497.4]
  wire [29:0] _T_574; // @[FixedPoint.scala 18:52:@31498.4]
  wire  _T_612; // @[package.scala 96:25:@31577.4 package.scala 96:25:@31578.4]
  wire  _T_614; // @[implicits.scala 55:10:@31579.4]
  wire  _T_615; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 215:194:@31580.4]
  wire  x796_x439_D1; // @[package.scala 96:25:@31563.4 package.scala 96:25:@31564.4]
  wire  _T_616; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 215:281:@31581.4]
  wire  x794_b384_D8; // @[package.scala 96:25:@31545.4 package.scala 96:25:@31546.4]
  wire  _T_617; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 215:289:@31582.4]
  wire  x793_b385_D8; // @[package.scala 96:25:@31536.4 package.scala 96:25:@31537.4]
  wire [31:0] x797_x416_rdcol_D6_number; // @[package.scala 96:25:@31598.4 package.scala 96:25:@31599.4]
  wire [31:0] _T_628; // @[Math.scala 465:37:@31604.4]
  wire  x448; // @[Math.scala 465:44:@31606.4]
  wire  x449; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 223:24:@31609.4]
  wire  _T_659; // @[package.scala 96:25:@31653.4 package.scala 96:25:@31654.4]
  wire  _T_661; // @[implicits.scala 55:10:@31655.4]
  wire  _T_662; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:194:@31656.4]
  wire  x799_x450_D1; // @[package.scala 96:25:@31639.4 package.scala 96:25:@31640.4]
  wire  _T_663; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:281:@31657.4]
  wire  _T_664; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:289:@31658.4]
  wire [31:0] x800_x407_rdcol_D6_number; // @[package.scala 96:25:@31674.4 package.scala 96:25:@31675.4]
  wire [31:0] _T_675; // @[Math.scala 465:37:@31680.4]
  wire  x456; // @[Math.scala 465:44:@31682.4]
  wire  x457; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 244:24:@31685.4]
  wire  _T_706; // @[package.scala 96:25:@31729.4 package.scala 96:25:@31730.4]
  wire  _T_708; // @[implicits.scala 55:10:@31731.4]
  wire  _T_709; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:194:@31732.4]
  wire  x802_x458_D1; // @[package.scala 96:25:@31715.4 package.scala 96:25:@31716.4]
  wire  _T_710; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:281:@31733.4]
  wire  _T_711; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:289:@31734.4]
  wire [31:0] x803_b383_D6_number; // @[package.scala 96:25:@31750.4 package.scala 96:25:@31751.4]
  wire [31:0] _T_722; // @[Math.scala 465:37:@31756.4]
  wire  x464; // @[Math.scala 465:44:@31758.4]
  wire  x465; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 265:59:@31761.4]
  wire  _T_756; // @[package.scala 96:25:@31814.4 package.scala 96:25:@31815.4]
  wire  _T_758; // @[implicits.scala 55:10:@31816.4]
  wire  _T_759; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:194:@31817.4]
  wire  x806_x466_D2; // @[package.scala 96:25:@31800.4 package.scala 96:25:@31801.4]
  wire  _T_760; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:281:@31818.4]
  wire  _T_761; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:289:@31819.4]
  wire [31:0] x472_rdcol_number; // @[Math.scala 154:22:@31838.4 Math.scala 155:14:@31839.4]
  wire [31:0] _T_776; // @[Math.scala 465:37:@31844.4]
  wire  x473; // @[Math.scala 465:44:@31846.4]
  wire  x474; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 288:24:@31849.4]
  wire  _T_786; // @[FixedPoint.scala 50:25:@31856.4]
  wire [1:0] _T_790; // @[Bitwise.scala 72:12:@31858.4]
  wire [29:0] _T_791; // @[FixedPoint.scala 18:52:@31859.4]
  wire  _T_814; // @[package.scala 96:25:@31893.4 package.scala 96:25:@31894.4]
  wire  _T_816; // @[implicits.scala 55:10:@31895.4]
  wire  _T_817; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:194:@31896.4]
  wire  x807_x475_D1; // @[package.scala 96:25:@31879.4 package.scala 96:25:@31880.4]
  wire  _T_818; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:281:@31897.4]
  wire  _T_819; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:289:@31898.4]
  wire [31:0] x484_rdcol_number; // @[Math.scala 154:22:@31919.4 Math.scala 155:14:@31920.4]
  wire [31:0] _T_836; // @[Math.scala 465:37:@31925.4]
  wire  x485; // @[Math.scala 465:44:@31927.4]
  wire  x486; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 317:59:@31930.4]
  wire  _T_846; // @[FixedPoint.scala 50:25:@31937.4]
  wire [1:0] _T_850; // @[Bitwise.scala 72:12:@31939.4]
  wire [29:0] _T_851; // @[FixedPoint.scala 18:52:@31940.4]
  wire  _T_874; // @[package.scala 96:25:@31974.4 package.scala 96:25:@31975.4]
  wire  _T_876; // @[implicits.scala 55:10:@31976.4]
  wire  _T_877; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 330:194:@31977.4]
  wire  x808_x487_D1; // @[package.scala 96:25:@31960.4 package.scala 96:25:@31961.4]
  wire  _T_878; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 330:281:@31978.4]
  wire  _T_879; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 330:289:@31979.4]
  wire [31:0] x496_rdrow_number; // @[Math.scala 195:22:@31998.4 Math.scala 196:14:@31999.4]
  wire [31:0] _T_896; // @[Math.scala 406:49:@32005.4]
  wire [31:0] _T_898; // @[Math.scala 406:56:@32007.4]
  wire [31:0] _T_899; // @[Math.scala 406:56:@32008.4]
  wire [31:0] x771_number; // @[implicits.scala 133:21:@32009.4]
  wire  x498; // @[Math.scala 465:44:@32017.4]
  wire  x499; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 340:24:@32020.4]
  wire [31:0] _T_920; // @[Math.scala 406:49:@32029.4]
  wire [31:0] _T_922; // @[Math.scala 406:56:@32031.4]
  wire [31:0] _T_923; // @[Math.scala 406:56:@32032.4]
  wire  _T_928; // @[FixedPoint.scala 50:25:@32038.4]
  wire [1:0] _T_932; // @[Bitwise.scala 72:12:@32040.4]
  wire [29:0] _T_933; // @[FixedPoint.scala 18:52:@32041.4]
  wire  _T_959; // @[package.scala 96:25:@32084.4 package.scala 96:25:@32085.4]
  wire  _T_961; // @[implicits.scala 55:10:@32086.4]
  wire  _T_962; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:194:@32087.4]
  wire  x809_x500_D1; // @[package.scala 96:25:@32061.4 package.scala 96:25:@32062.4]
  wire  _T_963; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:281:@32088.4]
  wire  _T_964; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:289:@32089.4]
  wire  x509; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 361:24:@32100.4]
  wire  _T_992; // @[package.scala 96:25:@32135.4 package.scala 96:25:@32136.4]
  wire  _T_994; // @[implicits.scala 55:10:@32137.4]
  wire  _T_995; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:194:@32138.4]
  wire  x811_x510_D1; // @[package.scala 96:25:@32121.4 package.scala 96:25:@32122.4]
  wire  _T_996; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:281:@32139.4]
  wire  _T_997; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:289:@32140.4]
  wire  x516; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 376:24:@32151.4]
  wire  _T_1025; // @[package.scala 96:25:@32186.4 package.scala 96:25:@32187.4]
  wire  _T_1027; // @[implicits.scala 55:10:@32188.4]
  wire  _T_1028; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:194:@32189.4]
  wire  x812_x517_D1; // @[package.scala 96:25:@32172.4 package.scala 96:25:@32173.4]
  wire  _T_1029; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:281:@32190.4]
  wire  _T_1030; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:289:@32191.4]
  wire  x813_x464_D1; // @[package.scala 96:25:@32207.4 package.scala 96:25:@32208.4]
  wire  x523; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 393:24:@32211.4]
  wire  _T_1064; // @[package.scala 96:25:@32255.4 package.scala 96:25:@32256.4]
  wire  _T_1066; // @[implicits.scala 55:10:@32257.4]
  wire  _T_1067; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:194:@32258.4]
  wire  x815_x524_D1; // @[package.scala 96:25:@32241.4 package.scala 96:25:@32242.4]
  wire  _T_1068; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:281:@32259.4]
  wire  _T_1069; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:289:@32260.4]
  wire  x530; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 410:24:@32271.4]
  wire  _T_1097; // @[package.scala 96:25:@32306.4 package.scala 96:25:@32307.4]
  wire  _T_1099; // @[implicits.scala 55:10:@32308.4]
  wire  _T_1100; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:194:@32309.4]
  wire  x816_x531_D1; // @[package.scala 96:25:@32292.4 package.scala 96:25:@32293.4]
  wire  _T_1101; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:281:@32310.4]
  wire  _T_1102; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:289:@32311.4]
  wire  x537; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 431:59:@32322.4]
  wire  _T_1132; // @[package.scala 96:25:@32359.4 package.scala 96:25:@32360.4]
  wire  _T_1134; // @[implicits.scala 55:10:@32361.4]
  wire  _T_1135; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:194:@32362.4]
  wire  x817_x538_D1; // @[package.scala 96:25:@32345.4 package.scala 96:25:@32346.4]
  wire  _T_1136; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:281:@32363.4]
  wire  _T_1137; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:289:@32364.4]
  wire [31:0] x544_rdrow_number; // @[Math.scala 195:22:@32383.4 Math.scala 196:14:@32384.4]
  wire [31:0] _T_1154; // @[Math.scala 406:49:@32390.4]
  wire [31:0] _T_1156; // @[Math.scala 406:56:@32392.4]
  wire [31:0] _T_1157; // @[Math.scala 406:56:@32393.4]
  wire [31:0] x773_number; // @[implicits.scala 133:21:@32394.4]
  wire  x546; // @[Math.scala 465:44:@32402.4]
  wire  x547; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 454:24:@32405.4]
  wire [31:0] _T_1178; // @[Math.scala 406:49:@32414.4]
  wire [31:0] _T_1180; // @[Math.scala 406:56:@32416.4]
  wire [31:0] _T_1181; // @[Math.scala 406:56:@32417.4]
  wire  _T_1186; // @[FixedPoint.scala 50:25:@32423.4]
  wire [1:0] _T_1190; // @[Bitwise.scala 72:12:@32425.4]
  wire [29:0] _T_1191; // @[FixedPoint.scala 18:52:@32426.4]
  wire  _T_1217; // @[package.scala 96:25:@32469.4 package.scala 96:25:@32470.4]
  wire  _T_1219; // @[implicits.scala 55:10:@32471.4]
  wire  _T_1220; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 471:194:@32472.4]
  wire  x819_x548_D1; // @[package.scala 96:25:@32455.4 package.scala 96:25:@32456.4]
  wire  _T_1221; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 471:281:@32473.4]
  wire  _T_1222; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 471:289:@32474.4]
  wire  x557; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 475:24:@32485.4]
  wire  _T_1250; // @[package.scala 96:25:@32520.4 package.scala 96:25:@32521.4]
  wire  _T_1252; // @[implicits.scala 55:10:@32522.4]
  wire  _T_1253; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:194:@32523.4]
  wire  x820_x558_D1; // @[package.scala 96:25:@32506.4 package.scala 96:25:@32507.4]
  wire  _T_1254; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:281:@32524.4]
  wire  _T_1255; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:289:@32525.4]
  wire  x564; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 490:24:@32536.4]
  wire  _T_1283; // @[package.scala 96:25:@32571.4 package.scala 96:25:@32572.4]
  wire  _T_1285; // @[implicits.scala 55:10:@32573.4]
  wire  _T_1286; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:194:@32574.4]
  wire  x821_x565_D1; // @[package.scala 96:25:@32557.4 package.scala 96:25:@32558.4]
  wire  _T_1287; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:281:@32575.4]
  wire  _T_1288; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:289:@32576.4]
  wire  x571; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 505:24:@32587.4]
  wire  _T_1316; // @[package.scala 96:25:@32622.4 package.scala 96:25:@32623.4]
  wire  _T_1318; // @[implicits.scala 55:10:@32624.4]
  wire  _T_1319; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:194:@32625.4]
  wire  x822_x572_D1; // @[package.scala 96:25:@32608.4 package.scala 96:25:@32609.4]
  wire  _T_1320; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:281:@32626.4]
  wire  _T_1321; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:289:@32627.4]
  wire  x578; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 520:24:@32638.4]
  wire  _T_1349; // @[package.scala 96:25:@32673.4 package.scala 96:25:@32674.4]
  wire  _T_1351; // @[implicits.scala 55:10:@32675.4]
  wire  _T_1352; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:194:@32676.4]
  wire  x823_x579_D1; // @[package.scala 96:25:@32659.4 package.scala 96:25:@32660.4]
  wire  _T_1353; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:281:@32677.4]
  wire  _T_1354; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:289:@32678.4]
  wire  x585; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 535:24:@32689.4]
  wire  _T_1382; // @[package.scala 96:25:@32724.4 package.scala 96:25:@32725.4]
  wire  _T_1384; // @[implicits.scala 55:10:@32726.4]
  wire  _T_1385; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 546:194:@32727.4]
  wire  x824_x586_D1; // @[package.scala 96:25:@32710.4 package.scala 96:25:@32711.4]
  wire  _T_1386; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 546:281:@32728.4]
  wire  _T_1387; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 546:289:@32729.4]
  wire [7:0] x454_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 232:29:@31642.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:336:@31665.4]
  wire [8:0] _GEN_0; // @[Math.scala 450:32:@32743.4]
  wire [8:0] _T_1395; // @[Math.scala 450:32:@32743.4]
  wire [7:0] x507_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 353:29:@32073.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:406:@32096.4]
  wire [8:0] _GEN_1; // @[Math.scala 450:32:@32748.4]
  wire [8:0] _T_1399; // @[Math.scala 450:32:@32748.4]
  wire [7:0] x514_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 368:29:@32124.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:406:@32147.4]
  wire [9:0] _GEN_2; // @[Math.scala 450:32:@32753.4]
  wire [9:0] _T_1403; // @[Math.scala 450:32:@32753.4]
  wire [7:0] x521_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 383:29:@32175.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:406:@32198.4]
  wire [8:0] _GEN_3; // @[Math.scala 450:32:@32758.4]
  wire [8:0] _T_1407; // @[Math.scala 450:32:@32758.4]
  wire [7:0] x562_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 482:29:@32509.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:406:@32532.4]
  wire [8:0] _GEN_4; // @[Math.scala 450:32:@32763.4]
  wire [8:0] _T_1411; // @[Math.scala 450:32:@32763.4]
  wire [7:0] x604_sum_number; // @[Math.scala 154:22:@32852.4 Math.scala 155:14:@32853.4]
  wire [3:0] _T_1447; // @[FixedPoint.scala 18:52:@32858.4]
  wire [7:0] x462_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 253:29:@31718.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:336:@31741.4]
  wire [8:0] _GEN_5; // @[Math.scala 450:32:@32871.4]
  wire [8:0] _T_1454; // @[Math.scala 450:32:@32871.4]
  wire [8:0] _GEN_6; // @[Math.scala 450:32:@32876.4]
  wire [8:0] _T_1458; // @[Math.scala 450:32:@32876.4]
  wire [9:0] _GEN_7; // @[Math.scala 450:32:@32881.4]
  wire [9:0] _T_1462; // @[Math.scala 450:32:@32881.4]
  wire [7:0] x528_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 402:29:@32244.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:406:@32267.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@32886.4]
  wire [8:0] _T_1466; // @[Math.scala 450:32:@32886.4]
  wire [7:0] x569_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 497:29:@32560.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:406:@32583.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@32891.4]
  wire [8:0] _T_1470; // @[Math.scala 450:32:@32891.4]
  wire [7:0] x618_sum_number; // @[Math.scala 154:22:@32980.4 Math.scala 155:14:@32981.4]
  wire [3:0] _T_1506; // @[FixedPoint.scala 18:52:@32986.4]
  wire [7:0] x470_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 276:29:@31803.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:336:@31826.4]
  wire [8:0] _GEN_10; // @[Math.scala 450:32:@32999.4]
  wire [8:0] _T_1513; // @[Math.scala 450:32:@32999.4]
  wire [9:0] _GEN_11; // @[Math.scala 450:32:@33004.4]
  wire [9:0] _T_1517; // @[Math.scala 450:32:@33004.4]
  wire [7:0] x535_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 417:29:@32295.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:406:@32318.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@33009.4]
  wire [8:0] _T_1521; // @[Math.scala 450:32:@33009.4]
  wire [7:0] x576_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 512:29:@32611.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:406:@32634.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@33014.4]
  wire [8:0] _T_1525; // @[Math.scala 450:32:@33014.4]
  wire [7:0] x631_sum_number; // @[Math.scala 154:22:@33103.4 Math.scala 155:14:@33104.4]
  wire [3:0] _T_1561; // @[FixedPoint.scala 18:52:@33109.4]
  wire [7:0] x482_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 303:29:@31882.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:406:@31905.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@33122.4]
  wire [8:0] _T_1568; // @[Math.scala 450:32:@33122.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@33127.4]
  wire [9:0] _T_1572; // @[Math.scala 450:32:@33127.4]
  wire [7:0] x542_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 440:29:@32348.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:406:@32371.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@33132.4]
  wire [8:0] _T_1576; // @[Math.scala 450:32:@33132.4]
  wire [7:0] x583_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 527:29:@32662.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:406:@32685.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@33137.4]
  wire [8:0] _T_1580; // @[Math.scala 450:32:@33137.4]
  wire [7:0] x644_sum_number; // @[Math.scala 154:22:@33228.4 Math.scala 155:14:@33229.4]
  wire [3:0] _T_1618; // @[FixedPoint.scala 18:52:@33234.4]
  wire  _T_1643; // @[package.scala 96:25:@33291.4 package.scala 96:25:@33292.4]
  wire  _T_1645; // @[implicits.scala 55:10:@33293.4]
  wire  _T_1646; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:167:@33294.4]
  wire  _T_1648; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:255:@33296.4]
  wire  _T_1649; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:274:@33297.4]
  wire  x830_b384_D12; // @[package.scala 96:25:@33260.4 package.scala 96:25:@33261.4]
  wire  _T_1650; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:300:@33298.4]
  wire  x829_b385_D12; // @[package.scala 96:25:@33251.4 package.scala 96:25:@33252.4]
  wire  _T_1664; // @[package.scala 96:25:@33325.4 package.scala 96:25:@33326.4]
  wire  _T_1666; // @[implicits.scala 55:10:@33327.4]
  wire  _T_1667; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:167:@33328.4]
  wire  _T_1669; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:255:@33330.4]
  wire  _T_1670; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:274:@33331.4]
  wire  _T_1671; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:300:@33332.4]
  wire  _T_1685; // @[package.scala 96:25:@33359.4 package.scala 96:25:@33360.4]
  wire  _T_1687; // @[implicits.scala 55:10:@33361.4]
  wire  _T_1688; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:167:@33362.4]
  wire  _T_1690; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:255:@33364.4]
  wire  _T_1691; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:274:@33365.4]
  wire  _T_1692; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:300:@33366.4]
  wire  _T_1706; // @[package.scala 96:25:@33393.4 package.scala 96:25:@33394.4]
  wire  _T_1708; // @[implicits.scala 55:10:@33395.4]
  wire  _T_1709; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:167:@33396.4]
  wire  _T_1711; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:255:@33398.4]
  wire  _T_1712; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:274:@33399.4]
  wire  _T_1713; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:300:@33400.4]
  wire  _T_1739; // @[package.scala 96:25:@33446.4 package.scala 96:25:@33447.4]
  wire  _T_1741; // @[implicits.scala 55:10:@33448.4]
  wire  _T_1742; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 727:195:@33449.4]
  wire  x837_x439_D5; // @[package.scala 96:25:@33423.4 package.scala 96:25:@33424.4]
  wire  _T_1743; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 727:283:@33450.4]
  wire  _T_1744; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 727:291:@33451.4]
  wire  _T_1768; // @[package.scala 96:25:@33490.4 package.scala 96:25:@33491.4]
  wire  _T_1770; // @[implicits.scala 55:10:@33492.4]
  wire  _T_1771; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:195:@33493.4]
  wire  x840_x450_D5; // @[package.scala 96:25:@33476.4 package.scala 96:25:@33477.4]
  wire  _T_1772; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:283:@33494.4]
  wire  _T_1773; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:291:@33495.4]
  wire  _T_1797; // @[package.scala 96:25:@33534.4 package.scala 96:25:@33535.4]
  wire  _T_1799; // @[implicits.scala 55:10:@33536.4]
  wire  _T_1800; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:195:@33537.4]
  wire  x841_x458_D5; // @[package.scala 96:25:@33511.4 package.scala 96:25:@33512.4]
  wire  _T_1801; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:283:@33538.4]
  wire  _T_1802; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:291:@33539.4]
  wire  _T_1826; // @[package.scala 96:25:@33578.4 package.scala 96:25:@33579.4]
  wire  _T_1828; // @[implicits.scala 55:10:@33580.4]
  wire  _T_1829; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:195:@33581.4]
  wire  x844_x466_D6; // @[package.scala 96:25:@33564.4 package.scala 96:25:@33565.4]
  wire  _T_1830; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:283:@33582.4]
  wire  _T_1831; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:291:@33583.4]
  wire  _T_1855; // @[package.scala 96:25:@33622.4 package.scala 96:25:@33623.4]
  wire  _T_1857; // @[implicits.scala 55:10:@33624.4]
  wire  _T_1858; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:195:@33625.4]
  wire  x845_x475_D5; // @[package.scala 96:25:@33599.4 package.scala 96:25:@33600.4]
  wire  _T_1859; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:283:@33626.4]
  wire  _T_1860; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:291:@33627.4]
  wire  _T_1887; // @[package.scala 96:25:@33675.4 package.scala 96:25:@33676.4]
  wire  _T_1889; // @[implicits.scala 55:10:@33677.4]
  wire  _T_1890; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:195:@33678.4]
  wire  x847_x500_D5; // @[package.scala 96:25:@33643.4 package.scala 96:25:@33644.4]
  wire  _T_1891; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:283:@33679.4]
  wire  _T_1892; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:291:@33680.4]
  wire  _T_1916; // @[package.scala 96:25:@33719.4 package.scala 96:25:@33720.4]
  wire  _T_1918; // @[implicits.scala 55:10:@33721.4]
  wire  _T_1919; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:195:@33722.4]
  wire  x851_x510_D5; // @[package.scala 96:25:@33705.4 package.scala 96:25:@33706.4]
  wire  _T_1920; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:283:@33723.4]
  wire  _T_1921; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:291:@33724.4]
  wire  _T_1945; // @[package.scala 96:25:@33763.4 package.scala 96:25:@33764.4]
  wire  _T_1947; // @[implicits.scala 55:10:@33765.4]
  wire  _T_1948; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:195:@33766.4]
  wire  x853_x517_D5; // @[package.scala 96:25:@33749.4 package.scala 96:25:@33750.4]
  wire  _T_1949; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:283:@33767.4]
  wire  _T_1950; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:291:@33768.4]
  wire  _T_1974; // @[package.scala 96:25:@33807.4 package.scala 96:25:@33808.4]
  wire  _T_1976; // @[implicits.scala 55:10:@33809.4]
  wire  _T_1977; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:195:@33810.4]
  wire  x855_x524_D5; // @[package.scala 96:25:@33793.4 package.scala 96:25:@33794.4]
  wire  _T_1978; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:283:@33811.4]
  wire  _T_1979; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:291:@33812.4]
  wire  _T_2003; // @[package.scala 96:25:@33851.4 package.scala 96:25:@33852.4]
  wire  _T_2005; // @[implicits.scala 55:10:@33853.4]
  wire  _T_2006; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 834:195:@33854.4]
  wire  x856_x531_D5; // @[package.scala 96:25:@33828.4 package.scala 96:25:@33829.4]
  wire  _T_2007; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 834:283:@33855.4]
  wire  _T_2008; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 834:291:@33856.4]
  wire [7:0] x654_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 734:29:@33479.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:338:@33502.4]
  wire [8:0] _GEN_18; // @[Math.scala 450:32:@33870.4]
  wire [8:0] _T_2016; // @[Math.scala 450:32:@33870.4]
  wire [7:0] x662_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 780:29:@33664.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:338:@33687.4]
  wire [8:0] _GEN_19; // @[Math.scala 450:32:@33875.4]
  wire [8:0] _T_2020; // @[Math.scala 450:32:@33875.4]
  wire [7:0] x656_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 745:29:@33523.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:338:@33546.4]
  wire [8:0] _GEN_20; // @[Math.scala 450:32:@33922.4]
  wire [8:0] _T_2040; // @[Math.scala 450:32:@33922.4]
  wire [7:0] x664_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 797:29:@33708.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:408:@33731.4]
  wire [8:0] _GEN_21; // @[Math.scala 450:32:@33927.4]
  wire [8:0] _T_2044; // @[Math.scala 450:32:@33927.4]
  wire [7:0] x658_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 756:29:@33567.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:338:@33590.4]
  wire [8:0] _GEN_22; // @[Math.scala 450:32:@33974.4]
  wire [8:0] _T_2064; // @[Math.scala 450:32:@33974.4]
  wire [7:0] x666_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 808:29:@33752.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:408:@33775.4]
  wire [8:0] _GEN_23; // @[Math.scala 450:32:@33979.4]
  wire [8:0] _T_2068; // @[Math.scala 450:32:@33979.4]
  wire [7:0] x660_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 767:29:@33611.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:338:@33634.4]
  wire [8:0] _GEN_24; // @[Math.scala 450:32:@34026.4]
  wire [8:0] _T_2088; // @[Math.scala 450:32:@34026.4]
  wire [7:0] x668_rd_0_number; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 819:29:@33796.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:408:@33819.4]
  wire [8:0] _GEN_25; // @[Math.scala 450:32:@34031.4]
  wire [8:0] _T_2092; // @[Math.scala 450:32:@34031.4]
  wire [7:0] x689_div_number; // @[Math.scala 331:22:@34021.4 Math.scala 332:14:@34022.4]
  wire [7:0] x695_div_number; // @[Math.scala 331:22:@34073.4 Math.scala 332:14:@34074.4]
  wire [15:0] _T_2120; // @[Cat.scala 30:58:@34082.4]
  wire [7:0] x677_div_number; // @[Math.scala 331:22:@33917.4 Math.scala 332:14:@33918.4]
  wire [7:0] x683_div_number; // @[Math.scala 331:22:@33969.4 Math.scala 332:14:@33970.4]
  wire [15:0] _T_2121; // @[Cat.scala 30:58:@34083.4]
  wire  _T_2134; // @[package.scala 96:25:@34119.4 package.scala 96:25:@34120.4]
  wire  _T_2136; // @[implicits.scala 55:10:@34121.4]
  wire  x858_b384_D22; // @[package.scala 96:25:@34101.4 package.scala 96:25:@34102.4]
  wire  _T_2137; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 896:116:@34122.4]
  wire  x859_b385_D22; // @[package.scala 96:25:@34110.4 package.scala 96:25:@34111.4]
  wire  _T_2138; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 896:122:@34123.4]
  wire [31:0] x779_x768_D4_number; // @[package.scala 96:25:@31148.4 package.scala 96:25:@31149.4]
  wire [31:0] x780_x401_sum_D3_number; // @[package.scala 96:25:@31157.4 package.scala 96:25:@31158.4]
  wire [31:0] x783_x411_sum_D2_number; // @[package.scala 96:25:@31242.4 package.scala 96:25:@31243.4]
  wire [31:0] x785_x420_sum_D2_number; // @[package.scala 96:25:@31318.4 package.scala 96:25:@31319.4]
  wire [31:0] x786_x429_sum_D2_number; // @[package.scala 96:25:@31385.4 package.scala 96:25:@31386.4]
  wire [31:0] x442_sum_number; // @[Math.scala 154:22:@31527.4 Math.scala 155:14:@31528.4]
  wire [31:0] x795_x770_D2_number; // @[package.scala 96:25:@31554.4 package.scala 96:25:@31555.4]
  wire [31:0] x451_sum_number; // @[Math.scala 154:22:@31630.4 Math.scala 155:14:@31631.4]
  wire [31:0] x459_sum_number; // @[Math.scala 154:22:@31706.4 Math.scala 155:14:@31707.4]
  wire [31:0] x805_x467_sum_D1_number; // @[package.scala 96:25:@31791.4 package.scala 96:25:@31792.4]
  wire [31:0] x478_sum_number; // @[Math.scala 154:22:@31870.4 Math.scala 155:14:@31871.4]
  wire [31:0] x490_sum_number; // @[Math.scala 154:22:@31951.4 Math.scala 155:14:@31952.4]
  wire [31:0] x503_sum_number; // @[Math.scala 154:22:@32052.4 Math.scala 155:14:@32053.4]
  wire [31:0] x810_x772_D1_number; // @[package.scala 96:25:@32070.4 package.scala 96:25:@32071.4]
  wire [31:0] x511_sum_number; // @[Math.scala 154:22:@32112.4 Math.scala 155:14:@32113.4]
  wire [31:0] x518_sum_number; // @[Math.scala 154:22:@32163.4 Math.scala 155:14:@32164.4]
  wire [31:0] x525_sum_number; // @[Math.scala 154:22:@32232.4 Math.scala 155:14:@32233.4]
  wire [31:0] x532_sum_number; // @[Math.scala 154:22:@32283.4 Math.scala 155:14:@32284.4]
  wire [31:0] x539_sum_number; // @[Math.scala 154:22:@32336.4 Math.scala 155:14:@32337.4]
  wire [31:0] x551_sum_number; // @[Math.scala 154:22:@32437.4 Math.scala 155:14:@32438.4]
  wire [31:0] x818_x774_D1_number; // @[package.scala 96:25:@32446.4 package.scala 96:25:@32447.4]
  wire [31:0] x559_sum_number; // @[Math.scala 154:22:@32497.4 Math.scala 155:14:@32498.4]
  wire [31:0] x566_sum_number; // @[Math.scala 154:22:@32548.4 Math.scala 155:14:@32549.4]
  wire [31:0] x573_sum_number; // @[Math.scala 154:22:@32599.4 Math.scala 155:14:@32600.4]
  wire [31:0] x580_sum_number; // @[Math.scala 154:22:@32650.4 Math.scala 155:14:@32651.4]
  wire [31:0] x587_sum_number; // @[Math.scala 154:22:@32701.4 Math.scala 155:14:@32702.4]
  wire [31:0] x831_x768_D12_number; // @[package.scala 96:25:@33269.4 package.scala 96:25:@33270.4]
  wire [31:0] x832_x401_sum_D11_number; // @[package.scala 96:25:@33278.4 package.scala 96:25:@33279.4]
  wire [31:0] x833_x411_sum_D10_number; // @[package.scala 96:25:@33312.4 package.scala 96:25:@33313.4]
  wire [31:0] x834_x420_sum_D10_number; // @[package.scala 96:25:@33346.4 package.scala 96:25:@33347.4]
  wire [31:0] x835_x429_sum_D10_number; // @[package.scala 96:25:@33380.4 package.scala 96:25:@33381.4]
  wire [31:0] x836_x770_D6_number; // @[package.scala 96:25:@33414.4 package.scala 96:25:@33415.4]
  wire [31:0] x838_x442_sum_D4_number; // @[package.scala 96:25:@33432.4 package.scala 96:25:@33433.4]
  wire [31:0] x839_x451_sum_D4_number; // @[package.scala 96:25:@33467.4 package.scala 96:25:@33468.4]
  wire [31:0] x842_x459_sum_D4_number; // @[package.scala 96:25:@33520.4 package.scala 96:25:@33521.4]
  wire [31:0] x843_x467_sum_D5_number; // @[package.scala 96:25:@33555.4 package.scala 96:25:@33556.4]
  wire [31:0] x846_x478_sum_D4_number; // @[package.scala 96:25:@33608.4 package.scala 96:25:@33609.4]
  wire [31:0] x848_x503_sum_D4_number; // @[package.scala 96:25:@33652.4 package.scala 96:25:@33653.4]
  wire [31:0] x849_x772_D5_number; // @[package.scala 96:25:@33661.4 package.scala 96:25:@33662.4]
  wire [31:0] x850_x511_sum_D4_number; // @[package.scala 96:25:@33696.4 package.scala 96:25:@33697.4]
  wire [31:0] x852_x518_sum_D4_number; // @[package.scala 96:25:@33740.4 package.scala 96:25:@33741.4]
  wire [31:0] x854_x525_sum_D4_number; // @[package.scala 96:25:@33784.4 package.scala 96:25:@33785.4]
  wire [31:0] x857_x532_sum_D4_number; // @[package.scala 96:25:@33837.4 package.scala 96:25:@33838.4]
  _ _ ( // @[Math.scala 709:24:@30729.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@30741.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x386_lb_0 x386_lb_0 ( // @[m_x386_lb_0.scala 47:17:@30751.4]
    .clock(x386_lb_0_clock),
    .reset(x386_lb_0_reset),
    .io_rPort_17_banks_0(x386_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x386_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x386_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x386_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x386_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_0(x386_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x386_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x386_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x386_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x386_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_0(x386_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x386_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x386_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x386_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x386_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_0(x386_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x386_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x386_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x386_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x386_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_0(x386_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x386_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x386_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x386_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x386_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_0(x386_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x386_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x386_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x386_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x386_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_0(x386_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x386_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x386_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x386_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x386_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_0(x386_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x386_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x386_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x386_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x386_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_0(x386_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x386_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x386_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x386_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x386_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x386_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x386_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x386_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x386_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x386_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x386_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x386_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x386_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x386_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x386_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x386_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x386_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x386_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x386_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x386_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x386_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x386_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x386_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x386_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x386_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x386_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x386_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x386_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x386_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x386_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x386_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x386_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x386_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x386_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x386_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x386_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x386_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x386_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x386_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x386_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x386_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x386_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x386_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x386_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x386_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x386_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x386_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x386_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x386_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x386_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_0(x386_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x386_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x386_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x386_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x386_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x386_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x386_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x386_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x386_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x386_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x386_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x386_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x386_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x386_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x386_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x386_lb_0_io_wPort_0_en_0)
  );
  x387_lb2_0 x387_lb2_0 ( // @[m_x387_lb2_0.scala 39:17:@30896.4]
    .clock(x387_lb2_0_clock),
    .reset(x387_lb2_0_reset),
    .io_rPort_9_banks_0(x387_lb2_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x387_lb2_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x387_lb2_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x387_lb2_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x387_lb2_0_io_rPort_9_output_0),
    .io_rPort_8_banks_0(x387_lb2_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x387_lb2_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x387_lb2_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x387_lb2_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x387_lb2_0_io_rPort_8_output_0),
    .io_rPort_7_banks_0(x387_lb2_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x387_lb2_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x387_lb2_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x387_lb2_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x387_lb2_0_io_rPort_7_output_0),
    .io_rPort_6_banks_0(x387_lb2_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x387_lb2_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x387_lb2_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x387_lb2_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x387_lb2_0_io_rPort_6_output_0),
    .io_rPort_5_banks_0(x387_lb2_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x387_lb2_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x387_lb2_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x387_lb2_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x387_lb2_0_io_rPort_5_output_0),
    .io_rPort_4_banks_0(x387_lb2_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x387_lb2_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x387_lb2_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x387_lb2_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x387_lb2_0_io_rPort_4_output_0),
    .io_rPort_3_banks_0(x387_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x387_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x387_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x387_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x387_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_0(x387_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x387_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x387_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x387_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x387_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_0(x387_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x387_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x387_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x387_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x387_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_0(x387_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x387_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x387_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x387_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x387_lb2_0_io_rPort_0_output_0),
    .io_wPort_3_banks_0(x387_lb2_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x387_lb2_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x387_lb2_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x387_lb2_0_io_wPort_3_en_0),
    .io_wPort_2_banks_0(x387_lb2_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x387_lb2_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x387_lb2_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x387_lb2_0_io_wPort_2_en_0),
    .io_wPort_1_banks_0(x387_lb2_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x387_lb2_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x387_lb2_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x387_lb2_0_io_wPort_1_en_0),
    .io_wPort_0_banks_0(x387_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x387_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x387_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x387_lb2_0_io_wPort_0_en_0)
  );
  RetimeWrapper_196 RetimeWrapper ( // @[package.scala 93:22:@31006.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x401_sum x401_sum_1 ( // @[Math.scala 150:24:@31106.4]
    .clock(x401_sum_1_clock),
    .reset(x401_sum_1_reset),
    .io_a(x401_sum_1_io_a),
    .io_b(x401_sum_1_io_b),
    .io_flow(x401_sum_1_io_flow),
    .io_result(x401_sum_1_io_result)
  );
  RetimeWrapper_198 RetimeWrapper_1 ( // @[package.scala 93:22:@31116.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_2 ( // @[package.scala 93:22:@31125.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_200 RetimeWrapper_3 ( // @[package.scala 93:22:@31134.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_4 ( // @[package.scala 93:22:@31143.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_202 RetimeWrapper_5 ( // @[package.scala 93:22:@31152.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_6 ( // @[package.scala 93:22:@31165.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x401_sum x407_rdcol_1 ( // @[Math.scala 150:24:@31188.4]
    .clock(x407_rdcol_1_clock),
    .reset(x407_rdcol_1_reset),
    .io_a(x407_rdcol_1_io_a),
    .io_b(x407_rdcol_1_io_b),
    .io_flow(x407_rdcol_1_io_flow),
    .io_result(x407_rdcol_1_io_result)
  );
  RetimeWrapper_196 RetimeWrapper_7 ( // @[package.scala 93:22:@31209.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x401_sum x411_sum_1 ( // @[Math.scala 150:24:@31218.4]
    .clock(x411_sum_1_clock),
    .reset(x411_sum_1_reset),
    .io_a(x411_sum_1_io_a),
    .io_b(x411_sum_1_io_b),
    .io_flow(x411_sum_1_io_flow),
    .io_result(x411_sum_1_io_result)
  );
  RetimeWrapper_200 RetimeWrapper_8 ( // @[package.scala 93:22:@31228.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_208 RetimeWrapper_9 ( // @[package.scala 93:22:@31237.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_10 ( // @[package.scala 93:22:@31250.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x401_sum x416_rdcol_1 ( // @[Math.scala 150:24:@31273.4]
    .clock(x416_rdcol_1_clock),
    .reset(x416_rdcol_1_reset),
    .io_a(x416_rdcol_1_io_a),
    .io_b(x416_rdcol_1_io_b),
    .io_flow(x416_rdcol_1_io_flow),
    .io_result(x416_rdcol_1_io_result)
  );
  x401_sum x420_sum_1 ( // @[Math.scala 150:24:@31294.4]
    .clock(x420_sum_1_clock),
    .reset(x420_sum_1_reset),
    .io_a(x420_sum_1_io_a),
    .io_b(x420_sum_1_io_b),
    .io_flow(x420_sum_1_io_flow),
    .io_result(x420_sum_1_io_result)
  );
  RetimeWrapper_200 RetimeWrapper_11 ( // @[package.scala 93:22:@31304.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_208 RetimeWrapper_12 ( // @[package.scala 93:22:@31313.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_13 ( // @[package.scala 93:22:@31326.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x401_sum x425_rdcol_1 ( // @[Math.scala 150:24:@31349.4]
    .clock(x425_rdcol_1_clock),
    .reset(x425_rdcol_1_reset),
    .io_a(x425_rdcol_1_io_a),
    .io_b(x425_rdcol_1_io_b),
    .io_flow(x425_rdcol_1_io_flow),
    .io_result(x425_rdcol_1_io_result)
  );
  x401_sum x429_sum_1 ( // @[Math.scala 150:24:@31370.4]
    .clock(x429_sum_1_clock),
    .reset(x429_sum_1_reset),
    .io_a(x429_sum_1_io_a),
    .io_b(x429_sum_1_io_b),
    .io_flow(x429_sum_1_io_flow),
    .io_result(x429_sum_1_io_result)
  );
  RetimeWrapper_208 RetimeWrapper_14 ( // @[package.scala 93:22:@31380.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_200 RetimeWrapper_15 ( // @[package.scala 93:22:@31389.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_16 ( // @[package.scala 93:22:@31402.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_17 ( // @[package.scala 93:22:@31423.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_18 ( // @[package.scala 93:22:@31450.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper RetimeWrapper_19 ( // @[package.scala 93:22:@31468.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_196 RetimeWrapper_20 ( // @[package.scala 93:22:@31503.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_21 ( // @[package.scala 93:22:@31512.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  x401_sum x442_sum_1 ( // @[Math.scala 150:24:@31521.4]
    .clock(x442_sum_1_clock),
    .reset(x442_sum_1_reset),
    .io_a(x442_sum_1_io_a),
    .io_b(x442_sum_1_io_b),
    .io_flow(x442_sum_1_io_flow),
    .io_result(x442_sum_1_io_result)
  );
  RetimeWrapper_226 RetimeWrapper_22 ( // @[package.scala 93:22:@31531.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_23 ( // @[package.scala 93:22:@31540.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_208 RetimeWrapper_24 ( // @[package.scala 93:22:@31549.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@31558.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_26 ( // @[package.scala 93:22:@31572.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_27 ( // @[package.scala 93:22:@31593.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_28 ( // @[package.scala 93:22:@31615.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x401_sum x451_sum_1 ( // @[Math.scala 150:24:@31624.4]
    .clock(x451_sum_1_clock),
    .reset(x451_sum_1_reset),
    .io_a(x451_sum_1_io_a),
    .io_b(x451_sum_1_io_b),
    .io_flow(x451_sum_1_io_flow),
    .io_result(x451_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@31634.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_30 ( // @[package.scala 93:22:@31648.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_31 ( // @[package.scala 93:22:@31669.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_32 ( // @[package.scala 93:22:@31691.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x401_sum x459_sum_1 ( // @[Math.scala 150:24:@31700.4]
    .clock(x459_sum_1_clock),
    .reset(x459_sum_1_reset),
    .io_a(x459_sum_1_io_a),
    .io_b(x459_sum_1_io_b),
    .io_flow(x459_sum_1_io_flow),
    .io_result(x459_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_33 ( // @[package.scala 93:22:@31710.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_34 ( // @[package.scala 93:22:@31724.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_35 ( // @[package.scala 93:22:@31745.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_36 ( // @[package.scala 93:22:@31767.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x401_sum x467_sum_1 ( // @[Math.scala 150:24:@31776.4]
    .clock(x467_sum_1_clock),
    .reset(x467_sum_1_reset),
    .io_a(x467_sum_1_io_a),
    .io_b(x467_sum_1_io_b),
    .io_flow(x467_sum_1_io_flow),
    .io_result(x467_sum_1_io_result)
  );
  RetimeWrapper_196 RetimeWrapper_37 ( // @[package.scala 93:22:@31786.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_52 RetimeWrapper_38 ( // @[package.scala 93:22:@31795.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_39 ( // @[package.scala 93:22:@31809.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x401_sum x472_rdcol_1 ( // @[Math.scala 150:24:@31832.4]
    .clock(x472_rdcol_1_clock),
    .reset(x472_rdcol_1_reset),
    .io_a(x472_rdcol_1_io_a),
    .io_b(x472_rdcol_1_io_b),
    .io_flow(x472_rdcol_1_io_flow),
    .io_result(x472_rdcol_1_io_result)
  );
  x401_sum x478_sum_1 ( // @[Math.scala 150:24:@31864.4]
    .clock(x478_sum_1_clock),
    .reset(x478_sum_1_reset),
    .io_a(x478_sum_1_io_a),
    .io_b(x478_sum_1_io_b),
    .io_flow(x478_sum_1_io_flow),
    .io_result(x478_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_40 ( // @[package.scala 93:22:@31874.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_41 ( // @[package.scala 93:22:@31888.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  x401_sum x484_rdcol_1 ( // @[Math.scala 150:24:@31913.4]
    .clock(x484_rdcol_1_clock),
    .reset(x484_rdcol_1_reset),
    .io_a(x484_rdcol_1_io_a),
    .io_b(x484_rdcol_1_io_b),
    .io_flow(x484_rdcol_1_io_flow),
    .io_result(x484_rdcol_1_io_result)
  );
  x401_sum x490_sum_1 ( // @[Math.scala 150:24:@31945.4]
    .clock(x490_sum_1_clock),
    .reset(x490_sum_1_reset),
    .io_a(x490_sum_1_io_a),
    .io_b(x490_sum_1_io_b),
    .io_flow(x490_sum_1_io_flow),
    .io_result(x490_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_42 ( // @[package.scala 93:22:@31955.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_43 ( // @[package.scala 93:22:@31969.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x496_rdrow x496_rdrow_1 ( // @[Math.scala 191:24:@31992.4]
    .clock(x496_rdrow_1_clock),
    .reset(x496_rdrow_1_reset),
    .io_a(x496_rdrow_1_io_a),
    .io_b(x496_rdrow_1_io_b),
    .io_flow(x496_rdrow_1_io_flow),
    .io_result(x496_rdrow_1_io_result)
  );
  x401_sum x503_sum_1 ( // @[Math.scala 150:24:@32046.4]
    .clock(x503_sum_1_clock),
    .reset(x503_sum_1_reset),
    .io_a(x503_sum_1_io_a),
    .io_b(x503_sum_1_io_b),
    .io_flow(x503_sum_1_io_flow),
    .io_result(x503_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@32056.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_196 RetimeWrapper_45 ( // @[package.scala 93:22:@32065.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_46 ( // @[package.scala 93:22:@32079.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  x401_sum x511_sum_1 ( // @[Math.scala 150:24:@32106.4]
    .clock(x511_sum_1_clock),
    .reset(x511_sum_1_reset),
    .io_a(x511_sum_1_io_a),
    .io_b(x511_sum_1_io_b),
    .io_flow(x511_sum_1_io_flow),
    .io_result(x511_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@32116.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_48 ( // @[package.scala 93:22:@32130.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x401_sum x518_sum_1 ( // @[Math.scala 150:24:@32157.4]
    .clock(x518_sum_1_clock),
    .reset(x518_sum_1_reset),
    .io_a(x518_sum_1_io_a),
    .io_b(x518_sum_1_io_b),
    .io_flow(x518_sum_1_io_flow),
    .io_result(x518_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_49 ( // @[package.scala 93:22:@32167.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_50 ( // @[package.scala 93:22:@32181.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper RetimeWrapper_51 ( // @[package.scala 93:22:@32202.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_267 RetimeWrapper_52 ( // @[package.scala 93:22:@32217.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x401_sum x525_sum_1 ( // @[Math.scala 150:24:@32226.4]
    .clock(x525_sum_1_clock),
    .reset(x525_sum_1_reset),
    .io_a(x525_sum_1_io_a),
    .io_b(x525_sum_1_io_b),
    .io_flow(x525_sum_1_io_flow),
    .io_result(x525_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_53 ( // @[package.scala 93:22:@32236.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_54 ( // @[package.scala 93:22:@32250.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x401_sum x532_sum_1 ( // @[Math.scala 150:24:@32277.4]
    .clock(x532_sum_1_clock),
    .reset(x532_sum_1_reset),
    .io_a(x532_sum_1_io_a),
    .io_b(x532_sum_1_io_b),
    .io_flow(x532_sum_1_io_flow),
    .io_result(x532_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_55 ( // @[package.scala 93:22:@32287.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_56 ( // @[package.scala 93:22:@32301.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x401_sum x539_sum_1 ( // @[Math.scala 150:24:@32330.4]
    .clock(x539_sum_1_clock),
    .reset(x539_sum_1_reset),
    .io_a(x539_sum_1_io_a),
    .io_b(x539_sum_1_io_b),
    .io_flow(x539_sum_1_io_flow),
    .io_result(x539_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@32340.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_58 ( // @[package.scala 93:22:@32354.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x496_rdrow x544_rdrow_1 ( // @[Math.scala 191:24:@32377.4]
    .clock(x544_rdrow_1_clock),
    .reset(x544_rdrow_1_reset),
    .io_a(x544_rdrow_1_io_a),
    .io_b(x544_rdrow_1_io_b),
    .io_flow(x544_rdrow_1_io_flow),
    .io_result(x544_rdrow_1_io_result)
  );
  x401_sum x551_sum_1 ( // @[Math.scala 150:24:@32431.4]
    .clock(x551_sum_1_clock),
    .reset(x551_sum_1_reset),
    .io_a(x551_sum_1_io_a),
    .io_b(x551_sum_1_io_b),
    .io_flow(x551_sum_1_io_flow),
    .io_result(x551_sum_1_io_result)
  );
  RetimeWrapper_196 RetimeWrapper_59 ( // @[package.scala 93:22:@32441.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper RetimeWrapper_60 ( // @[package.scala 93:22:@32450.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_61 ( // @[package.scala 93:22:@32464.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x401_sum x559_sum_1 ( // @[Math.scala 150:24:@32491.4]
    .clock(x559_sum_1_clock),
    .reset(x559_sum_1_reset),
    .io_a(x559_sum_1_io_a),
    .io_b(x559_sum_1_io_b),
    .io_flow(x559_sum_1_io_flow),
    .io_result(x559_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@32501.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_63 ( // @[package.scala 93:22:@32515.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x401_sum x566_sum_1 ( // @[Math.scala 150:24:@32542.4]
    .clock(x566_sum_1_clock),
    .reset(x566_sum_1_reset),
    .io_a(x566_sum_1_io_a),
    .io_b(x566_sum_1_io_b),
    .io_flow(x566_sum_1_io_flow),
    .io_result(x566_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_64 ( // @[package.scala 93:22:@32552.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_65 ( // @[package.scala 93:22:@32566.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x401_sum x573_sum_1 ( // @[Math.scala 150:24:@32593.4]
    .clock(x573_sum_1_clock),
    .reset(x573_sum_1_reset),
    .io_a(x573_sum_1_io_a),
    .io_b(x573_sum_1_io_b),
    .io_flow(x573_sum_1_io_flow),
    .io_result(x573_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_66 ( // @[package.scala 93:22:@32603.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_67 ( // @[package.scala 93:22:@32617.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x401_sum x580_sum_1 ( // @[Math.scala 150:24:@32644.4]
    .clock(x580_sum_1_clock),
    .reset(x580_sum_1_reset),
    .io_a(x580_sum_1_io_a),
    .io_b(x580_sum_1_io_b),
    .io_flow(x580_sum_1_io_flow),
    .io_result(x580_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_68 ( // @[package.scala 93:22:@32654.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_69 ( // @[package.scala 93:22:@32668.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x401_sum x587_sum_1 ( // @[Math.scala 150:24:@32695.4]
    .clock(x587_sum_1_clock),
    .reset(x587_sum_1_reset),
    .io_a(x587_sum_1_io_a),
    .io_b(x587_sum_1_io_b),
    .io_flow(x587_sum_1_io_flow),
    .io_result(x587_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_70 ( // @[package.scala 93:22:@32705.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_226 RetimeWrapper_71 ( // @[package.scala 93:22:@32719.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x597_x23 x597_x23_1 ( // @[Math.scala 150:24:@32767.4]
    .clock(x597_x23_1_clock),
    .reset(x597_x23_1_reset),
    .io_a(x597_x23_1_io_a),
    .io_b(x597_x23_1_io_b),
    .io_flow(x597_x23_1_io_flow),
    .io_result(x597_x23_1_io_result)
  );
  x597_x23 x598_x24_1 ( // @[Math.scala 150:24:@32777.4]
    .clock(x598_x24_1_clock),
    .reset(x598_x24_1_reset),
    .io_a(x598_x24_1_io_a),
    .io_b(x598_x24_1_io_b),
    .io_flow(x598_x24_1_io_flow),
    .io_result(x598_x24_1_io_result)
  );
  x597_x23 x599_x23_1 ( // @[Math.scala 150:24:@32787.4]
    .clock(x599_x23_1_clock),
    .reset(x599_x23_1_reset),
    .io_a(x599_x23_1_io_a),
    .io_b(x599_x23_1_io_b),
    .io_flow(x599_x23_1_io_flow),
    .io_result(x599_x23_1_io_result)
  );
  x597_x23 x600_x24_1 ( // @[Math.scala 150:24:@32797.4]
    .clock(x600_x24_1_clock),
    .reset(x600_x24_1_reset),
    .io_a(x600_x24_1_io_a),
    .io_b(x600_x24_1_io_b),
    .io_flow(x600_x24_1_io_flow),
    .io_result(x600_x24_1_io_result)
  );
  x601_x23 x601_x23_1 ( // @[Math.scala 150:24:@32807.4]
    .io_a(x601_x23_1_io_a),
    .io_b(x601_x23_1_io_b),
    .io_result(x601_x23_1_io_result)
  );
  x601_x23 x602_x24_1 ( // @[Math.scala 150:24:@32817.4]
    .io_a(x602_x24_1_io_a),
    .io_b(x602_x24_1_io_b),
    .io_result(x602_x24_1_io_result)
  );
  x601_x23 x603_x23_1 ( // @[Math.scala 150:24:@32827.4]
    .io_a(x603_x23_1_io_a),
    .io_b(x603_x23_1_io_b),
    .io_result(x603_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_72 ( // @[package.scala 93:22:@32837.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x601_x23 x604_sum_1 ( // @[Math.scala 150:24:@32846.4]
    .io_a(x604_sum_1_io_a),
    .io_b(x604_sum_1_io_b),
    .io_result(x604_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_73 ( // @[package.scala 93:22:@32860.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  x597_x23 x611_x23_1 ( // @[Math.scala 150:24:@32895.4]
    .clock(x611_x23_1_clock),
    .reset(x611_x23_1_reset),
    .io_a(x611_x23_1_io_a),
    .io_b(x611_x23_1_io_b),
    .io_flow(x611_x23_1_io_flow),
    .io_result(x611_x23_1_io_result)
  );
  x597_x23 x612_x24_1 ( // @[Math.scala 150:24:@32905.4]
    .clock(x612_x24_1_clock),
    .reset(x612_x24_1_reset),
    .io_a(x612_x24_1_io_a),
    .io_b(x612_x24_1_io_b),
    .io_flow(x612_x24_1_io_flow),
    .io_result(x612_x24_1_io_result)
  );
  x597_x23 x613_x23_1 ( // @[Math.scala 150:24:@32915.4]
    .clock(x613_x23_1_clock),
    .reset(x613_x23_1_reset),
    .io_a(x613_x23_1_io_a),
    .io_b(x613_x23_1_io_b),
    .io_flow(x613_x23_1_io_flow),
    .io_result(x613_x23_1_io_result)
  );
  x597_x23 x614_x24_1 ( // @[Math.scala 150:24:@32925.4]
    .clock(x614_x24_1_clock),
    .reset(x614_x24_1_reset),
    .io_a(x614_x24_1_io_a),
    .io_b(x614_x24_1_io_b),
    .io_flow(x614_x24_1_io_flow),
    .io_result(x614_x24_1_io_result)
  );
  x601_x23 x615_x23_1 ( // @[Math.scala 150:24:@32935.4]
    .io_a(x615_x23_1_io_a),
    .io_b(x615_x23_1_io_b),
    .io_result(x615_x23_1_io_result)
  );
  x601_x23 x616_x24_1 ( // @[Math.scala 150:24:@32945.4]
    .io_a(x616_x24_1_io_a),
    .io_b(x616_x24_1_io_b),
    .io_result(x616_x24_1_io_result)
  );
  x601_x23 x617_x23_1 ( // @[Math.scala 150:24:@32955.4]
    .io_a(x617_x23_1_io_a),
    .io_b(x617_x23_1_io_b),
    .io_result(x617_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_74 ( // @[package.scala 93:22:@32965.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x601_x23 x618_sum_1 ( // @[Math.scala 150:24:@32974.4]
    .io_a(x618_sum_1_io_a),
    .io_b(x618_sum_1_io_b),
    .io_result(x618_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_75 ( // @[package.scala 93:22:@32988.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  x597_x23 x624_x23_1 ( // @[Math.scala 150:24:@33018.4]
    .clock(x624_x23_1_clock),
    .reset(x624_x23_1_reset),
    .io_a(x624_x23_1_io_a),
    .io_b(x624_x23_1_io_b),
    .io_flow(x624_x23_1_io_flow),
    .io_result(x624_x23_1_io_result)
  );
  x597_x23 x625_x24_1 ( // @[Math.scala 150:24:@33028.4]
    .clock(x625_x24_1_clock),
    .reset(x625_x24_1_reset),
    .io_a(x625_x24_1_io_a),
    .io_b(x625_x24_1_io_b),
    .io_flow(x625_x24_1_io_flow),
    .io_result(x625_x24_1_io_result)
  );
  x597_x23 x626_x23_1 ( // @[Math.scala 150:24:@33038.4]
    .clock(x626_x23_1_clock),
    .reset(x626_x23_1_reset),
    .io_a(x626_x23_1_io_a),
    .io_b(x626_x23_1_io_b),
    .io_flow(x626_x23_1_io_flow),
    .io_result(x626_x23_1_io_result)
  );
  x597_x23 x627_x24_1 ( // @[Math.scala 150:24:@33048.4]
    .clock(x627_x24_1_clock),
    .reset(x627_x24_1_reset),
    .io_a(x627_x24_1_io_a),
    .io_b(x627_x24_1_io_b),
    .io_flow(x627_x24_1_io_flow),
    .io_result(x627_x24_1_io_result)
  );
  x601_x23 x628_x23_1 ( // @[Math.scala 150:24:@33058.4]
    .io_a(x628_x23_1_io_a),
    .io_b(x628_x23_1_io_b),
    .io_result(x628_x23_1_io_result)
  );
  x601_x23 x629_x24_1 ( // @[Math.scala 150:24:@33068.4]
    .io_a(x629_x24_1_io_a),
    .io_b(x629_x24_1_io_b),
    .io_result(x629_x24_1_io_result)
  );
  x601_x23 x630_x23_1 ( // @[Math.scala 150:24:@33078.4]
    .io_a(x630_x23_1_io_a),
    .io_b(x630_x23_1_io_b),
    .io_result(x630_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_76 ( // @[package.scala 93:22:@33088.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  x601_x23 x631_sum_1 ( // @[Math.scala 150:24:@33097.4]
    .io_a(x631_sum_1_io_a),
    .io_b(x631_sum_1_io_b),
    .io_result(x631_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_77 ( // @[package.scala 93:22:@33111.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x597_x23 x637_x23_1 ( // @[Math.scala 150:24:@33141.4]
    .clock(x637_x23_1_clock),
    .reset(x637_x23_1_reset),
    .io_a(x637_x23_1_io_a),
    .io_b(x637_x23_1_io_b),
    .io_flow(x637_x23_1_io_flow),
    .io_result(x637_x23_1_io_result)
  );
  x597_x23 x638_x24_1 ( // @[Math.scala 150:24:@33153.4]
    .clock(x638_x24_1_clock),
    .reset(x638_x24_1_reset),
    .io_a(x638_x24_1_io_a),
    .io_b(x638_x24_1_io_b),
    .io_flow(x638_x24_1_io_flow),
    .io_result(x638_x24_1_io_result)
  );
  x597_x23 x639_x23_1 ( // @[Math.scala 150:24:@33163.4]
    .clock(x639_x23_1_clock),
    .reset(x639_x23_1_reset),
    .io_a(x639_x23_1_io_a),
    .io_b(x639_x23_1_io_b),
    .io_flow(x639_x23_1_io_flow),
    .io_result(x639_x23_1_io_result)
  );
  x597_x23 x640_x24_1 ( // @[Math.scala 150:24:@33173.4]
    .clock(x640_x24_1_clock),
    .reset(x640_x24_1_reset),
    .io_a(x640_x24_1_io_a),
    .io_b(x640_x24_1_io_b),
    .io_flow(x640_x24_1_io_flow),
    .io_result(x640_x24_1_io_result)
  );
  x601_x23 x641_x23_1 ( // @[Math.scala 150:24:@33183.4]
    .io_a(x641_x23_1_io_a),
    .io_b(x641_x23_1_io_b),
    .io_result(x641_x23_1_io_result)
  );
  x601_x23 x642_x24_1 ( // @[Math.scala 150:24:@33193.4]
    .io_a(x642_x24_1_io_a),
    .io_b(x642_x24_1_io_b),
    .io_result(x642_x24_1_io_result)
  );
  x601_x23 x643_x23_1 ( // @[Math.scala 150:24:@33203.4]
    .io_a(x643_x23_1_io_a),
    .io_b(x643_x23_1_io_b),
    .io_result(x643_x23_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_78 ( // @[package.scala 93:22:@33213.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  x601_x23 x644_sum_1 ( // @[Math.scala 150:24:@33222.4]
    .io_a(x644_sum_1_io_a),
    .io_b(x644_sum_1_io_b),
    .io_result(x644_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_79 ( // @[package.scala 93:22:@33236.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_80 ( // @[package.scala 93:22:@33246.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_81 ( // @[package.scala 93:22:@33255.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_323 RetimeWrapper_82 ( // @[package.scala 93:22:@33264.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_324 RetimeWrapper_83 ( // @[package.scala 93:22:@33273.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_84 ( // @[package.scala 93:22:@33286.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_85 ( // @[package.scala 93:22:@33307.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_86 ( // @[package.scala 93:22:@33320.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_87 ( // @[package.scala 93:22:@33341.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_88 ( // @[package.scala 93:22:@33354.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_89 ( // @[package.scala 93:22:@33375.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_90 ( // @[package.scala 93:22:@33388.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_91 ( // @[package.scala 93:22:@33409.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_92 ( // @[package.scala 93:22:@33418.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_93 ( // @[package.scala 93:22:@33427.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_94 ( // @[package.scala 93:22:@33441.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_95 ( // @[package.scala 93:22:@33462.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_96 ( // @[package.scala 93:22:@33471.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_97 ( // @[package.scala 93:22:@33485.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_98 ( // @[package.scala 93:22:@33506.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_99 ( // @[package.scala 93:22:@33515.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_100 ( // @[package.scala 93:22:@33529.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_342 RetimeWrapper_101 ( // @[package.scala 93:22:@33550.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_343 RetimeWrapper_102 ( // @[package.scala 93:22:@33559.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_103 ( // @[package.scala 93:22:@33573.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_104 ( // @[package.scala 93:22:@33594.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_105 ( // @[package.scala 93:22:@33603.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_106 ( // @[package.scala 93:22:@33617.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_107 ( // @[package.scala 93:22:@33638.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_108 ( // @[package.scala 93:22:@33647.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_342 RetimeWrapper_109 ( // @[package.scala 93:22:@33656.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_110 ( // @[package.scala 93:22:@33670.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_111 ( // @[package.scala 93:22:@33691.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_112 ( // @[package.scala 93:22:@33700.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_113 ( // @[package.scala 93:22:@33714.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_114 ( // @[package.scala 93:22:@33735.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_115 ( // @[package.scala 93:22:@33744.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_116 ( // @[package.scala 93:22:@33758.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_117 ( // @[package.scala 93:22:@33779.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_118 ( // @[package.scala 93:22:@33788.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_119 ( // @[package.scala 93:22:@33802.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_120 ( // @[package.scala 93:22:@33823.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_121 ( // @[package.scala 93:22:@33832.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_321 RetimeWrapper_122 ( // @[package.scala 93:22:@33846.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  x601_x23 x674_x25_1 ( // @[Math.scala 150:24:@33879.4]
    .io_a(x674_x25_1_io_a),
    .io_b(x674_x25_1_io_b),
    .io_result(x674_x25_1_io_result)
  );
  x601_x23 x675_x26_1 ( // @[Math.scala 150:24:@33889.4]
    .io_a(x675_x26_1_io_a),
    .io_b(x675_x26_1_io_b),
    .io_result(x675_x26_1_io_result)
  );
  x601_x23 x676_sum_1 ( // @[Math.scala 150:24:@33899.4]
    .io_a(x676_sum_1_io_a),
    .io_b(x676_sum_1_io_b),
    .io_result(x676_sum_1_io_result)
  );
  x677_div x677_div_1 ( // @[Math.scala 327:24:@33911.4]
    .clock(x677_div_1_clock),
    .reset(x677_div_1_reset),
    .io_a(x677_div_1_io_a),
    .io_flow(x677_div_1_io_flow),
    .io_result(x677_div_1_io_result)
  );
  x601_x23 x680_x25_1 ( // @[Math.scala 150:24:@33931.4]
    .io_a(x680_x25_1_io_a),
    .io_b(x680_x25_1_io_b),
    .io_result(x680_x25_1_io_result)
  );
  x601_x23 x681_x26_1 ( // @[Math.scala 150:24:@33941.4]
    .io_a(x681_x26_1_io_a),
    .io_b(x681_x26_1_io_b),
    .io_result(x681_x26_1_io_result)
  );
  x601_x23 x682_sum_1 ( // @[Math.scala 150:24:@33951.4]
    .io_a(x682_sum_1_io_a),
    .io_b(x682_sum_1_io_b),
    .io_result(x682_sum_1_io_result)
  );
  x677_div x683_div_1 ( // @[Math.scala 327:24:@33963.4]
    .clock(x683_div_1_clock),
    .reset(x683_div_1_reset),
    .io_a(x683_div_1_io_a),
    .io_flow(x683_div_1_io_flow),
    .io_result(x683_div_1_io_result)
  );
  x601_x23 x686_x25_1 ( // @[Math.scala 150:24:@33983.4]
    .io_a(x686_x25_1_io_a),
    .io_b(x686_x25_1_io_b),
    .io_result(x686_x25_1_io_result)
  );
  x601_x23 x687_x26_1 ( // @[Math.scala 150:24:@33993.4]
    .io_a(x687_x26_1_io_a),
    .io_b(x687_x26_1_io_b),
    .io_result(x687_x26_1_io_result)
  );
  x601_x23 x688_sum_1 ( // @[Math.scala 150:24:@34003.4]
    .io_a(x688_sum_1_io_a),
    .io_b(x688_sum_1_io_b),
    .io_result(x688_sum_1_io_result)
  );
  x677_div x689_div_1 ( // @[Math.scala 327:24:@34015.4]
    .clock(x689_div_1_clock),
    .reset(x689_div_1_reset),
    .io_a(x689_div_1_io_a),
    .io_flow(x689_div_1_io_flow),
    .io_result(x689_div_1_io_result)
  );
  x601_x23 x692_x25_1 ( // @[Math.scala 150:24:@34035.4]
    .io_a(x692_x25_1_io_a),
    .io_b(x692_x25_1_io_b),
    .io_result(x692_x25_1_io_result)
  );
  x601_x23 x693_x26_1 ( // @[Math.scala 150:24:@34045.4]
    .io_a(x693_x26_1_io_a),
    .io_b(x693_x26_1_io_b),
    .io_result(x693_x26_1_io_result)
  );
  x601_x23 x694_sum_1 ( // @[Math.scala 150:24:@34055.4]
    .io_a(x694_sum_1_io_a),
    .io_b(x694_sum_1_io_b),
    .io_result(x694_sum_1_io_result)
  );
  x677_div x695_div_1 ( // @[Math.scala 327:24:@34067.4]
    .clock(x695_div_1_clock),
    .reset(x695_div_1_reset),
    .io_a(x695_div_1_io_a),
    .io_flow(x695_div_1_io_flow),
    .io_result(x695_div_1_io_result)
  );
  RetimeWrapper_202 RetimeWrapper_123 ( // @[package.scala 93:22:@34087.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_369 RetimeWrapper_124 ( // @[package.scala 93:22:@34096.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_369 RetimeWrapper_125 ( // @[package.scala 93:22:@34105.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_369 RetimeWrapper_126 ( // @[package.scala 93:22:@34114.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  assign b384 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 62:18:@30749.4]
  assign b385 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 63:18:@30750.4]
  assign _T_207 = b384 & b385; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 69:30:@30994.4]
  assign _T_208 = _T_207 & io_sigsIn_datapathEn; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 69:37:@30995.4]
  assign _T_212 = io_in_x373_TID == 8'h0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:76:@31000.4]
  assign _T_213 = _T_208 & _T_212; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:62:@31001.4]
  assign _T_215 = io_in_x373_TDEST == 8'h0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:101:@31002.4]
  assign x775_x388_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@31011.4 package.scala 96:25:@31012.4]
  assign b382_number = __io_result; // @[Math.scala 712:22:@30734.4 Math.scala 713:14:@30735.4]
  assign _T_247 = $signed(b382_number); // @[Math.scala 499:52:@31031.4]
  assign x392 = $signed(32'sh1) == $signed(_T_247); // @[Math.scala 499:44:@31039.4]
  assign x393 = $signed(32'sh2) == $signed(_T_247); // @[Math.scala 499:44:@31046.4]
  assign x394 = $signed(32'sh3) == $signed(_T_247); // @[Math.scala 499:44:@31053.4]
  assign _T_294 = x392 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@31065.4]
  assign _T_296 = x393 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@31066.4]
  assign _T_298 = x394 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@31067.4]
  assign _T_300 = _T_294 | _T_296; // @[Mux.scala 19:72:@31069.4]
  assign x395_number = _T_300 | _T_298; // @[Mux.scala 19:72:@31070.4]
  assign _T_312 = $signed(x395_number); // @[Math.scala 406:49:@31080.4]
  assign _T_314 = $signed(_T_312) & $signed(32'sh3); // @[Math.scala 406:56:@31082.4]
  assign _T_315 = $signed(_T_314); // @[Math.scala 406:56:@31083.4]
  assign _T_320 = x395_number[31]; // @[FixedPoint.scala 50:25:@31089.4]
  assign _T_324 = _T_320 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31091.4]
  assign _T_325 = x395_number[31:2]; // @[FixedPoint.scala 18:52:@31092.4]
  assign b383_number = __1_io_result; // @[Math.scala 712:22:@30746.4 Math.scala 713:14:@30747.4]
  assign _T_330 = b383_number[31]; // @[FixedPoint.scala 50:25:@31098.4]
  assign _T_334 = _T_330 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31100.4]
  assign _T_335 = b383_number[31:2]; // @[FixedPoint.scala 18:52:@31101.4]
  assign _T_360 = ~ io_sigsIn_break; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:101:@31162.4]
  assign _T_364 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@31170.4 package.scala 96:25:@31171.4]
  assign _T_366 = io_rr ? _T_364 : 1'h0; // @[implicits.scala 55:10:@31172.4]
  assign _T_367 = _T_360 & _T_366; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:118:@31173.4]
  assign _T_369 = _T_367 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:205:@31175.4]
  assign _T_370 = _T_369 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:224:@31176.4]
  assign x777_b384_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@31130.4 package.scala 96:25:@31131.4]
  assign _T_371 = _T_370 & x777_b384_D4; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 114:250:@31177.4]
  assign x776_b385_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31121.4 package.scala 96:25:@31122.4]
  assign x407_rdcol_number = x407_rdcol_1_io_result; // @[Math.scala 154:22:@31194.4 Math.scala 155:14:@31195.4]
  assign _T_384 = x407_rdcol_number[31]; // @[FixedPoint.scala 50:25:@31201.4]
  assign _T_388 = _T_384 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31203.4]
  assign _T_389 = x407_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@31204.4]
  assign _T_412 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@31255.4 package.scala 96:25:@31256.4]
  assign _T_414 = io_rr ? _T_412 : 1'h0; // @[implicits.scala 55:10:@31257.4]
  assign _T_415 = _T_360 & _T_414; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:118:@31258.4]
  assign _T_417 = _T_415 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:205:@31260.4]
  assign _T_418 = _T_417 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:224:@31261.4]
  assign _T_419 = _T_418 & x777_b384_D4; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 133:250:@31262.4]
  assign x416_rdcol_number = x416_rdcol_1_io_result; // @[Math.scala 154:22:@31279.4 Math.scala 155:14:@31280.4]
  assign _T_432 = x416_rdcol_number[31]; // @[FixedPoint.scala 50:25:@31286.4]
  assign _T_436 = _T_432 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31288.4]
  assign _T_437 = x416_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@31289.4]
  assign _T_457 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@31331.4 package.scala 96:25:@31332.4]
  assign _T_459 = io_rr ? _T_457 : 1'h0; // @[implicits.scala 55:10:@31333.4]
  assign _T_460 = _T_360 & _T_459; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:118:@31334.4]
  assign _T_462 = _T_460 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:205:@31336.4]
  assign _T_463 = _T_462 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:224:@31337.4]
  assign _T_464 = _T_463 & x777_b384_D4; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 150:250:@31338.4]
  assign x425_rdcol_number = x425_rdcol_1_io_result; // @[Math.scala 154:22:@31355.4 Math.scala 155:14:@31356.4]
  assign _T_477 = x425_rdcol_number[31]; // @[FixedPoint.scala 50:25:@31362.4]
  assign _T_481 = _T_477 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31364.4]
  assign _T_482 = x425_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@31365.4]
  assign _T_502 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@31407.4 package.scala 96:25:@31408.4]
  assign _T_504 = io_rr ? _T_502 : 1'h0; // @[implicits.scala 55:10:@31409.4]
  assign _T_505 = _T_360 & _T_504; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:118:@31410.4]
  assign _T_507 = _T_505 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:205:@31412.4]
  assign _T_508 = _T_507 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:224:@31413.4]
  assign _T_509 = _T_508 & x777_b384_D4; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 167:250:@31414.4]
  assign x788_b382_D6_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@31428.4 package.scala 96:25:@31429.4]
  assign _T_521 = $signed(x788_b382_D6_number); // @[Math.scala 406:49:@31435.4]
  assign _T_523 = $signed(_T_521) & $signed(32'sh3); // @[Math.scala 406:56:@31437.4]
  assign _T_524 = $signed(_T_523); // @[Math.scala 406:56:@31438.4]
  assign x769_number = $unsigned(_T_524); // @[implicits.scala 133:21:@31439.4]
  assign x436 = $signed(_T_521) < $signed(32'sh0); // @[Math.scala 465:44:@31447.4]
  assign x789_x425_rdcol_D6_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@31455.4 package.scala 96:25:@31456.4]
  assign _T_544 = $signed(x789_x425_rdcol_D6_number); // @[Math.scala 465:37:@31463.4]
  assign x437 = $signed(_T_544) < $signed(32'sh0); // @[Math.scala 465:44:@31465.4]
  assign x790_x436_D1 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@31473.4 package.scala 96:25:@31474.4]
  assign x438 = x790_x436_D1 | x437; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 190:24:@31477.4]
  assign _T_561 = $signed(x769_number); // @[Math.scala 406:49:@31486.4]
  assign _T_563 = $signed(_T_561) & $signed(32'sh3); // @[Math.scala 406:56:@31488.4]
  assign _T_564 = $signed(_T_563); // @[Math.scala 406:56:@31489.4]
  assign _T_569 = x769_number[31]; // @[FixedPoint.scala 50:25:@31495.4]
  assign _T_573 = _T_569 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31497.4]
  assign _T_574 = x769_number[31:2]; // @[FixedPoint.scala 18:52:@31498.4]
  assign _T_612 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@31577.4 package.scala 96:25:@31578.4]
  assign _T_614 = io_rr ? _T_612 : 1'h0; // @[implicits.scala 55:10:@31579.4]
  assign _T_615 = _T_360 & _T_614; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 215:194:@31580.4]
  assign x796_x439_D1 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@31563.4 package.scala 96:25:@31564.4]
  assign _T_616 = _T_615 & x796_x439_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 215:281:@31581.4]
  assign x794_b384_D8 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@31545.4 package.scala 96:25:@31546.4]
  assign _T_617 = _T_616 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 215:289:@31582.4]
  assign x793_b385_D8 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@31536.4 package.scala 96:25:@31537.4]
  assign x797_x416_rdcol_D6_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@31598.4 package.scala 96:25:@31599.4]
  assign _T_628 = $signed(x797_x416_rdcol_D6_number); // @[Math.scala 465:37:@31604.4]
  assign x448 = $signed(_T_628) < $signed(32'sh0); // @[Math.scala 465:44:@31606.4]
  assign x449 = x790_x436_D1 | x448; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 223:24:@31609.4]
  assign _T_659 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@31653.4 package.scala 96:25:@31654.4]
  assign _T_661 = io_rr ? _T_659 : 1'h0; // @[implicits.scala 55:10:@31655.4]
  assign _T_662 = _T_360 & _T_661; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:194:@31656.4]
  assign x799_x450_D1 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@31639.4 package.scala 96:25:@31640.4]
  assign _T_663 = _T_662 & x799_x450_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:281:@31657.4]
  assign _T_664 = _T_663 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:289:@31658.4]
  assign x800_x407_rdcol_D6_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@31674.4 package.scala 96:25:@31675.4]
  assign _T_675 = $signed(x800_x407_rdcol_D6_number); // @[Math.scala 465:37:@31680.4]
  assign x456 = $signed(_T_675) < $signed(32'sh0); // @[Math.scala 465:44:@31682.4]
  assign x457 = x790_x436_D1 | x456; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 244:24:@31685.4]
  assign _T_706 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@31729.4 package.scala 96:25:@31730.4]
  assign _T_708 = io_rr ? _T_706 : 1'h0; // @[implicits.scala 55:10:@31731.4]
  assign _T_709 = _T_360 & _T_708; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:194:@31732.4]
  assign x802_x458_D1 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@31715.4 package.scala 96:25:@31716.4]
  assign _T_710 = _T_709 & x802_x458_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:281:@31733.4]
  assign _T_711 = _T_710 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:289:@31734.4]
  assign x803_b383_D6_number = RetimeWrapper_35_io_out; // @[package.scala 96:25:@31750.4 package.scala 96:25:@31751.4]
  assign _T_722 = $signed(x803_b383_D6_number); // @[Math.scala 465:37:@31756.4]
  assign x464 = $signed(_T_722) < $signed(32'sh0); // @[Math.scala 465:44:@31758.4]
  assign x465 = x436 | x464; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 265:59:@31761.4]
  assign _T_756 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@31814.4 package.scala 96:25:@31815.4]
  assign _T_758 = io_rr ? _T_756 : 1'h0; // @[implicits.scala 55:10:@31816.4]
  assign _T_759 = _T_360 & _T_758; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:194:@31817.4]
  assign x806_x466_D2 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@31800.4 package.scala 96:25:@31801.4]
  assign _T_760 = _T_759 & x806_x466_D2; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:281:@31818.4]
  assign _T_761 = _T_760 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:289:@31819.4]
  assign x472_rdcol_number = x472_rdcol_1_io_result; // @[Math.scala 154:22:@31838.4 Math.scala 155:14:@31839.4]
  assign _T_776 = $signed(x472_rdcol_number); // @[Math.scala 465:37:@31844.4]
  assign x473 = $signed(_T_776) < $signed(32'sh0); // @[Math.scala 465:44:@31846.4]
  assign x474 = x790_x436_D1 | x473; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 288:24:@31849.4]
  assign _T_786 = x472_rdcol_number[31]; // @[FixedPoint.scala 50:25:@31856.4]
  assign _T_790 = _T_786 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31858.4]
  assign _T_791 = x472_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@31859.4]
  assign _T_814 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@31893.4 package.scala 96:25:@31894.4]
  assign _T_816 = io_rr ? _T_814 : 1'h0; // @[implicits.scala 55:10:@31895.4]
  assign _T_817 = _T_360 & _T_816; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:194:@31896.4]
  assign x807_x475_D1 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@31879.4 package.scala 96:25:@31880.4]
  assign _T_818 = _T_817 & x807_x475_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:281:@31897.4]
  assign _T_819 = _T_818 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:289:@31898.4]
  assign x484_rdcol_number = x484_rdcol_1_io_result; // @[Math.scala 154:22:@31919.4 Math.scala 155:14:@31920.4]
  assign _T_836 = $signed(x484_rdcol_number); // @[Math.scala 465:37:@31925.4]
  assign x485 = $signed(_T_836) < $signed(32'sh0); // @[Math.scala 465:44:@31927.4]
  assign x486 = x790_x436_D1 | x485; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 317:59:@31930.4]
  assign _T_846 = x484_rdcol_number[31]; // @[FixedPoint.scala 50:25:@31937.4]
  assign _T_850 = _T_846 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@31939.4]
  assign _T_851 = x484_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@31940.4]
  assign _T_874 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@31974.4 package.scala 96:25:@31975.4]
  assign _T_876 = io_rr ? _T_874 : 1'h0; // @[implicits.scala 55:10:@31976.4]
  assign _T_877 = _T_360 & _T_876; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 330:194:@31977.4]
  assign x808_x487_D1 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@31960.4 package.scala 96:25:@31961.4]
  assign _T_878 = _T_877 & x808_x487_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 330:281:@31978.4]
  assign _T_879 = _T_878 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 330:289:@31979.4]
  assign x496_rdrow_number = x496_rdrow_1_io_result; // @[Math.scala 195:22:@31998.4 Math.scala 196:14:@31999.4]
  assign _T_896 = $signed(x496_rdrow_number); // @[Math.scala 406:49:@32005.4]
  assign _T_898 = $signed(_T_896) & $signed(32'sh3); // @[Math.scala 406:56:@32007.4]
  assign _T_899 = $signed(_T_898); // @[Math.scala 406:56:@32008.4]
  assign x771_number = $unsigned(_T_899); // @[implicits.scala 133:21:@32009.4]
  assign x498 = $signed(_T_896) < $signed(32'sh0); // @[Math.scala 465:44:@32017.4]
  assign x499 = x498 | x437; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 340:24:@32020.4]
  assign _T_920 = $signed(x771_number); // @[Math.scala 406:49:@32029.4]
  assign _T_922 = $signed(_T_920) & $signed(32'sh3); // @[Math.scala 406:56:@32031.4]
  assign _T_923 = $signed(_T_922); // @[Math.scala 406:56:@32032.4]
  assign _T_928 = x771_number[31]; // @[FixedPoint.scala 50:25:@32038.4]
  assign _T_932 = _T_928 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32040.4]
  assign _T_933 = x771_number[31:2]; // @[FixedPoint.scala 18:52:@32041.4]
  assign _T_959 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@32084.4 package.scala 96:25:@32085.4]
  assign _T_961 = io_rr ? _T_959 : 1'h0; // @[implicits.scala 55:10:@32086.4]
  assign _T_962 = _T_360 & _T_961; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:194:@32087.4]
  assign x809_x500_D1 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@32061.4 package.scala 96:25:@32062.4]
  assign _T_963 = _T_962 & x809_x500_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:281:@32088.4]
  assign _T_964 = _T_963 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:289:@32089.4]
  assign x509 = x498 | x448; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 361:24:@32100.4]
  assign _T_992 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@32135.4 package.scala 96:25:@32136.4]
  assign _T_994 = io_rr ? _T_992 : 1'h0; // @[implicits.scala 55:10:@32137.4]
  assign _T_995 = _T_360 & _T_994; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:194:@32138.4]
  assign x811_x510_D1 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@32121.4 package.scala 96:25:@32122.4]
  assign _T_996 = _T_995 & x811_x510_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:281:@32139.4]
  assign _T_997 = _T_996 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:289:@32140.4]
  assign x516 = x498 | x456; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 376:24:@32151.4]
  assign _T_1025 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@32186.4 package.scala 96:25:@32187.4]
  assign _T_1027 = io_rr ? _T_1025 : 1'h0; // @[implicits.scala 55:10:@32188.4]
  assign _T_1028 = _T_360 & _T_1027; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:194:@32189.4]
  assign x812_x517_D1 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@32172.4 package.scala 96:25:@32173.4]
  assign _T_1029 = _T_1028 & x812_x517_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:281:@32190.4]
  assign _T_1030 = _T_1029 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:289:@32191.4]
  assign x813_x464_D1 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@32207.4 package.scala 96:25:@32208.4]
  assign x523 = x498 | x813_x464_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 393:24:@32211.4]
  assign _T_1064 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@32255.4 package.scala 96:25:@32256.4]
  assign _T_1066 = io_rr ? _T_1064 : 1'h0; // @[implicits.scala 55:10:@32257.4]
  assign _T_1067 = _T_360 & _T_1066; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:194:@32258.4]
  assign x815_x524_D1 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@32241.4 package.scala 96:25:@32242.4]
  assign _T_1068 = _T_1067 & x815_x524_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:281:@32259.4]
  assign _T_1069 = _T_1068 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:289:@32260.4]
  assign x530 = x498 | x473; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 410:24:@32271.4]
  assign _T_1097 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@32306.4 package.scala 96:25:@32307.4]
  assign _T_1099 = io_rr ? _T_1097 : 1'h0; // @[implicits.scala 55:10:@32308.4]
  assign _T_1100 = _T_360 & _T_1099; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:194:@32309.4]
  assign x816_x531_D1 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@32292.4 package.scala 96:25:@32293.4]
  assign _T_1101 = _T_1100 & x816_x531_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:281:@32310.4]
  assign _T_1102 = _T_1101 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:289:@32311.4]
  assign x537 = x498 | x485; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 431:59:@32322.4]
  assign _T_1132 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@32359.4 package.scala 96:25:@32360.4]
  assign _T_1134 = io_rr ? _T_1132 : 1'h0; // @[implicits.scala 55:10:@32361.4]
  assign _T_1135 = _T_360 & _T_1134; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:194:@32362.4]
  assign x817_x538_D1 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@32345.4 package.scala 96:25:@32346.4]
  assign _T_1136 = _T_1135 & x817_x538_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:281:@32363.4]
  assign _T_1137 = _T_1136 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:289:@32364.4]
  assign x544_rdrow_number = x544_rdrow_1_io_result; // @[Math.scala 195:22:@32383.4 Math.scala 196:14:@32384.4]
  assign _T_1154 = $signed(x544_rdrow_number); // @[Math.scala 406:49:@32390.4]
  assign _T_1156 = $signed(_T_1154) & $signed(32'sh3); // @[Math.scala 406:56:@32392.4]
  assign _T_1157 = $signed(_T_1156); // @[Math.scala 406:56:@32393.4]
  assign x773_number = $unsigned(_T_1157); // @[implicits.scala 133:21:@32394.4]
  assign x546 = $signed(_T_1154) < $signed(32'sh0); // @[Math.scala 465:44:@32402.4]
  assign x547 = x546 | x437; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 454:24:@32405.4]
  assign _T_1178 = $signed(x773_number); // @[Math.scala 406:49:@32414.4]
  assign _T_1180 = $signed(_T_1178) & $signed(32'sh3); // @[Math.scala 406:56:@32416.4]
  assign _T_1181 = $signed(_T_1180); // @[Math.scala 406:56:@32417.4]
  assign _T_1186 = x773_number[31]; // @[FixedPoint.scala 50:25:@32423.4]
  assign _T_1190 = _T_1186 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@32425.4]
  assign _T_1191 = x773_number[31:2]; // @[FixedPoint.scala 18:52:@32426.4]
  assign _T_1217 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@32469.4 package.scala 96:25:@32470.4]
  assign _T_1219 = io_rr ? _T_1217 : 1'h0; // @[implicits.scala 55:10:@32471.4]
  assign _T_1220 = _T_360 & _T_1219; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 471:194:@32472.4]
  assign x819_x548_D1 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@32455.4 package.scala 96:25:@32456.4]
  assign _T_1221 = _T_1220 & x819_x548_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 471:281:@32473.4]
  assign _T_1222 = _T_1221 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 471:289:@32474.4]
  assign x557 = x546 | x448; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 475:24:@32485.4]
  assign _T_1250 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@32520.4 package.scala 96:25:@32521.4]
  assign _T_1252 = io_rr ? _T_1250 : 1'h0; // @[implicits.scala 55:10:@32522.4]
  assign _T_1253 = _T_360 & _T_1252; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:194:@32523.4]
  assign x820_x558_D1 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@32506.4 package.scala 96:25:@32507.4]
  assign _T_1254 = _T_1253 & x820_x558_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:281:@32524.4]
  assign _T_1255 = _T_1254 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:289:@32525.4]
  assign x564 = x546 | x456; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 490:24:@32536.4]
  assign _T_1283 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@32571.4 package.scala 96:25:@32572.4]
  assign _T_1285 = io_rr ? _T_1283 : 1'h0; // @[implicits.scala 55:10:@32573.4]
  assign _T_1286 = _T_360 & _T_1285; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:194:@32574.4]
  assign x821_x565_D1 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@32557.4 package.scala 96:25:@32558.4]
  assign _T_1287 = _T_1286 & x821_x565_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:281:@32575.4]
  assign _T_1288 = _T_1287 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:289:@32576.4]
  assign x571 = x546 | x813_x464_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 505:24:@32587.4]
  assign _T_1316 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@32622.4 package.scala 96:25:@32623.4]
  assign _T_1318 = io_rr ? _T_1316 : 1'h0; // @[implicits.scala 55:10:@32624.4]
  assign _T_1319 = _T_360 & _T_1318; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:194:@32625.4]
  assign x822_x572_D1 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@32608.4 package.scala 96:25:@32609.4]
  assign _T_1320 = _T_1319 & x822_x572_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:281:@32626.4]
  assign _T_1321 = _T_1320 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:289:@32627.4]
  assign x578 = x546 | x473; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 520:24:@32638.4]
  assign _T_1349 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@32673.4 package.scala 96:25:@32674.4]
  assign _T_1351 = io_rr ? _T_1349 : 1'h0; // @[implicits.scala 55:10:@32675.4]
  assign _T_1352 = _T_360 & _T_1351; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:194:@32676.4]
  assign x823_x579_D1 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@32659.4 package.scala 96:25:@32660.4]
  assign _T_1353 = _T_1352 & x823_x579_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:281:@32677.4]
  assign _T_1354 = _T_1353 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:289:@32678.4]
  assign x585 = x546 | x485; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 535:24:@32689.4]
  assign _T_1382 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@32724.4 package.scala 96:25:@32725.4]
  assign _T_1384 = io_rr ? _T_1382 : 1'h0; // @[implicits.scala 55:10:@32726.4]
  assign _T_1385 = _T_360 & _T_1384; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 546:194:@32727.4]
  assign x824_x586_D1 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@32710.4 package.scala 96:25:@32711.4]
  assign _T_1386 = _T_1385 & x824_x586_D1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 546:281:@32728.4]
  assign _T_1387 = _T_1386 & x794_b384_D8; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 546:289:@32729.4]
  assign x454_rd_0_number = x386_lb_0_io_rPort_17_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 232:29:@31642.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 236:336:@31665.4]
  assign _GEN_0 = {{1'd0}, x454_rd_0_number}; // @[Math.scala 450:32:@32743.4]
  assign _T_1395 = _GEN_0 << 1; // @[Math.scala 450:32:@32743.4]
  assign x507_rd_0_number = x386_lb_0_io_rPort_3_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 353:29:@32073.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 357:406:@32096.4]
  assign _GEN_1 = {{1'd0}, x507_rd_0_number}; // @[Math.scala 450:32:@32748.4]
  assign _T_1399 = _GEN_1 << 1; // @[Math.scala 450:32:@32748.4]
  assign x514_rd_0_number = x386_lb_0_io_rPort_2_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 368:29:@32124.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 372:406:@32147.4]
  assign _GEN_2 = {{2'd0}, x514_rd_0_number}; // @[Math.scala 450:32:@32753.4]
  assign _T_1403 = _GEN_2 << 2; // @[Math.scala 450:32:@32753.4]
  assign x521_rd_0_number = x386_lb_0_io_rPort_11_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 383:29:@32175.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 387:406:@32198.4]
  assign _GEN_3 = {{1'd0}, x521_rd_0_number}; // @[Math.scala 450:32:@32758.4]
  assign _T_1407 = _GEN_3 << 1; // @[Math.scala 450:32:@32758.4]
  assign x562_rd_0_number = x386_lb_0_io_rPort_7_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 482:29:@32509.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 486:406:@32532.4]
  assign _GEN_4 = {{1'd0}, x562_rd_0_number}; // @[Math.scala 450:32:@32763.4]
  assign _T_1411 = _GEN_4 << 1; // @[Math.scala 450:32:@32763.4]
  assign x604_sum_number = x604_sum_1_io_result; // @[Math.scala 154:22:@32852.4 Math.scala 155:14:@32853.4]
  assign _T_1447 = x604_sum_number[7:4]; // @[FixedPoint.scala 18:52:@32858.4]
  assign x462_rd_0_number = x386_lb_0_io_rPort_10_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 253:29:@31718.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 257:336:@31741.4]
  assign _GEN_5 = {{1'd0}, x462_rd_0_number}; // @[Math.scala 450:32:@32871.4]
  assign _T_1454 = _GEN_5 << 1; // @[Math.scala 450:32:@32871.4]
  assign _GEN_6 = {{1'd0}, x514_rd_0_number}; // @[Math.scala 450:32:@32876.4]
  assign _T_1458 = _GEN_6 << 1; // @[Math.scala 450:32:@32876.4]
  assign _GEN_7 = {{2'd0}, x521_rd_0_number}; // @[Math.scala 450:32:@32881.4]
  assign _T_1462 = _GEN_7 << 2; // @[Math.scala 450:32:@32881.4]
  assign x528_rd_0_number = x386_lb_0_io_rPort_16_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 402:29:@32244.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 406:406:@32267.4]
  assign _GEN_8 = {{1'd0}, x528_rd_0_number}; // @[Math.scala 450:32:@32886.4]
  assign _T_1466 = _GEN_8 << 1; // @[Math.scala 450:32:@32886.4]
  assign x569_rd_0_number = x386_lb_0_io_rPort_6_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 497:29:@32560.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 501:406:@32583.4]
  assign _GEN_9 = {{1'd0}, x569_rd_0_number}; // @[Math.scala 450:32:@32891.4]
  assign _T_1470 = _GEN_9 << 1; // @[Math.scala 450:32:@32891.4]
  assign x618_sum_number = x618_sum_1_io_result; // @[Math.scala 154:22:@32980.4 Math.scala 155:14:@32981.4]
  assign _T_1506 = x618_sum_number[7:4]; // @[FixedPoint.scala 18:52:@32986.4]
  assign x470_rd_0_number = x386_lb_0_io_rPort_12_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 276:29:@31803.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 280:336:@31826.4]
  assign _GEN_10 = {{1'd0}, x470_rd_0_number}; // @[Math.scala 450:32:@32999.4]
  assign _T_1513 = _GEN_10 << 1; // @[Math.scala 450:32:@32999.4]
  assign _GEN_11 = {{2'd0}, x528_rd_0_number}; // @[Math.scala 450:32:@33004.4]
  assign _T_1517 = _GEN_11 << 2; // @[Math.scala 450:32:@33004.4]
  assign x535_rd_0_number = x386_lb_0_io_rPort_9_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 417:29:@32295.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 421:406:@32318.4]
  assign _GEN_12 = {{1'd0}, x535_rd_0_number}; // @[Math.scala 450:32:@33009.4]
  assign _T_1521 = _GEN_12 << 1; // @[Math.scala 450:32:@33009.4]
  assign x576_rd_0_number = x386_lb_0_io_rPort_13_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 512:29:@32611.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 516:406:@32634.4]
  assign _GEN_13 = {{1'd0}, x576_rd_0_number}; // @[Math.scala 450:32:@33014.4]
  assign _T_1525 = _GEN_13 << 1; // @[Math.scala 450:32:@33014.4]
  assign x631_sum_number = x631_sum_1_io_result; // @[Math.scala 154:22:@33103.4 Math.scala 155:14:@33104.4]
  assign _T_1561 = x631_sum_number[7:4]; // @[FixedPoint.scala 18:52:@33109.4]
  assign x482_rd_0_number = x386_lb_0_io_rPort_15_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 303:29:@31882.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 307:406:@31905.4]
  assign _GEN_14 = {{1'd0}, x482_rd_0_number}; // @[Math.scala 450:32:@33122.4]
  assign _T_1568 = _GEN_14 << 1; // @[Math.scala 450:32:@33122.4]
  assign _GEN_15 = {{2'd0}, x535_rd_0_number}; // @[Math.scala 450:32:@33127.4]
  assign _T_1572 = _GEN_15 << 2; // @[Math.scala 450:32:@33127.4]
  assign x542_rd_0_number = x386_lb_0_io_rPort_1_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 440:29:@32348.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 444:406:@32371.4]
  assign _GEN_16 = {{1'd0}, x542_rd_0_number}; // @[Math.scala 450:32:@33132.4]
  assign _T_1576 = _GEN_16 << 1; // @[Math.scala 450:32:@33132.4]
  assign x583_rd_0_number = x386_lb_0_io_rPort_4_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 527:29:@32662.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 531:406:@32685.4]
  assign _GEN_17 = {{1'd0}, x583_rd_0_number}; // @[Math.scala 450:32:@33137.4]
  assign _T_1580 = _GEN_17 << 1; // @[Math.scala 450:32:@33137.4]
  assign x644_sum_number = x644_sum_1_io_result; // @[Math.scala 154:22:@33228.4 Math.scala 155:14:@33229.4]
  assign _T_1618 = x644_sum_number[7:4]; // @[FixedPoint.scala 18:52:@33234.4]
  assign _T_1643 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@33291.4 package.scala 96:25:@33292.4]
  assign _T_1645 = io_rr ? _T_1643 : 1'h0; // @[implicits.scala 55:10:@33293.4]
  assign _T_1646 = _T_360 & _T_1645; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:167:@33294.4]
  assign _T_1648 = _T_1646 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:255:@33296.4]
  assign _T_1649 = _T_1648 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:274:@33297.4]
  assign x830_b384_D12 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@33260.4 package.scala 96:25:@33261.4]
  assign _T_1650 = _T_1649 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 694:300:@33298.4]
  assign x829_b385_D12 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@33251.4 package.scala 96:25:@33252.4]
  assign _T_1664 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@33325.4 package.scala 96:25:@33326.4]
  assign _T_1666 = io_rr ? _T_1664 : 1'h0; // @[implicits.scala 55:10:@33327.4]
  assign _T_1667 = _T_360 & _T_1666; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:167:@33328.4]
  assign _T_1669 = _T_1667 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:255:@33330.4]
  assign _T_1670 = _T_1669 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:274:@33331.4]
  assign _T_1671 = _T_1670 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 701:300:@33332.4]
  assign _T_1685 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@33359.4 package.scala 96:25:@33360.4]
  assign _T_1687 = io_rr ? _T_1685 : 1'h0; // @[implicits.scala 55:10:@33361.4]
  assign _T_1688 = _T_360 & _T_1687; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:167:@33362.4]
  assign _T_1690 = _T_1688 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:255:@33364.4]
  assign _T_1691 = _T_1690 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:274:@33365.4]
  assign _T_1692 = _T_1691 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 708:300:@33366.4]
  assign _T_1706 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@33393.4 package.scala 96:25:@33394.4]
  assign _T_1708 = io_rr ? _T_1706 : 1'h0; // @[implicits.scala 55:10:@33395.4]
  assign _T_1709 = _T_360 & _T_1708; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:167:@33396.4]
  assign _T_1711 = _T_1709 & _T_360; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:255:@33398.4]
  assign _T_1712 = _T_1711 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:274:@33399.4]
  assign _T_1713 = _T_1712 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 715:300:@33400.4]
  assign _T_1739 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@33446.4 package.scala 96:25:@33447.4]
  assign _T_1741 = io_rr ? _T_1739 : 1'h0; // @[implicits.scala 55:10:@33448.4]
  assign _T_1742 = _T_360 & _T_1741; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 727:195:@33449.4]
  assign x837_x439_D5 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@33423.4 package.scala 96:25:@33424.4]
  assign _T_1743 = _T_1742 & x837_x439_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 727:283:@33450.4]
  assign _T_1744 = _T_1743 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 727:291:@33451.4]
  assign _T_1768 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@33490.4 package.scala 96:25:@33491.4]
  assign _T_1770 = io_rr ? _T_1768 : 1'h0; // @[implicits.scala 55:10:@33492.4]
  assign _T_1771 = _T_360 & _T_1770; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:195:@33493.4]
  assign x840_x450_D5 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@33476.4 package.scala 96:25:@33477.4]
  assign _T_1772 = _T_1771 & x840_x450_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:283:@33494.4]
  assign _T_1773 = _T_1772 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:291:@33495.4]
  assign _T_1797 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@33534.4 package.scala 96:25:@33535.4]
  assign _T_1799 = io_rr ? _T_1797 : 1'h0; // @[implicits.scala 55:10:@33536.4]
  assign _T_1800 = _T_360 & _T_1799; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:195:@33537.4]
  assign x841_x458_D5 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@33511.4 package.scala 96:25:@33512.4]
  assign _T_1801 = _T_1800 & x841_x458_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:283:@33538.4]
  assign _T_1802 = _T_1801 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:291:@33539.4]
  assign _T_1826 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@33578.4 package.scala 96:25:@33579.4]
  assign _T_1828 = io_rr ? _T_1826 : 1'h0; // @[implicits.scala 55:10:@33580.4]
  assign _T_1829 = _T_360 & _T_1828; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:195:@33581.4]
  assign x844_x466_D6 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@33564.4 package.scala 96:25:@33565.4]
  assign _T_1830 = _T_1829 & x844_x466_D6; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:283:@33582.4]
  assign _T_1831 = _T_1830 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:291:@33583.4]
  assign _T_1855 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@33622.4 package.scala 96:25:@33623.4]
  assign _T_1857 = io_rr ? _T_1855 : 1'h0; // @[implicits.scala 55:10:@33624.4]
  assign _T_1858 = _T_360 & _T_1857; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:195:@33625.4]
  assign x845_x475_D5 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@33599.4 package.scala 96:25:@33600.4]
  assign _T_1859 = _T_1858 & x845_x475_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:283:@33626.4]
  assign _T_1860 = _T_1859 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:291:@33627.4]
  assign _T_1887 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@33675.4 package.scala 96:25:@33676.4]
  assign _T_1889 = io_rr ? _T_1887 : 1'h0; // @[implicits.scala 55:10:@33677.4]
  assign _T_1890 = _T_360 & _T_1889; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:195:@33678.4]
  assign x847_x500_D5 = RetimeWrapper_107_io_out; // @[package.scala 96:25:@33643.4 package.scala 96:25:@33644.4]
  assign _T_1891 = _T_1890 & x847_x500_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:283:@33679.4]
  assign _T_1892 = _T_1891 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:291:@33680.4]
  assign _T_1916 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@33719.4 package.scala 96:25:@33720.4]
  assign _T_1918 = io_rr ? _T_1916 : 1'h0; // @[implicits.scala 55:10:@33721.4]
  assign _T_1919 = _T_360 & _T_1918; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:195:@33722.4]
  assign x851_x510_D5 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@33705.4 package.scala 96:25:@33706.4]
  assign _T_1920 = _T_1919 & x851_x510_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:283:@33723.4]
  assign _T_1921 = _T_1920 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:291:@33724.4]
  assign _T_1945 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@33763.4 package.scala 96:25:@33764.4]
  assign _T_1947 = io_rr ? _T_1945 : 1'h0; // @[implicits.scala 55:10:@33765.4]
  assign _T_1948 = _T_360 & _T_1947; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:195:@33766.4]
  assign x853_x517_D5 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@33749.4 package.scala 96:25:@33750.4]
  assign _T_1949 = _T_1948 & x853_x517_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:283:@33767.4]
  assign _T_1950 = _T_1949 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:291:@33768.4]
  assign _T_1974 = RetimeWrapper_119_io_out; // @[package.scala 96:25:@33807.4 package.scala 96:25:@33808.4]
  assign _T_1976 = io_rr ? _T_1974 : 1'h0; // @[implicits.scala 55:10:@33809.4]
  assign _T_1977 = _T_360 & _T_1976; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:195:@33810.4]
  assign x855_x524_D5 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@33793.4 package.scala 96:25:@33794.4]
  assign _T_1978 = _T_1977 & x855_x524_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:283:@33811.4]
  assign _T_1979 = _T_1978 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:291:@33812.4]
  assign _T_2003 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@33851.4 package.scala 96:25:@33852.4]
  assign _T_2005 = io_rr ? _T_2003 : 1'h0; // @[implicits.scala 55:10:@33853.4]
  assign _T_2006 = _T_360 & _T_2005; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 834:195:@33854.4]
  assign x856_x531_D5 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@33828.4 package.scala 96:25:@33829.4]
  assign _T_2007 = _T_2006 & x856_x531_D5; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 834:283:@33855.4]
  assign _T_2008 = _T_2007 & x830_b384_D12; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 834:291:@33856.4]
  assign x654_rd_0_number = x387_lb2_0_io_rPort_3_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 734:29:@33479.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 738:338:@33502.4]
  assign _GEN_18 = {{1'd0}, x654_rd_0_number}; // @[Math.scala 450:32:@33870.4]
  assign _T_2016 = _GEN_18 << 1; // @[Math.scala 450:32:@33870.4]
  assign x662_rd_0_number = x387_lb2_0_io_rPort_4_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 780:29:@33664.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 784:338:@33687.4]
  assign _GEN_19 = {{1'd0}, x662_rd_0_number}; // @[Math.scala 450:32:@33875.4]
  assign _T_2020 = _GEN_19 << 1; // @[Math.scala 450:32:@33875.4]
  assign x656_rd_0_number = x387_lb2_0_io_rPort_7_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 745:29:@33523.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 749:338:@33546.4]
  assign _GEN_20 = {{1'd0}, x656_rd_0_number}; // @[Math.scala 450:32:@33922.4]
  assign _T_2040 = _GEN_20 << 1; // @[Math.scala 450:32:@33922.4]
  assign x664_rd_0_number = x387_lb2_0_io_rPort_9_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 797:29:@33708.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 801:408:@33731.4]
  assign _GEN_21 = {{1'd0}, x664_rd_0_number}; // @[Math.scala 450:32:@33927.4]
  assign _T_2044 = _GEN_21 << 1; // @[Math.scala 450:32:@33927.4]
  assign x658_rd_0_number = x387_lb2_0_io_rPort_6_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 756:29:@33567.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 760:338:@33590.4]
  assign _GEN_22 = {{1'd0}, x658_rd_0_number}; // @[Math.scala 450:32:@33974.4]
  assign _T_2064 = _GEN_22 << 1; // @[Math.scala 450:32:@33974.4]
  assign x666_rd_0_number = x387_lb2_0_io_rPort_0_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 808:29:@33752.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 812:408:@33775.4]
  assign _GEN_23 = {{1'd0}, x666_rd_0_number}; // @[Math.scala 450:32:@33979.4]
  assign _T_2068 = _GEN_23 << 1; // @[Math.scala 450:32:@33979.4]
  assign x660_rd_0_number = x387_lb2_0_io_rPort_2_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 767:29:@33611.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 771:338:@33634.4]
  assign _GEN_24 = {{1'd0}, x660_rd_0_number}; // @[Math.scala 450:32:@34026.4]
  assign _T_2088 = _GEN_24 << 1; // @[Math.scala 450:32:@34026.4]
  assign x668_rd_0_number = x387_lb2_0_io_rPort_5_output_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 819:29:@33796.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 823:408:@33819.4]
  assign _GEN_25 = {{1'd0}, x668_rd_0_number}; // @[Math.scala 450:32:@34031.4]
  assign _T_2092 = _GEN_25 << 1; // @[Math.scala 450:32:@34031.4]
  assign x689_div_number = x689_div_1_io_result; // @[Math.scala 331:22:@34021.4 Math.scala 332:14:@34022.4]
  assign x695_div_number = x695_div_1_io_result; // @[Math.scala 331:22:@34073.4 Math.scala 332:14:@34074.4]
  assign _T_2120 = {x689_div_number,x695_div_number}; // @[Cat.scala 30:58:@34082.4]
  assign x677_div_number = x677_div_1_io_result; // @[Math.scala 331:22:@33917.4 Math.scala 332:14:@33918.4]
  assign x683_div_number = x683_div_1_io_result; // @[Math.scala 331:22:@33969.4 Math.scala 332:14:@33970.4]
  assign _T_2121 = {x677_div_number,x683_div_number}; // @[Cat.scala 30:58:@34083.4]
  assign _T_2134 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@34119.4 package.scala 96:25:@34120.4]
  assign _T_2136 = io_rr ? _T_2134 : 1'h0; // @[implicits.scala 55:10:@34121.4]
  assign x858_b384_D22 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@34101.4 package.scala 96:25:@34102.4]
  assign _T_2137 = _T_2136 & x858_b384_D22; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 896:116:@34122.4]
  assign x859_b385_D22 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@34110.4 package.scala 96:25:@34111.4]
  assign _T_2138 = _T_2137 & x859_b385_D22; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 896:122:@34123.4]
  assign x779_x768_D4_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31148.4 package.scala 96:25:@31149.4]
  assign x780_x401_sum_D3_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@31157.4 package.scala 96:25:@31158.4]
  assign x783_x411_sum_D2_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@31242.4 package.scala 96:25:@31243.4]
  assign x785_x420_sum_D2_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@31318.4 package.scala 96:25:@31319.4]
  assign x786_x429_sum_D2_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@31385.4 package.scala 96:25:@31386.4]
  assign x442_sum_number = x442_sum_1_io_result; // @[Math.scala 154:22:@31527.4 Math.scala 155:14:@31528.4]
  assign x795_x770_D2_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@31554.4 package.scala 96:25:@31555.4]
  assign x451_sum_number = x451_sum_1_io_result; // @[Math.scala 154:22:@31630.4 Math.scala 155:14:@31631.4]
  assign x459_sum_number = x459_sum_1_io_result; // @[Math.scala 154:22:@31706.4 Math.scala 155:14:@31707.4]
  assign x805_x467_sum_D1_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@31791.4 package.scala 96:25:@31792.4]
  assign x478_sum_number = x478_sum_1_io_result; // @[Math.scala 154:22:@31870.4 Math.scala 155:14:@31871.4]
  assign x490_sum_number = x490_sum_1_io_result; // @[Math.scala 154:22:@31951.4 Math.scala 155:14:@31952.4]
  assign x503_sum_number = x503_sum_1_io_result; // @[Math.scala 154:22:@32052.4 Math.scala 155:14:@32053.4]
  assign x810_x772_D1_number = RetimeWrapper_45_io_out; // @[package.scala 96:25:@32070.4 package.scala 96:25:@32071.4]
  assign x511_sum_number = x511_sum_1_io_result; // @[Math.scala 154:22:@32112.4 Math.scala 155:14:@32113.4]
  assign x518_sum_number = x518_sum_1_io_result; // @[Math.scala 154:22:@32163.4 Math.scala 155:14:@32164.4]
  assign x525_sum_number = x525_sum_1_io_result; // @[Math.scala 154:22:@32232.4 Math.scala 155:14:@32233.4]
  assign x532_sum_number = x532_sum_1_io_result; // @[Math.scala 154:22:@32283.4 Math.scala 155:14:@32284.4]
  assign x539_sum_number = x539_sum_1_io_result; // @[Math.scala 154:22:@32336.4 Math.scala 155:14:@32337.4]
  assign x551_sum_number = x551_sum_1_io_result; // @[Math.scala 154:22:@32437.4 Math.scala 155:14:@32438.4]
  assign x818_x774_D1_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@32446.4 package.scala 96:25:@32447.4]
  assign x559_sum_number = x559_sum_1_io_result; // @[Math.scala 154:22:@32497.4 Math.scala 155:14:@32498.4]
  assign x566_sum_number = x566_sum_1_io_result; // @[Math.scala 154:22:@32548.4 Math.scala 155:14:@32549.4]
  assign x573_sum_number = x573_sum_1_io_result; // @[Math.scala 154:22:@32599.4 Math.scala 155:14:@32600.4]
  assign x580_sum_number = x580_sum_1_io_result; // @[Math.scala 154:22:@32650.4 Math.scala 155:14:@32651.4]
  assign x587_sum_number = x587_sum_1_io_result; // @[Math.scala 154:22:@32701.4 Math.scala 155:14:@32702.4]
  assign x831_x768_D12_number = RetimeWrapper_82_io_out; // @[package.scala 96:25:@33269.4 package.scala 96:25:@33270.4]
  assign x832_x401_sum_D11_number = RetimeWrapper_83_io_out; // @[package.scala 96:25:@33278.4 package.scala 96:25:@33279.4]
  assign x833_x411_sum_D10_number = RetimeWrapper_85_io_out; // @[package.scala 96:25:@33312.4 package.scala 96:25:@33313.4]
  assign x834_x420_sum_D10_number = RetimeWrapper_87_io_out; // @[package.scala 96:25:@33346.4 package.scala 96:25:@33347.4]
  assign x835_x429_sum_D10_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@33380.4 package.scala 96:25:@33381.4]
  assign x836_x770_D6_number = RetimeWrapper_91_io_out; // @[package.scala 96:25:@33414.4 package.scala 96:25:@33415.4]
  assign x838_x442_sum_D4_number = RetimeWrapper_93_io_out; // @[package.scala 96:25:@33432.4 package.scala 96:25:@33433.4]
  assign x839_x451_sum_D4_number = RetimeWrapper_95_io_out; // @[package.scala 96:25:@33467.4 package.scala 96:25:@33468.4]
  assign x842_x459_sum_D4_number = RetimeWrapper_99_io_out; // @[package.scala 96:25:@33520.4 package.scala 96:25:@33521.4]
  assign x843_x467_sum_D5_number = RetimeWrapper_101_io_out; // @[package.scala 96:25:@33555.4 package.scala 96:25:@33556.4]
  assign x846_x478_sum_D4_number = RetimeWrapper_105_io_out; // @[package.scala 96:25:@33608.4 package.scala 96:25:@33609.4]
  assign x848_x503_sum_D4_number = RetimeWrapper_108_io_out; // @[package.scala 96:25:@33652.4 package.scala 96:25:@33653.4]
  assign x849_x772_D5_number = RetimeWrapper_109_io_out; // @[package.scala 96:25:@33661.4 package.scala 96:25:@33662.4]
  assign x850_x511_sum_D4_number = RetimeWrapper_111_io_out; // @[package.scala 96:25:@33696.4 package.scala 96:25:@33697.4]
  assign x852_x518_sum_D4_number = RetimeWrapper_114_io_out; // @[package.scala 96:25:@33740.4 package.scala 96:25:@33741.4]
  assign x854_x525_sum_D4_number = RetimeWrapper_117_io_out; // @[package.scala 96:25:@33784.4 package.scala 96:25:@33785.4]
  assign x857_x532_sum_D4_number = RetimeWrapper_121_io_out; // @[package.scala 96:25:@33837.4 package.scala 96:25:@33838.4]
  assign io_in_x374_TVALID = _T_2138 & io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 896:22:@34125.4]
  assign io_in_x374_TDATA = {{224'd0}, RetimeWrapper_123_io_out}; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 897:24:@34126.4]
  assign io_in_x373_TREADY = _T_213 & _T_215; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 69:22:@30996.4 sm_x700_inr_Foreach_SAMPLER_BOX.scala 71:22:@31004.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@30732.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@30744.4]
  assign x386_lb_0_clock = clock; // @[:@30752.4]
  assign x386_lb_0_reset = reset; // @[:@30753.4]
  assign x386_lb_0_io_rPort_17_banks_0 = x795_x770_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@31660.4]
  assign x386_lb_0_io_rPort_17_ofs_0 = x451_sum_number[0]; // @[MemInterfaceType.scala 107:54:@31662.4]
  assign x386_lb_0_io_rPort_17_en_0 = _T_664 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@31664.4]
  assign x386_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31663.4]
  assign x386_lb_0_io_rPort_16_banks_0 = x810_x772_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32262.4]
  assign x386_lb_0_io_rPort_16_ofs_0 = x525_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32264.4]
  assign x386_lb_0_io_rPort_16_en_0 = _T_1069 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32266.4]
  assign x386_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32265.4]
  assign x386_lb_0_io_rPort_15_banks_0 = x795_x770_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@31900.4]
  assign x386_lb_0_io_rPort_15_ofs_0 = x478_sum_number[0]; // @[MemInterfaceType.scala 107:54:@31902.4]
  assign x386_lb_0_io_rPort_15_en_0 = _T_819 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@31904.4]
  assign x386_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31903.4]
  assign x386_lb_0_io_rPort_14_banks_0 = x795_x770_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@31584.4]
  assign x386_lb_0_io_rPort_14_ofs_0 = x442_sum_number[0]; // @[MemInterfaceType.scala 107:54:@31586.4]
  assign x386_lb_0_io_rPort_14_en_0 = _T_617 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@31588.4]
  assign x386_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31587.4]
  assign x386_lb_0_io_rPort_13_banks_0 = x818_x774_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32629.4]
  assign x386_lb_0_io_rPort_13_ofs_0 = x573_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32631.4]
  assign x386_lb_0_io_rPort_13_en_0 = _T_1321 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32633.4]
  assign x386_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32632.4]
  assign x386_lb_0_io_rPort_12_banks_0 = x795_x770_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@31821.4]
  assign x386_lb_0_io_rPort_12_ofs_0 = x805_x467_sum_D1_number[0]; // @[MemInterfaceType.scala 107:54:@31823.4]
  assign x386_lb_0_io_rPort_12_en_0 = _T_761 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@31825.4]
  assign x386_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31824.4]
  assign x386_lb_0_io_rPort_11_banks_0 = x810_x772_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32193.4]
  assign x386_lb_0_io_rPort_11_ofs_0 = x518_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32195.4]
  assign x386_lb_0_io_rPort_11_en_0 = _T_1030 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32197.4]
  assign x386_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32196.4]
  assign x386_lb_0_io_rPort_10_banks_0 = x795_x770_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@31736.4]
  assign x386_lb_0_io_rPort_10_ofs_0 = x459_sum_number[0]; // @[MemInterfaceType.scala 107:54:@31738.4]
  assign x386_lb_0_io_rPort_10_en_0 = _T_711 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@31740.4]
  assign x386_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31739.4]
  assign x386_lb_0_io_rPort_9_banks_0 = x810_x772_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32313.4]
  assign x386_lb_0_io_rPort_9_ofs_0 = x532_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32315.4]
  assign x386_lb_0_io_rPort_9_en_0 = _T_1102 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32317.4]
  assign x386_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32316.4]
  assign x386_lb_0_io_rPort_8_banks_0 = x795_x770_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@31981.4]
  assign x386_lb_0_io_rPort_8_ofs_0 = x490_sum_number[0]; // @[MemInterfaceType.scala 107:54:@31983.4]
  assign x386_lb_0_io_rPort_8_en_0 = _T_879 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@31985.4]
  assign x386_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@31984.4]
  assign x386_lb_0_io_rPort_7_banks_0 = x818_x774_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32527.4]
  assign x386_lb_0_io_rPort_7_ofs_0 = x559_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32529.4]
  assign x386_lb_0_io_rPort_7_en_0 = _T_1255 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32531.4]
  assign x386_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32530.4]
  assign x386_lb_0_io_rPort_6_banks_0 = x818_x774_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32578.4]
  assign x386_lb_0_io_rPort_6_ofs_0 = x566_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32580.4]
  assign x386_lb_0_io_rPort_6_en_0 = _T_1288 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32582.4]
  assign x386_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32581.4]
  assign x386_lb_0_io_rPort_5_banks_0 = x818_x774_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32731.4]
  assign x386_lb_0_io_rPort_5_ofs_0 = x587_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32733.4]
  assign x386_lb_0_io_rPort_5_en_0 = _T_1387 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32735.4]
  assign x386_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32734.4]
  assign x386_lb_0_io_rPort_4_banks_0 = x818_x774_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32680.4]
  assign x386_lb_0_io_rPort_4_ofs_0 = x580_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32682.4]
  assign x386_lb_0_io_rPort_4_en_0 = _T_1354 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32684.4]
  assign x386_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32683.4]
  assign x386_lb_0_io_rPort_3_banks_0 = x810_x772_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32091.4]
  assign x386_lb_0_io_rPort_3_ofs_0 = x503_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32093.4]
  assign x386_lb_0_io_rPort_3_en_0 = _T_964 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32095.4]
  assign x386_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32094.4]
  assign x386_lb_0_io_rPort_2_banks_0 = x810_x772_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32142.4]
  assign x386_lb_0_io_rPort_2_ofs_0 = x511_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32144.4]
  assign x386_lb_0_io_rPort_2_en_0 = _T_997 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32146.4]
  assign x386_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32145.4]
  assign x386_lb_0_io_rPort_1_banks_0 = x810_x772_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32366.4]
  assign x386_lb_0_io_rPort_1_ofs_0 = x539_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32368.4]
  assign x386_lb_0_io_rPort_1_en_0 = _T_1137 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32370.4]
  assign x386_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32369.4]
  assign x386_lb_0_io_rPort_0_banks_0 = x818_x774_D1_number[2:0]; // @[MemInterfaceType.scala 106:58:@32476.4]
  assign x386_lb_0_io_rPort_0_ofs_0 = x551_sum_number[0]; // @[MemInterfaceType.scala 107:54:@32478.4]
  assign x386_lb_0_io_rPort_0_en_0 = _T_1222 & x793_b385_D8; // @[MemInterfaceType.scala 110:79:@32480.4]
  assign x386_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32479.4]
  assign x386_lb_0_io_wPort_3_banks_0 = x779_x768_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@31416.4]
  assign x386_lb_0_io_wPort_3_ofs_0 = x786_x429_sum_D2_number[0]; // @[MemInterfaceType.scala 89:54:@31418.4]
  assign x386_lb_0_io_wPort_3_data_0 = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 90:56:@31419.4]
  assign x386_lb_0_io_wPort_3_en_0 = _T_509 & x776_b385_D4; // @[MemInterfaceType.scala 93:57:@31421.4]
  assign x386_lb_0_io_wPort_2_banks_0 = x779_x768_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@31340.4]
  assign x386_lb_0_io_wPort_2_ofs_0 = x785_x420_sum_D2_number[0]; // @[MemInterfaceType.scala 89:54:@31342.4]
  assign x386_lb_0_io_wPort_2_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@31343.4]
  assign x386_lb_0_io_wPort_2_en_0 = _T_464 & x776_b385_D4; // @[MemInterfaceType.scala 93:57:@31345.4]
  assign x386_lb_0_io_wPort_1_banks_0 = x779_x768_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@31264.4]
  assign x386_lb_0_io_wPort_1_ofs_0 = x783_x411_sum_D2_number[0]; // @[MemInterfaceType.scala 89:54:@31266.4]
  assign x386_lb_0_io_wPort_1_data_0 = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 90:56:@31267.4]
  assign x386_lb_0_io_wPort_1_en_0 = _T_419 & x776_b385_D4; // @[MemInterfaceType.scala 93:57:@31269.4]
  assign x386_lb_0_io_wPort_0_banks_0 = x779_x768_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@31179.4]
  assign x386_lb_0_io_wPort_0_ofs_0 = x780_x401_sum_D3_number[0]; // @[MemInterfaceType.scala 89:54:@31181.4]
  assign x386_lb_0_io_wPort_0_data_0 = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 90:56:@31182.4]
  assign x386_lb_0_io_wPort_0_en_0 = _T_371 & x776_b385_D4; // @[MemInterfaceType.scala 93:57:@31184.4]
  assign x387_lb2_0_clock = clock; // @[:@30897.4]
  assign x387_lb2_0_reset = reset; // @[:@30898.4]
  assign x387_lb2_0_io_rPort_9_banks_0 = x849_x772_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@33726.4]
  assign x387_lb2_0_io_rPort_9_ofs_0 = x850_x511_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33728.4]
  assign x387_lb2_0_io_rPort_9_en_0 = _T_1921 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33730.4]
  assign x387_lb2_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33729.4]
  assign x387_lb2_0_io_rPort_8_banks_0 = x836_x770_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@33453.4]
  assign x387_lb2_0_io_rPort_8_ofs_0 = x838_x442_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33455.4]
  assign x387_lb2_0_io_rPort_8_en_0 = _T_1744 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33457.4]
  assign x387_lb2_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33456.4]
  assign x387_lb2_0_io_rPort_7_banks_0 = x836_x770_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@33541.4]
  assign x387_lb2_0_io_rPort_7_ofs_0 = x842_x459_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33543.4]
  assign x387_lb2_0_io_rPort_7_en_0 = _T_1802 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33545.4]
  assign x387_lb2_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33544.4]
  assign x387_lb2_0_io_rPort_6_banks_0 = x836_x770_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@33585.4]
  assign x387_lb2_0_io_rPort_6_ofs_0 = x843_x467_sum_D5_number[0]; // @[MemInterfaceType.scala 107:54:@33587.4]
  assign x387_lb2_0_io_rPort_6_en_0 = _T_1831 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33589.4]
  assign x387_lb2_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33588.4]
  assign x387_lb2_0_io_rPort_5_banks_0 = x849_x772_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@33814.4]
  assign x387_lb2_0_io_rPort_5_ofs_0 = x854_x525_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33816.4]
  assign x387_lb2_0_io_rPort_5_en_0 = _T_1979 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33818.4]
  assign x387_lb2_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33817.4]
  assign x387_lb2_0_io_rPort_4_banks_0 = x849_x772_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@33682.4]
  assign x387_lb2_0_io_rPort_4_ofs_0 = x848_x503_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33684.4]
  assign x387_lb2_0_io_rPort_4_en_0 = _T_1892 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33686.4]
  assign x387_lb2_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33685.4]
  assign x387_lb2_0_io_rPort_3_banks_0 = x836_x770_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@33497.4]
  assign x387_lb2_0_io_rPort_3_ofs_0 = x839_x451_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33499.4]
  assign x387_lb2_0_io_rPort_3_en_0 = _T_1773 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33501.4]
  assign x387_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33500.4]
  assign x387_lb2_0_io_rPort_2_banks_0 = x836_x770_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@33629.4]
  assign x387_lb2_0_io_rPort_2_ofs_0 = x846_x478_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33631.4]
  assign x387_lb2_0_io_rPort_2_en_0 = _T_1860 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33633.4]
  assign x387_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33632.4]
  assign x387_lb2_0_io_rPort_1_banks_0 = x849_x772_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@33858.4]
  assign x387_lb2_0_io_rPort_1_ofs_0 = x857_x532_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33860.4]
  assign x387_lb2_0_io_rPort_1_en_0 = _T_2008 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33862.4]
  assign x387_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33861.4]
  assign x387_lb2_0_io_rPort_0_banks_0 = x849_x772_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@33770.4]
  assign x387_lb2_0_io_rPort_0_ofs_0 = x852_x518_sum_D4_number[0]; // @[MemInterfaceType.scala 107:54:@33772.4]
  assign x387_lb2_0_io_rPort_0_en_0 = _T_1950 & x829_b385_D12; // @[MemInterfaceType.scala 110:79:@33774.4]
  assign x387_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33773.4]
  assign x387_lb2_0_io_wPort_3_banks_0 = x831_x768_D12_number[2:0]; // @[MemInterfaceType.scala 88:58:@33402.4]
  assign x387_lb2_0_io_wPort_3_ofs_0 = x835_x429_sum_D10_number[0]; // @[MemInterfaceType.scala 89:54:@33404.4]
  assign x387_lb2_0_io_wPort_3_data_0 = RetimeWrapper_73_io_out; // @[MemInterfaceType.scala 90:56:@33405.4]
  assign x387_lb2_0_io_wPort_3_en_0 = _T_1713 & x829_b385_D12; // @[MemInterfaceType.scala 93:57:@33407.4]
  assign x387_lb2_0_io_wPort_2_banks_0 = x831_x768_D12_number[2:0]; // @[MemInterfaceType.scala 88:58:@33368.4]
  assign x387_lb2_0_io_wPort_2_ofs_0 = x834_x420_sum_D10_number[0]; // @[MemInterfaceType.scala 89:54:@33370.4]
  assign x387_lb2_0_io_wPort_2_data_0 = RetimeWrapper_75_io_out; // @[MemInterfaceType.scala 90:56:@33371.4]
  assign x387_lb2_0_io_wPort_2_en_0 = _T_1692 & x829_b385_D12; // @[MemInterfaceType.scala 93:57:@33373.4]
  assign x387_lb2_0_io_wPort_1_banks_0 = x831_x768_D12_number[2:0]; // @[MemInterfaceType.scala 88:58:@33334.4]
  assign x387_lb2_0_io_wPort_1_ofs_0 = x833_x411_sum_D10_number[0]; // @[MemInterfaceType.scala 89:54:@33336.4]
  assign x387_lb2_0_io_wPort_1_data_0 = RetimeWrapper_77_io_out; // @[MemInterfaceType.scala 90:56:@33337.4]
  assign x387_lb2_0_io_wPort_1_en_0 = _T_1671 & x829_b385_D12; // @[MemInterfaceType.scala 93:57:@33339.4]
  assign x387_lb2_0_io_wPort_0_banks_0 = x831_x768_D12_number[2:0]; // @[MemInterfaceType.scala 88:58:@33300.4]
  assign x387_lb2_0_io_wPort_0_ofs_0 = x832_x401_sum_D11_number[0]; // @[MemInterfaceType.scala 89:54:@33302.4]
  assign x387_lb2_0_io_wPort_0_data_0 = RetimeWrapper_79_io_out; // @[MemInterfaceType.scala 90:56:@33303.4]
  assign x387_lb2_0_io_wPort_0_en_0 = _T_1650 & x829_b385_D12; // @[MemInterfaceType.scala 93:57:@33305.4]
  assign RetimeWrapper_clock = clock; // @[:@31007.4]
  assign RetimeWrapper_reset = reset; // @[:@31008.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31010.4]
  assign RetimeWrapper_io_in = io_in_x373_TDATA[31:0]; // @[package.scala 94:16:@31009.4]
  assign x401_sum_1_clock = clock; // @[:@31107.4]
  assign x401_sum_1_reset = reset; // @[:@31108.4]
  assign x401_sum_1_io_a = {_T_324,_T_325}; // @[Math.scala 151:17:@31109.4]
  assign x401_sum_1_io_b = {_T_334,_T_335}; // @[Math.scala 152:17:@31110.4]
  assign x401_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31111.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31117.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31118.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31120.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@31119.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31126.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31127.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31129.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@31128.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31135.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31136.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31138.4]
  assign RetimeWrapper_3_io_in = x775_x388_D1_0_number[7:0]; // @[package.scala 94:16:@31137.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31144.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31145.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31147.4]
  assign RetimeWrapper_4_io_in = $unsigned(_T_315); // @[package.scala 94:16:@31146.4]
  assign RetimeWrapper_5_clock = clock; // @[:@31153.4]
  assign RetimeWrapper_5_reset = reset; // @[:@31154.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31156.4]
  assign RetimeWrapper_5_io_in = x401_sum_1_io_result; // @[package.scala 94:16:@31155.4]
  assign RetimeWrapper_6_clock = clock; // @[:@31166.4]
  assign RetimeWrapper_6_reset = reset; // @[:@31167.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31169.4]
  assign RetimeWrapper_6_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31168.4]
  assign x407_rdcol_1_clock = clock; // @[:@31189.4]
  assign x407_rdcol_1_reset = reset; // @[:@31190.4]
  assign x407_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@31191.4]
  assign x407_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@31192.4]
  assign x407_rdcol_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31193.4]
  assign RetimeWrapper_7_clock = clock; // @[:@31210.4]
  assign RetimeWrapper_7_reset = reset; // @[:@31211.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31213.4]
  assign RetimeWrapper_7_io_in = {_T_324,_T_325}; // @[package.scala 94:16:@31212.4]
  assign x411_sum_1_clock = clock; // @[:@31219.4]
  assign x411_sum_1_reset = reset; // @[:@31220.4]
  assign x411_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@31221.4]
  assign x411_sum_1_io_b = {_T_388,_T_389}; // @[Math.scala 152:17:@31222.4]
  assign x411_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31223.4]
  assign RetimeWrapper_8_clock = clock; // @[:@31229.4]
  assign RetimeWrapper_8_reset = reset; // @[:@31230.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31232.4]
  assign RetimeWrapper_8_io_in = x775_x388_D1_0_number[15:8]; // @[package.scala 94:16:@31231.4]
  assign RetimeWrapper_9_clock = clock; // @[:@31238.4]
  assign RetimeWrapper_9_reset = reset; // @[:@31239.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31241.4]
  assign RetimeWrapper_9_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@31240.4]
  assign RetimeWrapper_10_clock = clock; // @[:@31251.4]
  assign RetimeWrapper_10_reset = reset; // @[:@31252.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31254.4]
  assign RetimeWrapper_10_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31253.4]
  assign x416_rdcol_1_clock = clock; // @[:@31274.4]
  assign x416_rdcol_1_reset = reset; // @[:@31275.4]
  assign x416_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@31276.4]
  assign x416_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@31277.4]
  assign x416_rdcol_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31278.4]
  assign x420_sum_1_clock = clock; // @[:@31295.4]
  assign x420_sum_1_reset = reset; // @[:@31296.4]
  assign x420_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@31297.4]
  assign x420_sum_1_io_b = {_T_436,_T_437}; // @[Math.scala 152:17:@31298.4]
  assign x420_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31299.4]
  assign RetimeWrapper_11_clock = clock; // @[:@31305.4]
  assign RetimeWrapper_11_reset = reset; // @[:@31306.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31308.4]
  assign RetimeWrapper_11_io_in = x775_x388_D1_0_number[23:16]; // @[package.scala 94:16:@31307.4]
  assign RetimeWrapper_12_clock = clock; // @[:@31314.4]
  assign RetimeWrapper_12_reset = reset; // @[:@31315.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31317.4]
  assign RetimeWrapper_12_io_in = x420_sum_1_io_result; // @[package.scala 94:16:@31316.4]
  assign RetimeWrapper_13_clock = clock; // @[:@31327.4]
  assign RetimeWrapper_13_reset = reset; // @[:@31328.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31330.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31329.4]
  assign x425_rdcol_1_clock = clock; // @[:@31350.4]
  assign x425_rdcol_1_reset = reset; // @[:@31351.4]
  assign x425_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@31352.4]
  assign x425_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@31353.4]
  assign x425_rdcol_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31354.4]
  assign x429_sum_1_clock = clock; // @[:@31371.4]
  assign x429_sum_1_reset = reset; // @[:@31372.4]
  assign x429_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@31373.4]
  assign x429_sum_1_io_b = {_T_481,_T_482}; // @[Math.scala 152:17:@31374.4]
  assign x429_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31375.4]
  assign RetimeWrapper_14_clock = clock; // @[:@31381.4]
  assign RetimeWrapper_14_reset = reset; // @[:@31382.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31384.4]
  assign RetimeWrapper_14_io_in = x429_sum_1_io_result; // @[package.scala 94:16:@31383.4]
  assign RetimeWrapper_15_clock = clock; // @[:@31390.4]
  assign RetimeWrapper_15_reset = reset; // @[:@31391.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31393.4]
  assign RetimeWrapper_15_io_in = x775_x388_D1_0_number[31:24]; // @[package.scala 94:16:@31392.4]
  assign RetimeWrapper_16_clock = clock; // @[:@31403.4]
  assign RetimeWrapper_16_reset = reset; // @[:@31404.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31406.4]
  assign RetimeWrapper_16_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31405.4]
  assign RetimeWrapper_17_clock = clock; // @[:@31424.4]
  assign RetimeWrapper_17_reset = reset; // @[:@31425.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31427.4]
  assign RetimeWrapper_17_io_in = __io_result; // @[package.scala 94:16:@31426.4]
  assign RetimeWrapper_18_clock = clock; // @[:@31451.4]
  assign RetimeWrapper_18_reset = reset; // @[:@31452.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31454.4]
  assign RetimeWrapper_18_io_in = x425_rdcol_1_io_result; // @[package.scala 94:16:@31453.4]
  assign RetimeWrapper_19_clock = clock; // @[:@31469.4]
  assign RetimeWrapper_19_reset = reset; // @[:@31470.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31472.4]
  assign RetimeWrapper_19_io_in = $signed(_T_521) < $signed(32'sh0); // @[package.scala 94:16:@31471.4]
  assign RetimeWrapper_20_clock = clock; // @[:@31504.4]
  assign RetimeWrapper_20_reset = reset; // @[:@31505.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31507.4]
  assign RetimeWrapper_20_io_in = {_T_573,_T_574}; // @[package.scala 94:16:@31506.4]
  assign RetimeWrapper_21_clock = clock; // @[:@31513.4]
  assign RetimeWrapper_21_reset = reset; // @[:@31514.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31516.4]
  assign RetimeWrapper_21_io_in = {_T_481,_T_482}; // @[package.scala 94:16:@31515.4]
  assign x442_sum_1_clock = clock; // @[:@31522.4]
  assign x442_sum_1_reset = reset; // @[:@31523.4]
  assign x442_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@31524.4]
  assign x442_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@31525.4]
  assign x442_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31526.4]
  assign RetimeWrapper_22_clock = clock; // @[:@31532.4]
  assign RetimeWrapper_22_reset = reset; // @[:@31533.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31535.4]
  assign RetimeWrapper_22_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@31534.4]
  assign RetimeWrapper_23_clock = clock; // @[:@31541.4]
  assign RetimeWrapper_23_reset = reset; // @[:@31542.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31544.4]
  assign RetimeWrapper_23_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@31543.4]
  assign RetimeWrapper_24_clock = clock; // @[:@31550.4]
  assign RetimeWrapper_24_reset = reset; // @[:@31551.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31553.4]
  assign RetimeWrapper_24_io_in = $unsigned(_T_564); // @[package.scala 94:16:@31552.4]
  assign RetimeWrapper_25_clock = clock; // @[:@31559.4]
  assign RetimeWrapper_25_reset = reset; // @[:@31560.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31562.4]
  assign RetimeWrapper_25_io_in = ~ x438; // @[package.scala 94:16:@31561.4]
  assign RetimeWrapper_26_clock = clock; // @[:@31573.4]
  assign RetimeWrapper_26_reset = reset; // @[:@31574.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31576.4]
  assign RetimeWrapper_26_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31575.4]
  assign RetimeWrapper_27_clock = clock; // @[:@31594.4]
  assign RetimeWrapper_27_reset = reset; // @[:@31595.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31597.4]
  assign RetimeWrapper_27_io_in = x416_rdcol_1_io_result; // @[package.scala 94:16:@31596.4]
  assign RetimeWrapper_28_clock = clock; // @[:@31616.4]
  assign RetimeWrapper_28_reset = reset; // @[:@31617.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31619.4]
  assign RetimeWrapper_28_io_in = {_T_436,_T_437}; // @[package.scala 94:16:@31618.4]
  assign x451_sum_1_clock = clock; // @[:@31625.4]
  assign x451_sum_1_reset = reset; // @[:@31626.4]
  assign x451_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@31627.4]
  assign x451_sum_1_io_b = RetimeWrapper_28_io_out; // @[Math.scala 152:17:@31628.4]
  assign x451_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31629.4]
  assign RetimeWrapper_29_clock = clock; // @[:@31635.4]
  assign RetimeWrapper_29_reset = reset; // @[:@31636.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31638.4]
  assign RetimeWrapper_29_io_in = ~ x449; // @[package.scala 94:16:@31637.4]
  assign RetimeWrapper_30_clock = clock; // @[:@31649.4]
  assign RetimeWrapper_30_reset = reset; // @[:@31650.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31652.4]
  assign RetimeWrapper_30_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31651.4]
  assign RetimeWrapper_31_clock = clock; // @[:@31670.4]
  assign RetimeWrapper_31_reset = reset; // @[:@31671.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31673.4]
  assign RetimeWrapper_31_io_in = x407_rdcol_1_io_result; // @[package.scala 94:16:@31672.4]
  assign RetimeWrapper_32_clock = clock; // @[:@31692.4]
  assign RetimeWrapper_32_reset = reset; // @[:@31693.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31695.4]
  assign RetimeWrapper_32_io_in = {_T_388,_T_389}; // @[package.scala 94:16:@31694.4]
  assign x459_sum_1_clock = clock; // @[:@31701.4]
  assign x459_sum_1_reset = reset; // @[:@31702.4]
  assign x459_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@31703.4]
  assign x459_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@31704.4]
  assign x459_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31705.4]
  assign RetimeWrapper_33_clock = clock; // @[:@31711.4]
  assign RetimeWrapper_33_reset = reset; // @[:@31712.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31714.4]
  assign RetimeWrapper_33_io_in = ~ x457; // @[package.scala 94:16:@31713.4]
  assign RetimeWrapper_34_clock = clock; // @[:@31725.4]
  assign RetimeWrapper_34_reset = reset; // @[:@31726.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31728.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31727.4]
  assign RetimeWrapper_35_clock = clock; // @[:@31746.4]
  assign RetimeWrapper_35_reset = reset; // @[:@31747.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31749.4]
  assign RetimeWrapper_35_io_in = __1_io_result; // @[package.scala 94:16:@31748.4]
  assign RetimeWrapper_36_clock = clock; // @[:@31768.4]
  assign RetimeWrapper_36_reset = reset; // @[:@31769.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31771.4]
  assign RetimeWrapper_36_io_in = {_T_334,_T_335}; // @[package.scala 94:16:@31770.4]
  assign x467_sum_1_clock = clock; // @[:@31777.4]
  assign x467_sum_1_reset = reset; // @[:@31778.4]
  assign x467_sum_1_io_a = {_T_573,_T_574}; // @[Math.scala 151:17:@31779.4]
  assign x467_sum_1_io_b = RetimeWrapper_36_io_out; // @[Math.scala 152:17:@31780.4]
  assign x467_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31781.4]
  assign RetimeWrapper_37_clock = clock; // @[:@31787.4]
  assign RetimeWrapper_37_reset = reset; // @[:@31788.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31790.4]
  assign RetimeWrapper_37_io_in = x467_sum_1_io_result; // @[package.scala 94:16:@31789.4]
  assign RetimeWrapper_38_clock = clock; // @[:@31796.4]
  assign RetimeWrapper_38_reset = reset; // @[:@31797.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31799.4]
  assign RetimeWrapper_38_io_in = ~ x465; // @[package.scala 94:16:@31798.4]
  assign RetimeWrapper_39_clock = clock; // @[:@31810.4]
  assign RetimeWrapper_39_reset = reset; // @[:@31811.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31813.4]
  assign RetimeWrapper_39_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31812.4]
  assign x472_rdcol_1_clock = clock; // @[:@31833.4]
  assign x472_rdcol_1_reset = reset; // @[:@31834.4]
  assign x472_rdcol_1_io_a = RetimeWrapper_35_io_out; // @[Math.scala 151:17:@31835.4]
  assign x472_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@31836.4]
  assign x472_rdcol_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31837.4]
  assign x478_sum_1_clock = clock; // @[:@31865.4]
  assign x478_sum_1_reset = reset; // @[:@31866.4]
  assign x478_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@31867.4]
  assign x478_sum_1_io_b = {_T_790,_T_791}; // @[Math.scala 152:17:@31868.4]
  assign x478_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31869.4]
  assign RetimeWrapper_40_clock = clock; // @[:@31875.4]
  assign RetimeWrapper_40_reset = reset; // @[:@31876.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31878.4]
  assign RetimeWrapper_40_io_in = ~ x474; // @[package.scala 94:16:@31877.4]
  assign RetimeWrapper_41_clock = clock; // @[:@31889.4]
  assign RetimeWrapper_41_reset = reset; // @[:@31890.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31892.4]
  assign RetimeWrapper_41_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31891.4]
  assign x484_rdcol_1_clock = clock; // @[:@31914.4]
  assign x484_rdcol_1_reset = reset; // @[:@31915.4]
  assign x484_rdcol_1_io_a = RetimeWrapper_35_io_out; // @[Math.scala 151:17:@31916.4]
  assign x484_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@31917.4]
  assign x484_rdcol_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31918.4]
  assign x490_sum_1_clock = clock; // @[:@31946.4]
  assign x490_sum_1_reset = reset; // @[:@31947.4]
  assign x490_sum_1_io_a = RetimeWrapper_20_io_out; // @[Math.scala 151:17:@31948.4]
  assign x490_sum_1_io_b = {_T_850,_T_851}; // @[Math.scala 152:17:@31949.4]
  assign x490_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@31950.4]
  assign RetimeWrapper_42_clock = clock; // @[:@31956.4]
  assign RetimeWrapper_42_reset = reset; // @[:@31957.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31959.4]
  assign RetimeWrapper_42_io_in = ~ x486; // @[package.scala 94:16:@31958.4]
  assign RetimeWrapper_43_clock = clock; // @[:@31970.4]
  assign RetimeWrapper_43_reset = reset; // @[:@31971.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@31973.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@31972.4]
  assign x496_rdrow_1_clock = clock; // @[:@31993.4]
  assign x496_rdrow_1_reset = reset; // @[:@31994.4]
  assign x496_rdrow_1_io_a = RetimeWrapper_17_io_out; // @[Math.scala 192:17:@31995.4]
  assign x496_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@31996.4]
  assign x496_rdrow_1_io_flow = io_in_x374_TREADY; // @[Math.scala 194:20:@31997.4]
  assign x503_sum_1_clock = clock; // @[:@32047.4]
  assign x503_sum_1_reset = reset; // @[:@32048.4]
  assign x503_sum_1_io_a = {_T_932,_T_933}; // @[Math.scala 151:17:@32049.4]
  assign x503_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@32050.4]
  assign x503_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32051.4]
  assign RetimeWrapper_44_clock = clock; // @[:@32057.4]
  assign RetimeWrapper_44_reset = reset; // @[:@32058.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32060.4]
  assign RetimeWrapper_44_io_in = ~ x499; // @[package.scala 94:16:@32059.4]
  assign RetimeWrapper_45_clock = clock; // @[:@32066.4]
  assign RetimeWrapper_45_reset = reset; // @[:@32067.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32069.4]
  assign RetimeWrapper_45_io_in = $unsigned(_T_923); // @[package.scala 94:16:@32068.4]
  assign RetimeWrapper_46_clock = clock; // @[:@32080.4]
  assign RetimeWrapper_46_reset = reset; // @[:@32081.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32083.4]
  assign RetimeWrapper_46_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32082.4]
  assign x511_sum_1_clock = clock; // @[:@32107.4]
  assign x511_sum_1_reset = reset; // @[:@32108.4]
  assign x511_sum_1_io_a = {_T_932,_T_933}; // @[Math.scala 151:17:@32109.4]
  assign x511_sum_1_io_b = RetimeWrapper_28_io_out; // @[Math.scala 152:17:@32110.4]
  assign x511_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32111.4]
  assign RetimeWrapper_47_clock = clock; // @[:@32117.4]
  assign RetimeWrapper_47_reset = reset; // @[:@32118.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32120.4]
  assign RetimeWrapper_47_io_in = ~ x509; // @[package.scala 94:16:@32119.4]
  assign RetimeWrapper_48_clock = clock; // @[:@32131.4]
  assign RetimeWrapper_48_reset = reset; // @[:@32132.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32134.4]
  assign RetimeWrapper_48_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32133.4]
  assign x518_sum_1_clock = clock; // @[:@32158.4]
  assign x518_sum_1_reset = reset; // @[:@32159.4]
  assign x518_sum_1_io_a = {_T_932,_T_933}; // @[Math.scala 151:17:@32160.4]
  assign x518_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@32161.4]
  assign x518_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32162.4]
  assign RetimeWrapper_49_clock = clock; // @[:@32168.4]
  assign RetimeWrapper_49_reset = reset; // @[:@32169.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32171.4]
  assign RetimeWrapper_49_io_in = ~ x516; // @[package.scala 94:16:@32170.4]
  assign RetimeWrapper_50_clock = clock; // @[:@32182.4]
  assign RetimeWrapper_50_reset = reset; // @[:@32183.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32185.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32184.4]
  assign RetimeWrapper_51_clock = clock; // @[:@32203.4]
  assign RetimeWrapper_51_reset = reset; // @[:@32204.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32206.4]
  assign RetimeWrapper_51_io_in = $signed(_T_722) < $signed(32'sh0); // @[package.scala 94:16:@32205.4]
  assign RetimeWrapper_52_clock = clock; // @[:@32218.4]
  assign RetimeWrapper_52_reset = reset; // @[:@32219.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32221.4]
  assign RetimeWrapper_52_io_in = {_T_334,_T_335}; // @[package.scala 94:16:@32220.4]
  assign x525_sum_1_clock = clock; // @[:@32227.4]
  assign x525_sum_1_reset = reset; // @[:@32228.4]
  assign x525_sum_1_io_a = {_T_932,_T_933}; // @[Math.scala 151:17:@32229.4]
  assign x525_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@32230.4]
  assign x525_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32231.4]
  assign RetimeWrapper_53_clock = clock; // @[:@32237.4]
  assign RetimeWrapper_53_reset = reset; // @[:@32238.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32240.4]
  assign RetimeWrapper_53_io_in = ~ x523; // @[package.scala 94:16:@32239.4]
  assign RetimeWrapper_54_clock = clock; // @[:@32251.4]
  assign RetimeWrapper_54_reset = reset; // @[:@32252.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32254.4]
  assign RetimeWrapper_54_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32253.4]
  assign x532_sum_1_clock = clock; // @[:@32278.4]
  assign x532_sum_1_reset = reset; // @[:@32279.4]
  assign x532_sum_1_io_a = {_T_932,_T_933}; // @[Math.scala 151:17:@32280.4]
  assign x532_sum_1_io_b = {_T_790,_T_791}; // @[Math.scala 152:17:@32281.4]
  assign x532_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32282.4]
  assign RetimeWrapper_55_clock = clock; // @[:@32288.4]
  assign RetimeWrapper_55_reset = reset; // @[:@32289.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32291.4]
  assign RetimeWrapper_55_io_in = ~ x530; // @[package.scala 94:16:@32290.4]
  assign RetimeWrapper_56_clock = clock; // @[:@32302.4]
  assign RetimeWrapper_56_reset = reset; // @[:@32303.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32305.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32304.4]
  assign x539_sum_1_clock = clock; // @[:@32331.4]
  assign x539_sum_1_reset = reset; // @[:@32332.4]
  assign x539_sum_1_io_a = {_T_932,_T_933}; // @[Math.scala 151:17:@32333.4]
  assign x539_sum_1_io_b = {_T_850,_T_851}; // @[Math.scala 152:17:@32334.4]
  assign x539_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32335.4]
  assign RetimeWrapper_57_clock = clock; // @[:@32341.4]
  assign RetimeWrapper_57_reset = reset; // @[:@32342.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32344.4]
  assign RetimeWrapper_57_io_in = ~ x537; // @[package.scala 94:16:@32343.4]
  assign RetimeWrapper_58_clock = clock; // @[:@32355.4]
  assign RetimeWrapper_58_reset = reset; // @[:@32356.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32358.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32357.4]
  assign x544_rdrow_1_clock = clock; // @[:@32378.4]
  assign x544_rdrow_1_reset = reset; // @[:@32379.4]
  assign x544_rdrow_1_io_a = RetimeWrapper_17_io_out; // @[Math.scala 192:17:@32380.4]
  assign x544_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@32381.4]
  assign x544_rdrow_1_io_flow = io_in_x374_TREADY; // @[Math.scala 194:20:@32382.4]
  assign x551_sum_1_clock = clock; // @[:@32432.4]
  assign x551_sum_1_reset = reset; // @[:@32433.4]
  assign x551_sum_1_io_a = {_T_1190,_T_1191}; // @[Math.scala 151:17:@32434.4]
  assign x551_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@32435.4]
  assign x551_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32436.4]
  assign RetimeWrapper_59_clock = clock; // @[:@32442.4]
  assign RetimeWrapper_59_reset = reset; // @[:@32443.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32445.4]
  assign RetimeWrapper_59_io_in = $unsigned(_T_1181); // @[package.scala 94:16:@32444.4]
  assign RetimeWrapper_60_clock = clock; // @[:@32451.4]
  assign RetimeWrapper_60_reset = reset; // @[:@32452.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32454.4]
  assign RetimeWrapper_60_io_in = ~ x547; // @[package.scala 94:16:@32453.4]
  assign RetimeWrapper_61_clock = clock; // @[:@32465.4]
  assign RetimeWrapper_61_reset = reset; // @[:@32466.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32468.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32467.4]
  assign x559_sum_1_clock = clock; // @[:@32492.4]
  assign x559_sum_1_reset = reset; // @[:@32493.4]
  assign x559_sum_1_io_a = {_T_1190,_T_1191}; // @[Math.scala 151:17:@32494.4]
  assign x559_sum_1_io_b = RetimeWrapper_28_io_out; // @[Math.scala 152:17:@32495.4]
  assign x559_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32496.4]
  assign RetimeWrapper_62_clock = clock; // @[:@32502.4]
  assign RetimeWrapper_62_reset = reset; // @[:@32503.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32505.4]
  assign RetimeWrapper_62_io_in = ~ x557; // @[package.scala 94:16:@32504.4]
  assign RetimeWrapper_63_clock = clock; // @[:@32516.4]
  assign RetimeWrapper_63_reset = reset; // @[:@32517.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32519.4]
  assign RetimeWrapper_63_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32518.4]
  assign x566_sum_1_clock = clock; // @[:@32543.4]
  assign x566_sum_1_reset = reset; // @[:@32544.4]
  assign x566_sum_1_io_a = {_T_1190,_T_1191}; // @[Math.scala 151:17:@32545.4]
  assign x566_sum_1_io_b = RetimeWrapper_32_io_out; // @[Math.scala 152:17:@32546.4]
  assign x566_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32547.4]
  assign RetimeWrapper_64_clock = clock; // @[:@32553.4]
  assign RetimeWrapper_64_reset = reset; // @[:@32554.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32556.4]
  assign RetimeWrapper_64_io_in = ~ x564; // @[package.scala 94:16:@32555.4]
  assign RetimeWrapper_65_clock = clock; // @[:@32567.4]
  assign RetimeWrapper_65_reset = reset; // @[:@32568.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32570.4]
  assign RetimeWrapper_65_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32569.4]
  assign x573_sum_1_clock = clock; // @[:@32594.4]
  assign x573_sum_1_reset = reset; // @[:@32595.4]
  assign x573_sum_1_io_a = {_T_1190,_T_1191}; // @[Math.scala 151:17:@32596.4]
  assign x573_sum_1_io_b = RetimeWrapper_52_io_out; // @[Math.scala 152:17:@32597.4]
  assign x573_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32598.4]
  assign RetimeWrapper_66_clock = clock; // @[:@32604.4]
  assign RetimeWrapper_66_reset = reset; // @[:@32605.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32607.4]
  assign RetimeWrapper_66_io_in = ~ x571; // @[package.scala 94:16:@32606.4]
  assign RetimeWrapper_67_clock = clock; // @[:@32618.4]
  assign RetimeWrapper_67_reset = reset; // @[:@32619.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32621.4]
  assign RetimeWrapper_67_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32620.4]
  assign x580_sum_1_clock = clock; // @[:@32645.4]
  assign x580_sum_1_reset = reset; // @[:@32646.4]
  assign x580_sum_1_io_a = {_T_1190,_T_1191}; // @[Math.scala 151:17:@32647.4]
  assign x580_sum_1_io_b = {_T_790,_T_791}; // @[Math.scala 152:17:@32648.4]
  assign x580_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32649.4]
  assign RetimeWrapper_68_clock = clock; // @[:@32655.4]
  assign RetimeWrapper_68_reset = reset; // @[:@32656.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32658.4]
  assign RetimeWrapper_68_io_in = ~ x578; // @[package.scala 94:16:@32657.4]
  assign RetimeWrapper_69_clock = clock; // @[:@32669.4]
  assign RetimeWrapper_69_reset = reset; // @[:@32670.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32672.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32671.4]
  assign x587_sum_1_clock = clock; // @[:@32696.4]
  assign x587_sum_1_reset = reset; // @[:@32697.4]
  assign x587_sum_1_io_a = {_T_1190,_T_1191}; // @[Math.scala 151:17:@32698.4]
  assign x587_sum_1_io_b = {_T_850,_T_851}; // @[Math.scala 152:17:@32699.4]
  assign x587_sum_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32700.4]
  assign RetimeWrapper_70_clock = clock; // @[:@32706.4]
  assign RetimeWrapper_70_reset = reset; // @[:@32707.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32709.4]
  assign RetimeWrapper_70_io_in = ~ x585; // @[package.scala 94:16:@32708.4]
  assign RetimeWrapper_71_clock = clock; // @[:@32720.4]
  assign RetimeWrapper_71_reset = reset; // @[:@32721.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32723.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32722.4]
  assign x597_x23_1_clock = clock; // @[:@32768.4]
  assign x597_x23_1_reset = reset; // @[:@32769.4]
  assign x597_x23_1_io_a = x386_lb_0_io_rPort_14_output_0; // @[Math.scala 151:17:@32770.4]
  assign x597_x23_1_io_b = _T_1395[7:0]; // @[Math.scala 152:17:@32771.4]
  assign x597_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32772.4]
  assign x598_x24_1_clock = clock; // @[:@32778.4]
  assign x598_x24_1_reset = reset; // @[:@32779.4]
  assign x598_x24_1_io_a = x386_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@32780.4]
  assign x598_x24_1_io_b = _T_1399[7:0]; // @[Math.scala 152:17:@32781.4]
  assign x598_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32782.4]
  assign x599_x23_1_clock = clock; // @[:@32788.4]
  assign x599_x23_1_reset = reset; // @[:@32789.4]
  assign x599_x23_1_io_a = _T_1403[7:0]; // @[Math.scala 151:17:@32790.4]
  assign x599_x23_1_io_b = _T_1407[7:0]; // @[Math.scala 152:17:@32791.4]
  assign x599_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32792.4]
  assign x600_x24_1_clock = clock; // @[:@32798.4]
  assign x600_x24_1_reset = reset; // @[:@32799.4]
  assign x600_x24_1_io_a = x386_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@32800.4]
  assign x600_x24_1_io_b = _T_1411[7:0]; // @[Math.scala 152:17:@32801.4]
  assign x600_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32802.4]
  assign x601_x23_1_io_a = x597_x23_1_io_result; // @[Math.scala 151:17:@32810.4]
  assign x601_x23_1_io_b = x598_x24_1_io_result; // @[Math.scala 152:17:@32811.4]
  assign x602_x24_1_io_a = x599_x23_1_io_result; // @[Math.scala 151:17:@32820.4]
  assign x602_x24_1_io_b = x600_x24_1_io_result; // @[Math.scala 152:17:@32821.4]
  assign x603_x23_1_io_a = x601_x23_1_io_result; // @[Math.scala 151:17:@32830.4]
  assign x603_x23_1_io_b = x602_x24_1_io_result; // @[Math.scala 152:17:@32831.4]
  assign RetimeWrapper_72_clock = clock; // @[:@32838.4]
  assign RetimeWrapper_72_reset = reset; // @[:@32839.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32841.4]
  assign RetimeWrapper_72_io_in = x386_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@32840.4]
  assign x604_sum_1_io_a = x603_x23_1_io_result; // @[Math.scala 151:17:@32849.4]
  assign x604_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@32850.4]
  assign RetimeWrapper_73_clock = clock; // @[:@32861.4]
  assign RetimeWrapper_73_reset = reset; // @[:@32862.4]
  assign RetimeWrapper_73_io_flow = io_in_x374_TREADY; // @[package.scala 95:18:@32864.4]
  assign RetimeWrapper_73_io_in = {4'h0,_T_1447}; // @[package.scala 94:16:@32863.4]
  assign x611_x23_1_clock = clock; // @[:@32896.4]
  assign x611_x23_1_reset = reset; // @[:@32897.4]
  assign x611_x23_1_io_a = x386_lb_0_io_rPort_17_output_0; // @[Math.scala 151:17:@32898.4]
  assign x611_x23_1_io_b = _T_1454[7:0]; // @[Math.scala 152:17:@32899.4]
  assign x611_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32900.4]
  assign x612_x24_1_clock = clock; // @[:@32906.4]
  assign x612_x24_1_reset = reset; // @[:@32907.4]
  assign x612_x24_1_io_a = x386_lb_0_io_rPort_12_output_0; // @[Math.scala 151:17:@32908.4]
  assign x612_x24_1_io_b = _T_1458[7:0]; // @[Math.scala 152:17:@32909.4]
  assign x612_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32910.4]
  assign x613_x23_1_clock = clock; // @[:@32916.4]
  assign x613_x23_1_reset = reset; // @[:@32917.4]
  assign x613_x23_1_io_a = _T_1462[7:0]; // @[Math.scala 151:17:@32918.4]
  assign x613_x23_1_io_b = _T_1466[7:0]; // @[Math.scala 152:17:@32919.4]
  assign x613_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32920.4]
  assign x614_x24_1_clock = clock; // @[:@32926.4]
  assign x614_x24_1_reset = reset; // @[:@32927.4]
  assign x614_x24_1_io_a = x386_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@32928.4]
  assign x614_x24_1_io_b = _T_1470[7:0]; // @[Math.scala 152:17:@32929.4]
  assign x614_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@32930.4]
  assign x615_x23_1_io_a = x611_x23_1_io_result; // @[Math.scala 151:17:@32938.4]
  assign x615_x23_1_io_b = x612_x24_1_io_result; // @[Math.scala 152:17:@32939.4]
  assign x616_x24_1_io_a = x613_x23_1_io_result; // @[Math.scala 151:17:@32948.4]
  assign x616_x24_1_io_b = x614_x24_1_io_result; // @[Math.scala 152:17:@32949.4]
  assign x617_x23_1_io_a = x615_x23_1_io_result; // @[Math.scala 151:17:@32958.4]
  assign x617_x23_1_io_b = x616_x24_1_io_result; // @[Math.scala 152:17:@32959.4]
  assign RetimeWrapper_74_clock = clock; // @[:@32966.4]
  assign RetimeWrapper_74_reset = reset; // @[:@32967.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32969.4]
  assign RetimeWrapper_74_io_in = x386_lb_0_io_rPort_13_output_0; // @[package.scala 94:16:@32968.4]
  assign x618_sum_1_io_a = x617_x23_1_io_result; // @[Math.scala 151:17:@32977.4]
  assign x618_sum_1_io_b = RetimeWrapper_74_io_out; // @[Math.scala 152:17:@32978.4]
  assign RetimeWrapper_75_clock = clock; // @[:@32989.4]
  assign RetimeWrapper_75_reset = reset; // @[:@32990.4]
  assign RetimeWrapper_75_io_flow = io_in_x374_TREADY; // @[package.scala 95:18:@32992.4]
  assign RetimeWrapper_75_io_in = {4'h0,_T_1506}; // @[package.scala 94:16:@32991.4]
  assign x624_x23_1_clock = clock; // @[:@33019.4]
  assign x624_x23_1_reset = reset; // @[:@33020.4]
  assign x624_x23_1_io_a = x386_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@33021.4]
  assign x624_x23_1_io_b = _T_1513[7:0]; // @[Math.scala 152:17:@33022.4]
  assign x624_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33023.4]
  assign x625_x24_1_clock = clock; // @[:@33029.4]
  assign x625_x24_1_reset = reset; // @[:@33030.4]
  assign x625_x24_1_io_a = x386_lb_0_io_rPort_15_output_0; // @[Math.scala 151:17:@33031.4]
  assign x625_x24_1_io_b = _T_1407[7:0]; // @[Math.scala 152:17:@33032.4]
  assign x625_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33033.4]
  assign x626_x23_1_clock = clock; // @[:@33039.4]
  assign x626_x23_1_reset = reset; // @[:@33040.4]
  assign x626_x23_1_io_a = _T_1517[7:0]; // @[Math.scala 151:17:@33041.4]
  assign x626_x23_1_io_b = _T_1521[7:0]; // @[Math.scala 152:17:@33042.4]
  assign x626_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33043.4]
  assign x627_x24_1_clock = clock; // @[:@33049.4]
  assign x627_x24_1_reset = reset; // @[:@33050.4]
  assign x627_x24_1_io_a = x386_lb_0_io_rPort_6_output_0; // @[Math.scala 151:17:@33051.4]
  assign x627_x24_1_io_b = _T_1525[7:0]; // @[Math.scala 152:17:@33052.4]
  assign x627_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33053.4]
  assign x628_x23_1_io_a = x624_x23_1_io_result; // @[Math.scala 151:17:@33061.4]
  assign x628_x23_1_io_b = x625_x24_1_io_result; // @[Math.scala 152:17:@33062.4]
  assign x629_x24_1_io_a = x626_x23_1_io_result; // @[Math.scala 151:17:@33071.4]
  assign x629_x24_1_io_b = x627_x24_1_io_result; // @[Math.scala 152:17:@33072.4]
  assign x630_x23_1_io_a = x628_x23_1_io_result; // @[Math.scala 151:17:@33081.4]
  assign x630_x23_1_io_b = x629_x24_1_io_result; // @[Math.scala 152:17:@33082.4]
  assign RetimeWrapper_76_clock = clock; // @[:@33089.4]
  assign RetimeWrapper_76_reset = reset; // @[:@33090.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33092.4]
  assign RetimeWrapper_76_io_in = x386_lb_0_io_rPort_4_output_0; // @[package.scala 94:16:@33091.4]
  assign x631_sum_1_io_a = x630_x23_1_io_result; // @[Math.scala 151:17:@33100.4]
  assign x631_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@33101.4]
  assign RetimeWrapper_77_clock = clock; // @[:@33112.4]
  assign RetimeWrapper_77_reset = reset; // @[:@33113.4]
  assign RetimeWrapper_77_io_flow = io_in_x374_TREADY; // @[package.scala 95:18:@33115.4]
  assign RetimeWrapper_77_io_in = {4'h0,_T_1561}; // @[package.scala 94:16:@33114.4]
  assign x637_x23_1_clock = clock; // @[:@33142.4]
  assign x637_x23_1_reset = reset; // @[:@33143.4]
  assign x637_x23_1_io_a = x386_lb_0_io_rPort_12_output_0; // @[Math.scala 151:17:@33144.4]
  assign x637_x23_1_io_b = _T_1568[7:0]; // @[Math.scala 152:17:@33145.4]
  assign x637_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33146.4]
  assign x638_x24_1_clock = clock; // @[:@33154.4]
  assign x638_x24_1_reset = reset; // @[:@33155.4]
  assign x638_x24_1_io_a = x386_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@33156.4]
  assign x638_x24_1_io_b = _T_1466[7:0]; // @[Math.scala 152:17:@33157.4]
  assign x638_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33158.4]
  assign x639_x23_1_clock = clock; // @[:@33164.4]
  assign x639_x23_1_reset = reset; // @[:@33165.4]
  assign x639_x23_1_io_a = _T_1572[7:0]; // @[Math.scala 151:17:@33166.4]
  assign x639_x23_1_io_b = _T_1576[7:0]; // @[Math.scala 152:17:@33167.4]
  assign x639_x23_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33168.4]
  assign x640_x24_1_clock = clock; // @[:@33174.4]
  assign x640_x24_1_reset = reset; // @[:@33175.4]
  assign x640_x24_1_io_a = x386_lb_0_io_rPort_13_output_0; // @[Math.scala 151:17:@33176.4]
  assign x640_x24_1_io_b = _T_1580[7:0]; // @[Math.scala 152:17:@33177.4]
  assign x640_x24_1_io_flow = io_in_x374_TREADY; // @[Math.scala 153:20:@33178.4]
  assign x641_x23_1_io_a = x637_x23_1_io_result; // @[Math.scala 151:17:@33186.4]
  assign x641_x23_1_io_b = x638_x24_1_io_result; // @[Math.scala 152:17:@33187.4]
  assign x642_x24_1_io_a = x639_x23_1_io_result; // @[Math.scala 151:17:@33196.4]
  assign x642_x24_1_io_b = x640_x24_1_io_result; // @[Math.scala 152:17:@33197.4]
  assign x643_x23_1_io_a = x641_x23_1_io_result; // @[Math.scala 151:17:@33206.4]
  assign x643_x23_1_io_b = x642_x24_1_io_result; // @[Math.scala 152:17:@33207.4]
  assign RetimeWrapper_78_clock = clock; // @[:@33214.4]
  assign RetimeWrapper_78_reset = reset; // @[:@33215.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33217.4]
  assign RetimeWrapper_78_io_in = x386_lb_0_io_rPort_5_output_0; // @[package.scala 94:16:@33216.4]
  assign x644_sum_1_io_a = x643_x23_1_io_result; // @[Math.scala 151:17:@33225.4]
  assign x644_sum_1_io_b = RetimeWrapper_78_io_out; // @[Math.scala 152:17:@33226.4]
  assign RetimeWrapper_79_clock = clock; // @[:@33237.4]
  assign RetimeWrapper_79_reset = reset; // @[:@33238.4]
  assign RetimeWrapper_79_io_flow = io_in_x374_TREADY; // @[package.scala 95:18:@33240.4]
  assign RetimeWrapper_79_io_in = {4'h0,_T_1618}; // @[package.scala 94:16:@33239.4]
  assign RetimeWrapper_80_clock = clock; // @[:@33247.4]
  assign RetimeWrapper_80_reset = reset; // @[:@33248.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33250.4]
  assign RetimeWrapper_80_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33249.4]
  assign RetimeWrapper_81_clock = clock; // @[:@33256.4]
  assign RetimeWrapper_81_reset = reset; // @[:@33257.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33259.4]
  assign RetimeWrapper_81_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33258.4]
  assign RetimeWrapper_82_clock = clock; // @[:@33265.4]
  assign RetimeWrapper_82_reset = reset; // @[:@33266.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33268.4]
  assign RetimeWrapper_82_io_in = $unsigned(_T_315); // @[package.scala 94:16:@33267.4]
  assign RetimeWrapper_83_clock = clock; // @[:@33274.4]
  assign RetimeWrapper_83_reset = reset; // @[:@33275.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33277.4]
  assign RetimeWrapper_83_io_in = x401_sum_1_io_result; // @[package.scala 94:16:@33276.4]
  assign RetimeWrapper_84_clock = clock; // @[:@33287.4]
  assign RetimeWrapper_84_reset = reset; // @[:@33288.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33290.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33289.4]
  assign RetimeWrapper_85_clock = clock; // @[:@33308.4]
  assign RetimeWrapper_85_reset = reset; // @[:@33309.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33311.4]
  assign RetimeWrapper_85_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@33310.4]
  assign RetimeWrapper_86_clock = clock; // @[:@33321.4]
  assign RetimeWrapper_86_reset = reset; // @[:@33322.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33324.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33323.4]
  assign RetimeWrapper_87_clock = clock; // @[:@33342.4]
  assign RetimeWrapper_87_reset = reset; // @[:@33343.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33345.4]
  assign RetimeWrapper_87_io_in = x420_sum_1_io_result; // @[package.scala 94:16:@33344.4]
  assign RetimeWrapper_88_clock = clock; // @[:@33355.4]
  assign RetimeWrapper_88_reset = reset; // @[:@33356.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33358.4]
  assign RetimeWrapper_88_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33357.4]
  assign RetimeWrapper_89_clock = clock; // @[:@33376.4]
  assign RetimeWrapper_89_reset = reset; // @[:@33377.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33379.4]
  assign RetimeWrapper_89_io_in = x429_sum_1_io_result; // @[package.scala 94:16:@33378.4]
  assign RetimeWrapper_90_clock = clock; // @[:@33389.4]
  assign RetimeWrapper_90_reset = reset; // @[:@33390.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33392.4]
  assign RetimeWrapper_90_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33391.4]
  assign RetimeWrapper_91_clock = clock; // @[:@33410.4]
  assign RetimeWrapper_91_reset = reset; // @[:@33411.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33413.4]
  assign RetimeWrapper_91_io_in = $unsigned(_T_564); // @[package.scala 94:16:@33412.4]
  assign RetimeWrapper_92_clock = clock; // @[:@33419.4]
  assign RetimeWrapper_92_reset = reset; // @[:@33420.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33422.4]
  assign RetimeWrapper_92_io_in = ~ x438; // @[package.scala 94:16:@33421.4]
  assign RetimeWrapper_93_clock = clock; // @[:@33428.4]
  assign RetimeWrapper_93_reset = reset; // @[:@33429.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33431.4]
  assign RetimeWrapper_93_io_in = x442_sum_1_io_result; // @[package.scala 94:16:@33430.4]
  assign RetimeWrapper_94_clock = clock; // @[:@33442.4]
  assign RetimeWrapper_94_reset = reset; // @[:@33443.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33445.4]
  assign RetimeWrapper_94_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33444.4]
  assign RetimeWrapper_95_clock = clock; // @[:@33463.4]
  assign RetimeWrapper_95_reset = reset; // @[:@33464.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33466.4]
  assign RetimeWrapper_95_io_in = x451_sum_1_io_result; // @[package.scala 94:16:@33465.4]
  assign RetimeWrapper_96_clock = clock; // @[:@33472.4]
  assign RetimeWrapper_96_reset = reset; // @[:@33473.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33475.4]
  assign RetimeWrapper_96_io_in = ~ x449; // @[package.scala 94:16:@33474.4]
  assign RetimeWrapper_97_clock = clock; // @[:@33486.4]
  assign RetimeWrapper_97_reset = reset; // @[:@33487.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33489.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33488.4]
  assign RetimeWrapper_98_clock = clock; // @[:@33507.4]
  assign RetimeWrapper_98_reset = reset; // @[:@33508.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33510.4]
  assign RetimeWrapper_98_io_in = ~ x457; // @[package.scala 94:16:@33509.4]
  assign RetimeWrapper_99_clock = clock; // @[:@33516.4]
  assign RetimeWrapper_99_reset = reset; // @[:@33517.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33519.4]
  assign RetimeWrapper_99_io_in = x459_sum_1_io_result; // @[package.scala 94:16:@33518.4]
  assign RetimeWrapper_100_clock = clock; // @[:@33530.4]
  assign RetimeWrapper_100_reset = reset; // @[:@33531.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33533.4]
  assign RetimeWrapper_100_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33532.4]
  assign RetimeWrapper_101_clock = clock; // @[:@33551.4]
  assign RetimeWrapper_101_reset = reset; // @[:@33552.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33554.4]
  assign RetimeWrapper_101_io_in = x467_sum_1_io_result; // @[package.scala 94:16:@33553.4]
  assign RetimeWrapper_102_clock = clock; // @[:@33560.4]
  assign RetimeWrapper_102_reset = reset; // @[:@33561.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33563.4]
  assign RetimeWrapper_102_io_in = ~ x465; // @[package.scala 94:16:@33562.4]
  assign RetimeWrapper_103_clock = clock; // @[:@33574.4]
  assign RetimeWrapper_103_reset = reset; // @[:@33575.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33577.4]
  assign RetimeWrapper_103_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33576.4]
  assign RetimeWrapper_104_clock = clock; // @[:@33595.4]
  assign RetimeWrapper_104_reset = reset; // @[:@33596.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33598.4]
  assign RetimeWrapper_104_io_in = ~ x474; // @[package.scala 94:16:@33597.4]
  assign RetimeWrapper_105_clock = clock; // @[:@33604.4]
  assign RetimeWrapper_105_reset = reset; // @[:@33605.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33607.4]
  assign RetimeWrapper_105_io_in = x478_sum_1_io_result; // @[package.scala 94:16:@33606.4]
  assign RetimeWrapper_106_clock = clock; // @[:@33618.4]
  assign RetimeWrapper_106_reset = reset; // @[:@33619.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33621.4]
  assign RetimeWrapper_106_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33620.4]
  assign RetimeWrapper_107_clock = clock; // @[:@33639.4]
  assign RetimeWrapper_107_reset = reset; // @[:@33640.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33642.4]
  assign RetimeWrapper_107_io_in = ~ x499; // @[package.scala 94:16:@33641.4]
  assign RetimeWrapper_108_clock = clock; // @[:@33648.4]
  assign RetimeWrapper_108_reset = reset; // @[:@33649.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33651.4]
  assign RetimeWrapper_108_io_in = x503_sum_1_io_result; // @[package.scala 94:16:@33650.4]
  assign RetimeWrapper_109_clock = clock; // @[:@33657.4]
  assign RetimeWrapper_109_reset = reset; // @[:@33658.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33660.4]
  assign RetimeWrapper_109_io_in = $unsigned(_T_923); // @[package.scala 94:16:@33659.4]
  assign RetimeWrapper_110_clock = clock; // @[:@33671.4]
  assign RetimeWrapper_110_reset = reset; // @[:@33672.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33674.4]
  assign RetimeWrapper_110_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33673.4]
  assign RetimeWrapper_111_clock = clock; // @[:@33692.4]
  assign RetimeWrapper_111_reset = reset; // @[:@33693.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33695.4]
  assign RetimeWrapper_111_io_in = x511_sum_1_io_result; // @[package.scala 94:16:@33694.4]
  assign RetimeWrapper_112_clock = clock; // @[:@33701.4]
  assign RetimeWrapper_112_reset = reset; // @[:@33702.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33704.4]
  assign RetimeWrapper_112_io_in = ~ x509; // @[package.scala 94:16:@33703.4]
  assign RetimeWrapper_113_clock = clock; // @[:@33715.4]
  assign RetimeWrapper_113_reset = reset; // @[:@33716.4]
  assign RetimeWrapper_113_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33718.4]
  assign RetimeWrapper_113_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33717.4]
  assign RetimeWrapper_114_clock = clock; // @[:@33736.4]
  assign RetimeWrapper_114_reset = reset; // @[:@33737.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33739.4]
  assign RetimeWrapper_114_io_in = x518_sum_1_io_result; // @[package.scala 94:16:@33738.4]
  assign RetimeWrapper_115_clock = clock; // @[:@33745.4]
  assign RetimeWrapper_115_reset = reset; // @[:@33746.4]
  assign RetimeWrapper_115_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33748.4]
  assign RetimeWrapper_115_io_in = ~ x516; // @[package.scala 94:16:@33747.4]
  assign RetimeWrapper_116_clock = clock; // @[:@33759.4]
  assign RetimeWrapper_116_reset = reset; // @[:@33760.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33762.4]
  assign RetimeWrapper_116_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33761.4]
  assign RetimeWrapper_117_clock = clock; // @[:@33780.4]
  assign RetimeWrapper_117_reset = reset; // @[:@33781.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33783.4]
  assign RetimeWrapper_117_io_in = x525_sum_1_io_result; // @[package.scala 94:16:@33782.4]
  assign RetimeWrapper_118_clock = clock; // @[:@33789.4]
  assign RetimeWrapper_118_reset = reset; // @[:@33790.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33792.4]
  assign RetimeWrapper_118_io_in = ~ x523; // @[package.scala 94:16:@33791.4]
  assign RetimeWrapper_119_clock = clock; // @[:@33803.4]
  assign RetimeWrapper_119_reset = reset; // @[:@33804.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33806.4]
  assign RetimeWrapper_119_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33805.4]
  assign RetimeWrapper_120_clock = clock; // @[:@33824.4]
  assign RetimeWrapper_120_reset = reset; // @[:@33825.4]
  assign RetimeWrapper_120_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33827.4]
  assign RetimeWrapper_120_io_in = ~ x530; // @[package.scala 94:16:@33826.4]
  assign RetimeWrapper_121_clock = clock; // @[:@33833.4]
  assign RetimeWrapper_121_reset = reset; // @[:@33834.4]
  assign RetimeWrapper_121_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33836.4]
  assign RetimeWrapper_121_io_in = x532_sum_1_io_result; // @[package.scala 94:16:@33835.4]
  assign RetimeWrapper_122_clock = clock; // @[:@33847.4]
  assign RetimeWrapper_122_reset = reset; // @[:@33848.4]
  assign RetimeWrapper_122_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33850.4]
  assign RetimeWrapper_122_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33849.4]
  assign x674_x25_1_io_a = x387_lb2_0_io_rPort_8_output_0; // @[Math.scala 151:17:@33882.4]
  assign x674_x25_1_io_b = _T_2016[7:0]; // @[Math.scala 152:17:@33883.4]
  assign x675_x26_1_io_a = _T_2020[7:0]; // @[Math.scala 151:17:@33892.4]
  assign x675_x26_1_io_b = x387_lb2_0_io_rPort_9_output_0; // @[Math.scala 152:17:@33893.4]
  assign x676_sum_1_io_a = x674_x25_1_io_result; // @[Math.scala 151:17:@33902.4]
  assign x676_sum_1_io_b = x675_x26_1_io_result; // @[Math.scala 152:17:@33903.4]
  assign x677_div_1_clock = clock; // @[:@33912.4]
  assign x677_div_1_reset = reset; // @[:@33913.4]
  assign x677_div_1_io_a = x676_sum_1_io_result; // @[Math.scala 328:17:@33914.4]
  assign x677_div_1_io_flow = io_in_x374_TREADY; // @[Math.scala 330:20:@33916.4]
  assign x680_x25_1_io_a = x387_lb2_0_io_rPort_3_output_0; // @[Math.scala 151:17:@33934.4]
  assign x680_x25_1_io_b = _T_2040[7:0]; // @[Math.scala 152:17:@33935.4]
  assign x681_x26_1_io_a = _T_2044[7:0]; // @[Math.scala 151:17:@33944.4]
  assign x681_x26_1_io_b = x387_lb2_0_io_rPort_0_output_0; // @[Math.scala 152:17:@33945.4]
  assign x682_sum_1_io_a = x680_x25_1_io_result; // @[Math.scala 151:17:@33954.4]
  assign x682_sum_1_io_b = x681_x26_1_io_result; // @[Math.scala 152:17:@33955.4]
  assign x683_div_1_clock = clock; // @[:@33964.4]
  assign x683_div_1_reset = reset; // @[:@33965.4]
  assign x683_div_1_io_a = x682_sum_1_io_result; // @[Math.scala 328:17:@33966.4]
  assign x683_div_1_io_flow = io_in_x374_TREADY; // @[Math.scala 330:20:@33968.4]
  assign x686_x25_1_io_a = x387_lb2_0_io_rPort_7_output_0; // @[Math.scala 151:17:@33986.4]
  assign x686_x25_1_io_b = _T_2064[7:0]; // @[Math.scala 152:17:@33987.4]
  assign x687_x26_1_io_a = _T_2068[7:0]; // @[Math.scala 151:17:@33996.4]
  assign x687_x26_1_io_b = x387_lb2_0_io_rPort_5_output_0; // @[Math.scala 152:17:@33997.4]
  assign x688_sum_1_io_a = x686_x25_1_io_result; // @[Math.scala 151:17:@34006.4]
  assign x688_sum_1_io_b = x687_x26_1_io_result; // @[Math.scala 152:17:@34007.4]
  assign x689_div_1_clock = clock; // @[:@34016.4]
  assign x689_div_1_reset = reset; // @[:@34017.4]
  assign x689_div_1_io_a = x688_sum_1_io_result; // @[Math.scala 328:17:@34018.4]
  assign x689_div_1_io_flow = io_in_x374_TREADY; // @[Math.scala 330:20:@34020.4]
  assign x692_x25_1_io_a = x387_lb2_0_io_rPort_6_output_0; // @[Math.scala 151:17:@34038.4]
  assign x692_x25_1_io_b = _T_2088[7:0]; // @[Math.scala 152:17:@34039.4]
  assign x693_x26_1_io_a = _T_2092[7:0]; // @[Math.scala 151:17:@34048.4]
  assign x693_x26_1_io_b = x387_lb2_0_io_rPort_1_output_0; // @[Math.scala 152:17:@34049.4]
  assign x694_sum_1_io_a = x692_x25_1_io_result; // @[Math.scala 151:17:@34058.4]
  assign x694_sum_1_io_b = x693_x26_1_io_result; // @[Math.scala 152:17:@34059.4]
  assign x695_div_1_clock = clock; // @[:@34068.4]
  assign x695_div_1_reset = reset; // @[:@34069.4]
  assign x695_div_1_io_a = x694_sum_1_io_result; // @[Math.scala 328:17:@34070.4]
  assign x695_div_1_io_flow = io_in_x374_TREADY; // @[Math.scala 330:20:@34072.4]
  assign RetimeWrapper_123_clock = clock; // @[:@34088.4]
  assign RetimeWrapper_123_reset = reset; // @[:@34089.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34091.4]
  assign RetimeWrapper_123_io_in = {_T_2121,_T_2120}; // @[package.scala 94:16:@34090.4]
  assign RetimeWrapper_124_clock = clock; // @[:@34097.4]
  assign RetimeWrapper_124_reset = reset; // @[:@34098.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34100.4]
  assign RetimeWrapper_124_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@34099.4]
  assign RetimeWrapper_125_clock = clock; // @[:@34106.4]
  assign RetimeWrapper_125_reset = reset; // @[:@34107.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34109.4]
  assign RetimeWrapper_125_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@34108.4]
  assign RetimeWrapper_126_clock = clock; // @[:@34115.4]
  assign RetimeWrapper_126_reset = reset; // @[:@34116.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34118.4]
  assign RetimeWrapper_126_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34117.4]
endmodule
module x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1( // @[:@34136.2]
  input          clock, // @[:@34137.4]
  input          reset, // @[:@34138.4]
  output         io_in_x374_TVALID, // @[:@34139.4]
  input          io_in_x374_TREADY, // @[:@34139.4]
  output [255:0] io_in_x374_TDATA, // @[:@34139.4]
  input          io_in_x373_TVALID, // @[:@34139.4]
  output         io_in_x373_TREADY, // @[:@34139.4]
  input  [255:0] io_in_x373_TDATA, // @[:@34139.4]
  input  [7:0]   io_in_x373_TID, // @[:@34139.4]
  input  [7:0]   io_in_x373_TDEST, // @[:@34139.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@34139.4]
  input          io_sigsIn_smChildAcks_0, // @[:@34139.4]
  output         io_sigsOut_smDoneIn_0, // @[:@34139.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@34139.4]
  input          io_rr // @[:@34139.4]
);
  wire  x381_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x381_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x381_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x381_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire [31:0] x381_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire [31:0] x381_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x381_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x381_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x381_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@34149.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34236.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34236.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34236.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34236.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34236.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@34286.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@34286.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@34286.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@34286.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@34286.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TVALID; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TREADY; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire [255:0] x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TDATA; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TREADY; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire [255:0] x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TDATA; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire [7:0] x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TID; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire [7:0] x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TDEST; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire [31:0] x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire [31:0] x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
  wire  _T_239; // @[package.scala 96:25:@34241.4 package.scala 96:25:@34242.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x701_outr_UnitPipe.scala 68:66:@34247.4]
  wire  _T_252; // @[package.scala 96:25:@34283.4 package.scala 96:25:@34284.4]
  wire  _T_258; // @[package.scala 96:25:@34291.4 package.scala 96:25:@34292.4]
  wire  _T_261; // @[SpatialBlocks.scala 110:93:@34294.4]
  wire  x700_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 110:90:@34295.4]
  wire  _T_263; // @[SpatialBlocks.scala 128:36:@34303.4]
  wire  _T_264; // @[SpatialBlocks.scala 128:78:@34304.4]
  wire  _T_269; // @[SpatialBlocks.scala 130:61:@34313.4]
  x381_ctrchain x381_ctrchain ( // @[SpatialBlocks.scala 37:22:@34149.4]
    .clock(x381_ctrchain_clock),
    .reset(x381_ctrchain_reset),
    .io_input_reset(x381_ctrchain_io_input_reset),
    .io_input_enable(x381_ctrchain_io_input_enable),
    .io_output_counts_1(x381_ctrchain_io_output_counts_1),
    .io_output_counts_0(x381_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x381_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x381_ctrchain_io_output_oobs_1),
    .io_output_done(x381_ctrchain_io_output_done)
  );
  x700_inr_Foreach_SAMPLER_BOX_sm x700_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 32:18:@34208.4]
    .clock(x700_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x700_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x700_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x700_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x700_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x700_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x700_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x700_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x700_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34236.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34278.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@34286.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1 x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 909:24:@34318.4]
    .clock(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x374_TVALID(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TVALID),
    .io_in_x374_TREADY(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TREADY),
    .io_in_x374_TDATA(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TDATA),
    .io_in_x373_TREADY(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TREADY),
    .io_in_x373_TDATA(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TDATA),
    .io_in_x373_TID(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TID),
    .io_in_x373_TDEST(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TDEST),
    .io_sigsIn_backpressure(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_239 = RetimeWrapper_io_out; // @[package.scala 96:25:@34241.4 package.scala 96:25:@34242.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x373_TVALID | x700_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x701_outr_UnitPipe.scala 68:66:@34247.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34283.4 package.scala 96:25:@34284.4]
  assign _T_258 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@34291.4 package.scala 96:25:@34292.4]
  assign _T_261 = ~ _T_258; // @[SpatialBlocks.scala 110:93:@34294.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_252 & _T_261; // @[SpatialBlocks.scala 110:90:@34295.4]
  assign _T_263 = x700_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 128:36:@34303.4]
  assign _T_264 = ~ x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 128:78:@34304.4]
  assign _T_269 = x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 130:61:@34313.4]
  assign io_in_x374_TVALID = x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TVALID; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 48:23:@34376.4]
  assign io_in_x374_TDATA = x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TDATA; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 48:23:@34374.4]
  assign io_in_x373_TREADY = x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TREADY; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 49:23:@34384.4]
  assign io_sigsOut_smDoneIn_0 = x700_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 127:53:@34301.4]
  assign io_sigsOut_smCtrCopyDone_0 = x700_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 139:125:@34317.4]
  assign x381_ctrchain_clock = clock; // @[:@34150.4]
  assign x381_ctrchain_reset = reset; // @[:@34151.4]
  assign x381_ctrchain_io_input_reset = x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 130:103:@34316.4]
  assign x381_ctrchain_io_input_enable = _T_269 & x700_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 104:75:@34271.4 SpatialBlocks.scala 130:45:@34315.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@34209.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@34210.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_io_enable = x700_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x700_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 112:18:@34298.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_239 : 1'h0; // @[sm_x701_outr_UnitPipe.scala 66:50:@34244.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@34300.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x374_TREADY | x700_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 105:24:@34272.4]
  assign x700_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x701_outr_UnitPipe.scala 70:48:@34250.4]
  assign RetimeWrapper_clock = clock; // @[:@34237.4]
  assign RetimeWrapper_reset = reset; // @[:@34238.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34240.4]
  assign RetimeWrapper_io_in = x381_ctrchain_io_output_done; // @[package.scala 94:16:@34239.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34279.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34280.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34282.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@34281.4]
  assign RetimeWrapper_2_clock = clock; // @[:@34287.4]
  assign RetimeWrapper_2_reset = reset; // @[:@34288.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@34290.4]
  assign RetimeWrapper_2_io_in = x700_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@34289.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@34319.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@34320.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x374_TREADY = io_in_x374_TREADY; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 48:23:@34375.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TDATA = io_in_x373_TDATA; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 49:23:@34383.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TID = io_in_x373_TID; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 49:23:@34379.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x373_TDEST = io_in_x373_TDEST; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 49:23:@34378.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x374_TREADY | x700_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34402.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_263 & _T_264; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34400.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x700_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34398.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = x381_ctrchain_io_output_counts_1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34393.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = x381_ctrchain_io_output_counts_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34392.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x381_ctrchain_io_output_oobs_0; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34390.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x381_ctrchain_io_output_oobs_1; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 913:22:@34391.4]
  assign x700_inr_Foreach_SAMPLER_BOX_kernelx700_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x700_inr_Foreach_SAMPLER_BOX.scala 912:18:@34386.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@34415.2]
  input          clock, // @[:@34416.4]
  input          reset, // @[:@34417.4]
  output         io_in_x374_TVALID, // @[:@34418.4]
  input          io_in_x374_TREADY, // @[:@34418.4]
  output [255:0] io_in_x374_TDATA, // @[:@34418.4]
  input          io_in_x373_TVALID, // @[:@34418.4]
  output         io_in_x373_TREADY, // @[:@34418.4]
  input  [255:0] io_in_x373_TDATA, // @[:@34418.4]
  input  [7:0]   io_in_x373_TID, // @[:@34418.4]
  input  [7:0]   io_in_x373_TDEST, // @[:@34418.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@34418.4]
  input          io_sigsIn_smChildAcks_0, // @[:@34418.4]
  output         io_sigsOut_smDoneIn_0, // @[:@34418.4]
  input          io_rr // @[:@34418.4]
);
  wire  x701_outr_UnitPipe_sm_clock; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_reset; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_enable; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_done; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_parentAck; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_childAck_0; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  x701_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34611.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34611.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34611.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34611.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34611.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34619.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34619.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34619.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34619.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34619.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_clock; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_reset; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TVALID; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TREADY; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire [255:0] x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TDATA; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TVALID; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TREADY; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire [255:0] x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TDATA; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire [7:0] x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TID; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire [7:0] x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TDEST; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_rr; // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
  wire  _T_246; // @[package.scala 96:25:@34616.4 package.scala 96:25:@34617.4]
  wire  _T_252; // @[package.scala 96:25:@34624.4 package.scala 96:25:@34625.4]
  wire  _T_255; // @[SpatialBlocks.scala 110:93:@34627.4]
  x701_outr_UnitPipe_sm x701_outr_UnitPipe_sm ( // @[sm_x701_outr_UnitPipe.scala 32:18:@34559.4]
    .clock(x701_outr_UnitPipe_sm_clock),
    .reset(x701_outr_UnitPipe_sm_reset),
    .io_enable(x701_outr_UnitPipe_sm_io_enable),
    .io_done(x701_outr_UnitPipe_sm_io_done),
    .io_parentAck(x701_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x701_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x701_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x701_outr_UnitPipe_sm_io_childAck_0),
    .io_ctrCopyDone_0(x701_outr_UnitPipe_sm_io_ctrCopyDone_0)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34611.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34619.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1 x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1 ( // @[sm_x701_outr_UnitPipe.scala 75:24:@34646.4]
    .clock(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_clock),
    .reset(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_reset),
    .io_in_x374_TVALID(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TVALID),
    .io_in_x374_TREADY(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TREADY),
    .io_in_x374_TDATA(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TDATA),
    .io_in_x373_TVALID(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TVALID),
    .io_in_x373_TREADY(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TREADY),
    .io_in_x373_TDATA(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TDATA),
    .io_in_x373_TID(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TID),
    .io_in_x373_TDEST(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TDEST),
    .io_sigsIn_smEnableOuts_0(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smCtrCopyDone_0(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_rr(x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_246 = RetimeWrapper_io_out; // @[package.scala 96:25:@34616.4 package.scala 96:25:@34617.4]
  assign _T_252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34624.4 package.scala 96:25:@34625.4]
  assign _T_255 = ~ _T_252; // @[SpatialBlocks.scala 110:93:@34627.4]
  assign io_in_x374_TVALID = x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TVALID; // @[sm_x701_outr_UnitPipe.scala 48:23:@34702.4]
  assign io_in_x374_TDATA = x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TDATA; // @[sm_x701_outr_UnitPipe.scala 48:23:@34700.4]
  assign io_in_x373_TREADY = x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TREADY; // @[sm_x701_outr_UnitPipe.scala 49:23:@34710.4]
  assign io_sigsOut_smDoneIn_0 = x701_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 127:53:@34634.4]
  assign x701_outr_UnitPipe_sm_clock = clock; // @[:@34560.4]
  assign x701_outr_UnitPipe_sm_reset = reset; // @[:@34561.4]
  assign x701_outr_UnitPipe_sm_io_enable = _T_246 & _T_255; // @[SpatialBlocks.scala 112:18:@34631.4]
  assign x701_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 114:21:@34633.4]
  assign x701_outr_UnitPipe_sm_io_doneIn_0 = x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@34603.4]
  assign x701_outr_UnitPipe_sm_io_ctrCopyDone_0 = x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 132:80:@34645.4]
  assign RetimeWrapper_clock = clock; // @[:@34612.4]
  assign RetimeWrapper_reset = reset; // @[:@34613.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34615.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@34614.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34620.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34621.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34623.4]
  assign RetimeWrapper_1_io_in = x701_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@34622.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_clock = clock; // @[:@34647.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_reset = reset; // @[:@34648.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x374_TREADY = io_in_x374_TREADY; // @[sm_x701_outr_UnitPipe.scala 48:23:@34701.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TVALID = io_in_x373_TVALID; // @[sm_x701_outr_UnitPipe.scala 49:23:@34711.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TDATA = io_in_x373_TDATA; // @[sm_x701_outr_UnitPipe.scala 49:23:@34709.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TID = io_in_x373_TID; // @[sm_x701_outr_UnitPipe.scala 49:23:@34705.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_in_x373_TDEST = io_in_x373_TDEST; // @[sm_x701_outr_UnitPipe.scala 49:23:@34704.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x701_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x701_outr_UnitPipe.scala 79:22:@34720.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x701_outr_UnitPipe_sm_io_childAck_0; // @[sm_x701_outr_UnitPipe.scala 79:22:@34718.4]
  assign x701_outr_UnitPipe_kernelx701_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x701_outr_UnitPipe.scala 78:18:@34712.4]
endmodule
module AccelUnit( // @[:@34739.2]
  input          clock, // @[:@34740.4]
  input          reset, // @[:@34741.4]
  input          io_enable, // @[:@34742.4]
  output         io_done, // @[:@34742.4]
  input          io_reset, // @[:@34742.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@34742.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@34742.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@34742.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@34742.4]
  output         io_memStreams_loads_0_data_ready, // @[:@34742.4]
  input          io_memStreams_loads_0_data_valid, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@34742.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@34742.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@34742.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@34742.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@34742.4]
  input          io_memStreams_stores_0_data_ready, // @[:@34742.4]
  output         io_memStreams_stores_0_data_valid, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_1, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_2, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_3, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_4, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_5, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_6, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_7, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_8, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_9, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_10, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_11, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_12, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_13, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_14, // @[:@34742.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_15, // @[:@34742.4]
  output [15:0]  io_memStreams_stores_0_data_bits_wstrb, // @[:@34742.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@34742.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@34742.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@34742.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@34742.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@34742.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@34742.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@34742.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@34742.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@34742.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@34742.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@34742.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@34742.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@34742.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@34742.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@34742.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@34742.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@34742.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@34742.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@34742.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@34742.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@34742.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@34742.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@34742.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@34742.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@34742.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@34742.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@34742.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@34742.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@34742.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@34742.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@34742.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@34742.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@34742.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@34742.4]
  output         io_heap_0_req_valid, // @[:@34742.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@34742.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@34742.4]
  input          io_heap_0_resp_valid, // @[:@34742.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@34742.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@34742.4]
  input  [63:0]  io_argIns_0, // @[:@34742.4]
  input  [63:0]  io_argIns_1, // @[:@34742.4]
  input          io_argOuts_0_port_ready, // @[:@34742.4]
  output         io_argOuts_0_port_valid, // @[:@34742.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@34742.4]
  input  [63:0]  io_argOuts_0_echo // @[:@34742.4]
);
  wire  SingleCounter_clock; // @[Main.scala 35:32:@34905.4]
  wire  SingleCounter_reset; // @[Main.scala 35:32:@34905.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 35:32:@34905.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 35:32:@34905.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34923.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34923.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34923.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34923.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34923.4]
  wire  SRFF_clock; // @[Main.scala 39:28:@34932.4]
  wire  SRFF_reset; // @[Main.scala 39:28:@34932.4]
  wire  SRFF_io_input_set; // @[Main.scala 39:28:@34932.4]
  wire  SRFF_io_input_reset; // @[Main.scala 39:28:@34932.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 39:28:@34932.4]
  wire  SRFF_io_output; // @[Main.scala 39:28:@34932.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 32:18:@34970.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@35002.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@35002.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@35002.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@35002.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@35002.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_in_x374_TVALID; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_in_x374_TREADY; // @[sm_RootController.scala 73:24:@35061.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x374_TDATA; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_in_x373_TVALID; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_in_x373_TREADY; // @[sm_RootController.scala 73:24:@35061.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x373_TDATA; // @[sm_RootController.scala 73:24:@35061.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x373_TID; // @[sm_RootController.scala 73:24:@35061.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x373_TDEST; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 73:24:@35061.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 73:24:@35061.4]
  wire  _T_599; // @[package.scala 96:25:@34928.4 package.scala 96:25:@34929.4]
  wire  _T_664; // @[Main.scala 41:50:@34998.4]
  wire  _T_665; // @[Main.scala 41:59:@34999.4]
  wire  _T_677; // @[package.scala 100:49:@35019.4]
  reg  _T_680; // @[package.scala 48:56:@35020.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 35:32:@34905.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34923.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 39:28:@34932.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 32:18:@34970.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@35002.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 73:24:@35061.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x374_TVALID(RootController_kernelRootController_concrete1_io_in_x374_TVALID),
    .io_in_x374_TREADY(RootController_kernelRootController_concrete1_io_in_x374_TREADY),
    .io_in_x374_TDATA(RootController_kernelRootController_concrete1_io_in_x374_TDATA),
    .io_in_x373_TVALID(RootController_kernelRootController_concrete1_io_in_x373_TVALID),
    .io_in_x373_TREADY(RootController_kernelRootController_concrete1_io_in_x373_TREADY),
    .io_in_x373_TDATA(RootController_kernelRootController_concrete1_io_in_x373_TDATA),
    .io_in_x373_TID(RootController_kernelRootController_concrete1_io_in_x373_TID),
    .io_in_x373_TDEST(RootController_kernelRootController_concrete1_io_in_x373_TDEST),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@34928.4 package.scala 96:25:@34929.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 41:50:@34998.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 41:59:@34999.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@35019.4]
  assign io_done = SRFF_io_output; // @[Main.scala 48:23:@35018.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = 1'h0;
  assign io_memStreams_stores_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_stores_0_cmd_bits_size = 32'h0;
  assign io_memStreams_stores_0_data_valid = 1'h0;
  assign io_memStreams_stores_0_data_bits_wdata_0 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_1 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_2 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_3 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_4 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_5 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_6 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_7 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_8 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_9 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_10 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_11 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_12 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_13 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_14 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wdata_15 = 32'h0;
  assign io_memStreams_stores_0_data_bits_wstrb = 16'h0;
  assign io_memStreams_stores_0_wresp_ready = 1'h0;
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x373_TREADY; // @[sm_RootController.scala 49:23:@35125.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x374_TVALID; // @[sm_RootController.scala 48:23:@35117.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x374_TDATA; // @[sm_RootController.scala 48:23:@35115.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 48:23:@35114.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 48:23:@35113.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 48:23:@35112.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 48:23:@35111.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 48:23:@35110.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 48:23:@35109.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@34906.4]
  assign SingleCounter_reset = reset; // @[:@34907.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 36:79:@34921.4]
  assign RetimeWrapper_clock = clock; // @[:@34924.4]
  assign RetimeWrapper_reset = reset; // @[:@34925.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34927.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@34926.4]
  assign SRFF_clock = clock; // @[:@34933.4]
  assign SRFF_reset = reset; // @[:@34934.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 57:29:@35153.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 46:31:@35016.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 47:36:@35017.4]
  assign RootController_sm_clock = clock; // @[:@34971.4]
  assign RootController_sm_reset = reset; // @[:@34972.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 45:33:@35015.4 SpatialBlocks.scala 112:18:@35049.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 106:15:@35043.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 49:34:@35023.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 102:67:@35040.4]
  assign RetimeWrapper_1_clock = clock; // @[:@35003.4]
  assign RetimeWrapper_1_reset = reset; // @[:@35004.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@35006.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@35005.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@35062.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@35063.4]
  assign RootController_kernelRootController_concrete1_io_in_x374_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 48:23:@35116.4]
  assign RootController_kernelRootController_concrete1_io_in_x373_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 49:23:@35126.4]
  assign RootController_kernelRootController_concrete1_io_in_x373_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 49:23:@35124.4]
  assign RootController_kernelRootController_concrete1_io_in_x373_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 49:23:@35120.4]
  assign RootController_kernelRootController_concrete1_io_in_x373_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 49:23:@35119.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 77:22:@35135.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 77:22:@35133.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 76:18:@35127.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@35155.2]
  input         clock, // @[:@35156.4]
  input         reset, // @[:@35157.4]
  input  [31:0] io_raddr, // @[:@35158.4]
  input         io_wen, // @[:@35158.4]
  input  [31:0] io_waddr, // @[:@35158.4]
  input  [63:0] io_wdata, // @[:@35158.4]
  output [63:0] io_rdata // @[:@35158.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_1; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_2; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_3; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_4; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_5; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_6; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_7; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_8; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_9; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_10; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_11; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_12; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_13; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_14; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_15; // @[Instantiator.scala 53:44:@35160.4]
  wire [15:0] accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@35160.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@35160.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@35160.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@35160.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@35160.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@35160.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@35160.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@35160.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@35160.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@35160.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@35160.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wdata_1(accel_io_memStreams_stores_0_data_bits_wdata_1),
    .io_memStreams_stores_0_data_bits_wdata_2(accel_io_memStreams_stores_0_data_bits_wdata_2),
    .io_memStreams_stores_0_data_bits_wdata_3(accel_io_memStreams_stores_0_data_bits_wdata_3),
    .io_memStreams_stores_0_data_bits_wdata_4(accel_io_memStreams_stores_0_data_bits_wdata_4),
    .io_memStreams_stores_0_data_bits_wdata_5(accel_io_memStreams_stores_0_data_bits_wdata_5),
    .io_memStreams_stores_0_data_bits_wdata_6(accel_io_memStreams_stores_0_data_bits_wdata_6),
    .io_memStreams_stores_0_data_bits_wdata_7(accel_io_memStreams_stores_0_data_bits_wdata_7),
    .io_memStreams_stores_0_data_bits_wdata_8(accel_io_memStreams_stores_0_data_bits_wdata_8),
    .io_memStreams_stores_0_data_bits_wdata_9(accel_io_memStreams_stores_0_data_bits_wdata_9),
    .io_memStreams_stores_0_data_bits_wdata_10(accel_io_memStreams_stores_0_data_bits_wdata_10),
    .io_memStreams_stores_0_data_bits_wdata_11(accel_io_memStreams_stores_0_data_bits_wdata_11),
    .io_memStreams_stores_0_data_bits_wdata_12(accel_io_memStreams_stores_0_data_bits_wdata_12),
    .io_memStreams_stores_0_data_bits_wdata_13(accel_io_memStreams_stores_0_data_bits_wdata_13),
    .io_memStreams_stores_0_data_bits_wdata_14(accel_io_memStreams_stores_0_data_bits_wdata_14),
    .io_memStreams_stores_0_data_bits_wdata_15(accel_io_memStreams_stores_0_data_bits_wdata_15),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@35161.4]
  assign accel_reset = reset; // @[:@35162.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
